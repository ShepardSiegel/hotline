`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dS3v13m91EKVaf1cZDQOl5PZ9hu6M+f6vs0XE6ZWvu4T+k+BsaDsfXtA5ihuy5KziaNkS6EeNW9N
qq6Cir15IA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dFoKncYoLhQCFssB/O8LBGVZl2al/XtfGRmTA9WNIm+9uudHEd9VUzCdMJ9WAcxdxzsCxxkCXmG4
HHDzyCVhRZTSBEhDdB/aCFxrhNPYuuQz88IhJrhQ5IAlVl2BpBx2UdUIvlkGeX+KMSQB5YIlcwx+
mnw81zKOcZmKX8fMv3U=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xV6WOVKrkapwirPsVwTBBGAm4R4ZV9aoZSJ56oXmvm86Dn/qFUcnCnU3+EAVe37pLI2Jw4ylE2Xx
jd2bSJzVYPThJaH9QfEpaC+XnByGv9t/GnuHEEe5VrT6Dhvm3e1QbKksSIyRPhJlca4zTb0MT5/f
DDrJQuRgaLo+lvWycaJKiwDZgc9ZemDCJvRcVMywJvS92cs5yb4Ney6Zart7AvERqsFQdrxzzx1x
RfHrSi+eppLUo3JcwherB2dtyfudAMUj8d3GJ3lYlbEd0Zw75posY3L5nuZirVPQyjcPl9PQq2Cf
K4/dmfiasVrAt9hBbZaBipwzr09v2R36A/nwpg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HRhmdAtVhEQ1M+I+vih2I0W88e57CdYxytHMiv4Xhi1gvAIxup4cMyjnXNJ+fDagL5OxI68A8OBw
zxtR5N0hgCJhG2RFvqkd+lszkT9Y2KJSjB/t9QpxwxSV1eCqtO8KDjxK71E42KfXKd2xT+wg71hn
BY4r2rK9oc9nmpB4fhQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EYyOedtb8XVpgZbnIQAahg10Xuc2KzLM/2egI9YvLUKuuzec9slr30sgN0FyyaXLvZb7qsRUVEGK
Qc5hvWnTPE3AxEzb2iwwFuREOKtxDofKrV0lLddr3YksTw0HfIY2EzFLdF9yu+hYe8/LURWW0q0k
SFa9WehtkhguB8K4NaVwSfIoblptpJo77evw7UGQcGjobWTaN/a1My7w/ME82SFsPa/aRucJjOqY
D/Xmc39BLi/dfsLnsE0oNpGSAiplCnl6tMBUH0cmsVsQ5NGfGnfhLLfleT5u3KdbnRpKzQTtcQwm
gLIaq+iYNKYSrt50K9Ayc4rZJrtErg8ahUFWRQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9408)
`protect data_block
azzS8fpJbwF1jVym66XZy+Oend1bu9aOxANoikgF3M0RmY4CEWjT8aZYy/Ezd8w/ev9AG1iApClz
nKx7FOffLfeINoraoYtIe5VHqH8diCff9+JxwmhBbs55gVivjOY00osJYNcQHnbuwWBiGTZaL0Sr
K8dE/b1GTWP5sPZb1ImWaHPaqBkQeSbmORuMaTZ/myVOFTwVq/2BpOgtewAK2pBaoBSmpTf2cDI0
rVRom93YEOfLRTSdieYeOI8CeujXPEQYzb1VQWgRb5rqOyWmg6lkezb1+lk2iTpSmDklEfBJJMlb
dI72TNvljcjelCw9cadGGgxaBUnQPynXY+WdzsjKWJYkwqiJa97orXyYeqC+kCt2B2gAKQNbdaSR
q3Td8xk755bDjowakrPAUKO0K7HgC6ZIoKrdjUvQyMfk9uFstAkI0zpbwqDdTt5LchFlQAUMfGZH
JcmYyVRVJha6QQEE2QvJtN754gruofGHTx8Nlws0rxPBT4+2asT29P7nnzgfBDSNcrbYsQ0XOupw
pZtKylaIf6xjlDyE0RrMxpyjRzN4TqUMCLPTPldaa1p/RUAzT19XKR0PLQGBfTgBQz9rMiUm4MBZ
GicBIfJeqT2NGyKjNb+lLkR8HYzTJv6RLsi3WW9fIaGgX2AIaSGsThq9SwwuBd8mbeR9rVm0UKwY
uS0TpbKfcThRJFt/ZOAbM/BJDp5waLxRS1K6NeNqoSptTotSC+otWzaB7iN84e8sT7OHK4qGOZc9
6i6RjhlVInTVpE2TVK87nB7Aj9HfNcQAMVe+0w8ZOH8tbqCL56WpQtjNSAmKw8lBf3flu9DUwpl8
jw+TJQUpmSO2JVv3Xhl5SOvw0ix7zKdOkItNxXLzf8FX1VjnNJvuqfd/r24pXbfpJ0nI9OVQU2Vs
F7i7oMIH9sSx1cavrRUCgt3iEu8d3hnovpeURrxPIfxlhh6wLf2WYEW0BirhRqsukyzZVYOdyQ59
ScS77YUZfn7vR0Pzvtkrw2Pc05UdbUV7nlSI7UZMgQU9H3OzIv+G3qL/wsDcs/UTFjF097Bx+S23
Tjxci5LzQgPT2BPBvUxOxENJwea+5y5v9Vmi71RUln+zzLTOIj38g+EaPkchLF5RLAucE3BPuid5
Blc7NgOTnEpGLyfp9aa8Jsk+BcX1R3msNZHymMDW0jIu4jKL9gXfU6UqitODRabdHE47zXKXrsDE
HSMFLXMwa4Mzs5AHqnT7tyfu7eT/U6TvFjPJej8hLjNxpTQ13az4NWCZLrDq858RdukyHAujZR3w
CCMR/XFmR5FwvUtcUujz7pGer2qbDJWM0fsrhbDyIV0fKXICZMH56exsHGvC2sSCLo+NC+iFGS7H
SdPg2sVhUzaOJc7PPJF4ybR/MJbZFnJb9xjEU+gay78XYTqicINAlTfSOTCyNrP+++PZeSd5Anei
58o1OGl8u7Jlf4ss1jnrdh9z1vegyaQHFap3Yb27GDW0LMc6tjjUnfnIxUcu5O4D3sAWd65DyKJP
xpUhEbsojPr9OZUr5FosMA5Y4I8xLstlX+N+Jdsoc7pGNlyl2Nf50r+efVYQtl9SVGTERXDyrF22
pg8F+syKtzmOAj340M7gfkdqRHgLfzTtlPTQONu1K9nc5L6lZ1N/StoCm8HHTXK/U2fiduq/BcsW
1LbuRNFdN69SNU57LJ7JbCQgQuS/3yn8LIv5Md5jRzl823EDxSKJt3Z1cEeg17Era8fhUVJSlG5n
5vDYBSB1+nTcI1hkO5o4sXwVzD2c44OleYTHkq2acAYmrdHRHzBl/b9egu9g+neEvEdRmqjws/Sf
W7PD2hv9t+h7DJ4im7TX3x4T2vP3xyMKXmxHTwDLUYHFvrRNEhnIVWqHzH4ik1j3MVCRrrZEUJhS
w8TPgorQORk4pAWyqIlmQ+saArPBOMRWmOL5EymxvQC7HcNje1mbuOWIV2DDUthXZbDyyNaDnJvW
zm+fcbKkmYut+jaGJwqvr7O6C8z97ABsGk2r6cPKhqdoedurBU1uAa5BlHsh3RdShTmpD8rdaYad
+yfoohTffkT57QfikLbPDdmNHMX26rchstKzI/mY6MJeFy/FHmI/E19NmYKWsyxCrnxnofOwWGQh
+KH41/pgaf8dfkmE5vl20sUNMsP/uUiZ+GkC+C3Ok8StT9CjbkUH/EnIDMONS5xLKy5HUHZzYzfq
EGzvvo9ORE7CMsLpb20OIUABC6rnwlvYSDgOMCgB6ij2AW95uR4wL9/SKX2bWg30dxji3D4j2xLS
Qm34COPANyegiuVVNBLrgBnrPo3QjuJatFe5HxQVGFF40GrzwjH+A6mEdlau3gHA3CvbUUjc6pPj
S+jwxxho50NbcrwSgi1nywl8nNupGldER9GJ4OHAtNiQFYwGZP+cHmnsCKEGolIhwsB3ZyiqW9N7
fbxIEed23zCFInRhegnM+u5zxxypqmrsYq0iXzoyClxjZlMzieWYDQGXR85+WRw49wwHQi28lYet
JVbDE7TyXDCQ219hPS2oe5hsJYA+QBB0UCnUJ5mlr6E+R3A/TBQjF25civrvEQ/dDDn7Gb5IXjWU
xlZeZQBEZb0vBJNK+BzIhDvGz/RmRbwsKloCfdTJ4hVualN/aYqulYUryI2R6Hl4SgeM2TAXKAtP
78KWI1iJyfQ335zso7Uw78lTf9KQvhdRlmpwKXKxKVzhr/w/3CbyV+stkKAr2Q3ZCVW6HONVIuch
2ssvHSnG7ISWXoOu508Pyh/fMamk7Wr/Hx6To79LD+IM6ek/WXhDTJk6m5FW5ZaxTB9Ib9VBtGrc
q1mnt7pyW/HSKDFl1HelvO0k/3psgQzRk0uT34I3V/y1WwMY5CKledXsFUjjHOez6BicYT4btWMh
Oru/5cAPIrs9QVUoM49Oh4Xi8+vpjWydTH+XLfT3U/DAQjurg82y0suD618oEtpV2qSp118T4qwY
wsv3HZd8oyxTJQjoQeJbn0f7BKNoxoCaft5pb3TQ0/zDUUcLAV1abu577yycxyGkIVXm6smtZmVE
CWk0QLPNDTbyVOqx9PshtLTXjp23R2DVwlM3TteaqqBT0QAmTdcf09qt8ItwTP6qnwNLatWEBtlK
jWEcwsAO61aYTwe6Uye5sPhead4v8NC/38myqh4ceu9bT91503QvWeizy9UmVT6KKuSnP6vHmVDL
nAdupDwDskipG67oDe4dj4bCeovpb4DhBQXESKMzD0/spE/marBbGwj0qnUoT086OvPVN2TXxGv6
Ve7m7XyEtJkm70Hr1N01sYAmXEbA45Ke6DNhDZyT9LpWNjhA0gtSY8t1/XbRdLzpq+Z4o2z2Xdpq
ROx7+k50T00oN67rHZGQbB07uHXs6/VVXtG6XxfUDuq0JQUb1gDc6Vew/FZ3LEgjdMGxDfycJe+8
zdY9QhRaPQ6Op0edE4xkJ+pOb/agj6IMute2UTmZifnZl5T40TI6+xpX2oB5l/gbyLgH9q2txaul
WWXK3Jda8dyTVQfmspyn+tzbIh5/LsTYq2JkFYvVva1PN8JNR1DUUFNMnXsSyRgygUFwnS4PbA8s
FlQtuzUed5y4SEI0vibTebGrMt5tEX1k7Sn8fXJSdB/PfyEww55tyL66eZoszoQVG/YZ6PAfxa8r
OiJqL8coQkJBXOpLaoKkZOB7vPYO+Rv7NdCKxxle03JNQdnmdki//+0qHXI2E5iNGGHxS2m2CMu5
QD7X8KDm5dKcISxjv3T9McL2UWPyiyfr3v21hX2KLYbpHUhU5tD9mNWnSSUFYWqLRv+pucTlqKh0
1vpU8lEy4uFwDCW3CqBKJFRrrbc+wdT+oO/fLzVcC8VTsGWIrg/ip/Gl6xZVQxN4V/q5bB57zAJ4
5nZBiDLti5BHJ+Gk6cWw7+VIKZt5m4++aIqMzFl+VjlSkCO8Ru3B+V4jHFBnz4Fnpqq4x+cpjPFV
c7P7buaBpJNDHTz6cvaP/mgmS1DRmMwKAA+o6E7EqfaOSX77TqXDO+5Xp9yqbxXQOU8h5JYZwaDc
py0BS8sKlY7OQ6tkg9vsLUSk0lM4VhvYp/sTBQNqxN10fO1i9X0Yuju33Fw9oCpWAiJsuTAGN2RO
NBPffMgwLJYLg1xxtzPF3SLcSh0W2NwEdnhPE1OLnHKmZsQWcy1Nrm/mGtryxAmk3zewQz3Y6piz
JTzmkkytMuxQ/H9QZMhyk7eJrYqShLACONsZMD6fo76Ts6Yne07SgOHeVlks7XC6VgP8eaBJ6hEO
Kbx/ocxFBR/zqkfhORvHtyR7WhFRIOWnQ7jd9x5Jqv+TaSzFVe9dIamTcgZVhwE6cD9k3BH0PBEb
gRLnwnQhc2WccihBWF6lWAcKXqV0Tie9ipLFs4FaeaonlE8amtYUuZYg6QLLoZgMeyvkaHholjFp
wmcCQ+0fH4d7G8Q1+aaJeV2H8f2+eXf73l6DdjID3Tcds46mKL5KKClCLXOgSL5i3zz2RCQtMhhQ
94Kcs3cjmtcrO+OZihrsRRGvCB7HosknhnEnAi8FMJhlCuRDTE2FPZ0LPURFxtHvtr5s8aT3Pg3w
nMBHliGTPOzN+qQTX+7un7eF2hasli95nuENOBkBthmMRc3gXzP9Eqg64to20QmQ93vd0jRed2iV
ttYjqW75dKoJ3ag6lq0SdnEq1nR5frEUZXOfaAfPbD1OVcfTWbyK0BolQw4+W8PJbg/13Rj/YCN1
OCQ7t6JWlr67mGW6aIMPGNSpRWIPeH/7ZW2tCZupoJ5gxwB0QPS+R31FfifRZxDGAST7+KYmSDGu
xkn/keAJ2kGZL7sRFTYnH0EfcALNL646YRVAZC5j0SQncSCopX88Q0IGsHd8oDIFTkmiAm8tvmFx
b0Yb0hOWyK6DuWlcCb4T0e/XLGMsymH+PT21UJVVVyn336/gHlk8yP8c4UlknZcqCmAItevMoeuk
owk+UxSsQtT8v0FUHluE7T1AYJ+sWd+PFj53mPT2L0eT0ycBRQ/HYzBxh1RYziLOeJzkRxVI6zDH
YaoHAd3ozc5fOxiFyNFRNEP0vRbpq5VkpbYi00PZ0LhCpfujP03ClZ51uGUg8bADF6wiLxofecBU
snSkXaq3Vk2n2OXytoyTbcSSafzAUW/BUA76y9kZ/ViMIdLAA1d5eOKxRzXizYemvyCVDaUnulZ2
8x0nbi5fmTts3W+quNpzPoKSdVrHBJrbkKL42WuirdayysSFCD5cMJF3IrfYM7DI9conH5Em2JYR
FXWga+3I3/TguOyPaGOdL1wgE/7rXMG0zJKNuXY+kYNRVeTgQilUisHRMieF4AgQJjD/xRbkUbXK
YywvRLMLgnfgKPcEAMpLBBqJt+wCuEmIW0giWgrreDqVLqxdJZ4eIwhPSFVWnXe+QGkGJYAowwrm
n8V72IDgC7hMKpTE/Pxkqj40lfCY4kzXIFhKf8kJP//adBNdr4GpEieIcCWFR6EhtUL+p5QYmHsJ
+GTA998fmMHgGOqTTyPtnh5fgAYPn/j9Avm8lsleji8SgK0Tf7PNAj78+xxHbEkqOFtV7ipR8H5J
RISF+Bk84x9CN4P4km4KAw7h4eVeVfPFv0UVx9qg8+3gwvE+hcKtWM1sj08em7zPIHvn30afGj+b
jUS2iV9vgjJ9w49sPQCwuAcPwNl8ndHefyMSrfBjpQE1ljdL8NMeQXyzzrdz3GJNHTB75f9fzHTf
VTRh4gj4/5m+OICAnroDAm61MLZJtNK2+QGdyfG04MWj/x4snNM0EHM6xaJUAkoid/G9fzoQmbY3
8Hy0LE29eaa7spK5sHJn+r1AIETFUjvkrkMwDvBkTrHPo3d+yAyX7FB9tkJS61iRuZycbsYvjto/
gpqp3GHAWsxT53ZYN7Ug9xqVya9xOhm2tzYDNUmcrkqmkv3iYKwxiHZs/AA4g1lnJDlFQDTmqUtr
BGKpdmo6kM87TyZCiTJFSGG9fhjZVMyAAkAD2F2t0jHzxLjiz73o54dYQnaXAy9ECjpVueOGZTTQ
juqOKxH5c/80xTyJ7+J749ND5uykphje8M4gML3cuV0xUvwlk4xiKAp7Imd+phFiLMNBPFdvC2dH
+FM6YJPdLrTjc6PWhiwAmaNzOEao5CO86v5M2Vc0E8S1mfr5PdK5Kj984ctgsxTFdSu3E1EI592i
uyYjbuMNsNWKpp45dckz72cVmjupHicDdwrvNLDaeNwQ8Y7mfRoqB5t/UPUkifvHoAR3fuy44Qlh
yyB/oMTkgGH+TTNqGUcU8f5bTn+vzKa/llljMa1MK3JPuTDessrMdPKaNuTlGBHduYPUKWjKjmt0
RP3aTSUD7BzL8pNkSSyEzaHv8IbDq+Imt2VrRaQD7WZGoyondsT6jTiWKiTFo4BcXNkxMTgo45na
n5++DfQNfG0cR2sCVkpdYo1OJt56uNyXX70ZG3get3jd5+fKhFm8SXUVB9Wg2+Oax46dZdiUKFdb
m4A+4Wmis0eu2gfEDYWaLJ2n9PXG6oRKaPrfnZwRG6rsAwmtWg6ouHuH74cti5+HyiouyWlgG2pO
IK3/gIv020rriTqYSSHUlMUfjmGSBLR1Nu6lPLxgiELS7N0IoqpuMratLus0MOPhB75lR117bjwN
1JHuoaZ5PYXwqWQhZ693ROJt3KAcn49WdlFWLcItCviRs9PDtnkME1cdIW11SJscsx5tEx3KyX24
r+292FzrZ0si7VvhZJnMcnWRAdPgyhjlIFbn+49xTmzek9rqGhBP3Qpf30tmPnBWUmdmFDlUHGNL
ysYcpEs1KbfqMXNj52SDf7j0WKM/takvTpsgkgmWA3I1AoyqK3aKliAf0HKG2SSViVdg0Rj1+QP7
iwNVaTpQXjEVyLj1/3sBGmbA9SxtewGWChMZFnMCTUOtq2S/SZB/g0SpZ7GikTaCFQXUFGFb2CK9
U/pYvRM2N4XcHK+xfqjVU9eb1HSlAhv7n9ulMDWV1TdBdAXg44Fmrc9WpFX5kzG4LdtT4cMj4BI4
K2gFjvRgVAjBKfIIOzt7ccLbY3yfy8h30KOb0VYRUD5kYeUxupdIcVXDg736o0Q+0+qr7RvpW4NM
vl2EmRu/hrZbPwCFoLHd3QaLzZ/Di7xjXlnKgFsf/DcTuwuz/L+6Bwe1nKupH6z/6NK5BIzx9GSJ
cOuXrGFE+toWW4pCSug6ftHhvvZ6AVtnekJi+s9kXb7jbPV+OdkgnQdXtLSjB172OZx4MuRgq64q
6jjI3Te3fMW8kG+fWi1YlRFJiWzB+tpu5WghMfSnx+0GQd+ZwFQwjJSI1/vxdcoyfOBnzqzLAn9p
0tj8iIOs02W8zPwQWKXrhx+3gHmzAJ3OKMIWWU1GzOTpteO/qJVdt9JkaEK7QBHgHqdyys29jA9W
qfvxNIiQnEwPGKQTGyg0ayLM+Fm8cO14b/FKCMLnjT0SgAp9TE+3yBYJS9exMbYD34FJMwgImM2y
VCkFLOpxvJspBLTQB4aioSUc+u1BS9HWtbyO1VN1ExMV4uy8iiq9Vwu43WVMKnIqpLvCrnDqoDdD
aUaj7bZdho9rq4odNCEvG6gQfyBXVZRN70uOjbbXFcKE4scbc/qWqRtQOYi2sulJ3DGoEuHqkkHz
+T3CyI5/p7DKj3rCCzYlb2ffhgt12FwE8klb/ZPJZJYsiNXEsqVF0ESef699PBEEX5LQNEmBdweg
vZVMnokbY/dBaafOHuN860tQVUazrJV7ZxH1FO0xtI3IjTfGJW9aC+Rlibsj390WEL/mFVg2t3s5
+f0plJU9syxMU/rABoOlj4Gi+ThWrUl5vk8u/clEVhlYfCImqnoF149xEufwxPYJIAJPJk/9K/1S
G81ySDeFgeDlytJo5NpMVQ66HomFps+V45UgyWOpt0G5iIs1AtfWB2HBS6PXXuEVJ4rbS4pzl3Mq
2QGKl6kBBTsFwMeJzMy7ZoW3QGoX+iQrXL8laZiBDza7m/GKM27tn/Fm5Z5MpgH2h3ca/eZHq4jQ
wF9L4yXCt8WMY20sEdrjzmKBCqt1cisUNZQisezz61DTgJOV385qSHFpCnd/CJaUcaqzfL5XL/+R
7sHCHB3OWT9NLKP1Ymr4l473k0aZU3KEWIiPntvIwoyaJ2p0icwtQl6KGXNPxQp4WUnda274AGLR
UpjlKFWcti8/0MmzL8iZJqLceC+6gfVZZAJYlAIzLluHzhW+2WhUEBEMJhkpvy1/1prJGU9mcPAA
KeESUIPvp44crX3PruGmeJwHJVnTKMDex6YijjMHXwqUwvgQ1LI77RtcsquPwTWqWaLr4k8UEDhO
b3NOSyHytDSkSLYijj+9SLdwg4soGzRwooS13eCf8pZmp0YiFR1iNOsFih2cDnbZep+Hig92P5Pp
LS6/HEP5JHbssdi8h7fYKyLMl1vVNwkF4PG4ErAUq4vm3X0ykoKLofnn2mOLouijc90PiCTzk/6t
VA4u/W/sx5b99k7iLUOvJv3RzweMGEew2VAC7a3RPz7ha75jYx/HscC61eBhMF6dQriUSkz908NT
WwYge26JIJsmOSDM559F2THNaQdYZOlxCVD8z0m3UJS5osMWmYssl+FBXbO8dLIaaohSK5CJ+6Hj
LbGUM/CbIbwE2gT/G/HaXx6RwIxkFO2H3nZO5i1SlNHCkvBPV6cJbAPn8FFoju+Jp3MOydDHUqK4
rGqtFrBuTkSLGbfLJmk/YwxdCCCh/gDWRV6koxq6KzDwvluivoWh1ujCDn2i6Lhynl1W44BqKKxw
2IB58zC40On8l6dkfxbhGSOk1fujrTPU+vNIdetKDyZrIjaf7xLaDtV2FoWiLtr3qH/0m20ga97F
C/0ET+4ffwHdgSPjmeBM2hP6J8xMn/SuHr9Un8RruShKWX/jRFpDnPPZiX9rwVC2mXnRDzbx2kzB
J4lrN2vg4BvF+8iygS2V+m88UFesSpwoPZj5oxmNOVmBo/iHxHOdKypDBRnewvzZ9JWCfAP62N82
+6I4o9b5VwQSiFXNXRGv/8ye0drSvHi7isbGErAEoztPGOwtgkeBXk4Hf533ukfGnAXAkNw8m+xY
UFg5ehHpHeU5duQHQh+zM/URPa4HGMpFcK19ENF438BVflHkrvhDxE2LQxPyMqBxezTwGuCmPI7T
BsR+jxdaAl5oCFtqLQvkpwTCFQ+MW/c3Y55Io+vMw7IBjpvdSYjjbp9cQrBMdnqJdpD6dqlyN7eH
ZWJ2xmfqcIdDQiNMgdUoMOsuVPyR5KR4e7E6Q67D1StRmE30AcXnmc2s3y9S6qutq4fcmU6G/vP1
dnyRPbbtiLQ7AweEVDY+SDqBRiAAtrJAiuh876ze/5X4vABtsihvyEdQ6sFO8uxfmqRnEnEQbhFV
+nnvIN7pITNgfH7pNfHGi48JIigxJCoRUMWsBza+V9vO7+WC4ZC0AlOHwm5rTfzgkRr2DRfvk/d4
2NxeaC2WPj+hkPq7NgnOdOqTzEyW0wof05cI/37OGNIMSZUSwbyGTQ21P3HwcbSnqzwSx1Qj+MAa
mHHVZOaAmVR1yFj1ICjBT6Ti5+mV+kEpFKV5xcThBW/hJyfY82uJEv5+lWqB+RDqSftKi5KwUGaH
eh1uYq93W8T8p0R53clhhBp07xpDeuuDQv99DnSEkQv+ktyJbaHj+CZzwFqID+/H+h6Gvg2bvEDv
FgC5KJO6st0DutZC9dRgYWsHbgLR6v4VWN+bbAziOqwu1AYsjc1pNimAGcx/hFVkVhLPEEemlGUG
QEj3FeeaGE5VbCiNi0Aj5kPrViMKUD1ahbyPqzSCI9lpPsvwtZuEP3DyyEcRHrrlROMaW0EqnSJj
vRrl2WTa8CYSxqyhWvhzI1PqXmWq9GN8wZNcS/JpZxWJuIpJENhwtscKF33aKBpALCB92opbHj24
O0h78k/Ht+/Bv/nJNAPJT/JppDH4VuVCvWiRsIOMXhYJEeJxcwwRawnlSHYNNrM28dm4EoG2bAyz
dhjkTcaHrzr2Mp8aYsmnK4vQL1DGiDzDgS4DvWdEIFFJaffDSdBpDvGBnJTUWJ3vTiZxTktuVgQl
ijUKFVmij98/AkFWLK/7dh6ysjYD69pgI0uFOqrmUPwEiwHLtyIYvyefKIXKu9jvE5YsJa6lHUN1
CfHNjk+Tmtr7XUcXbuTDNcO6soFW4tWyNQ1tb9fLTChWUuwk+c8EpE7j4c+G1YzSZ16i4K/RmJlK
KK5guJAK5t1uBBVhuLnPNcEthlBjUeifTRCp8SwW1Nuov5yY8T7Squ8KpQrSkSP9rdAamKSjwIzF
8uXFaW7vb8an8XaUXO+UKTeJxUVToIbZLyhShNBBvdIDC7is7D133CZDSAY1ZCoCUgMtEzWuJSIC
tqmG7OXVVGXj+9MFw3SZsGE8wTIxeOpig5l/X6/oDj02g+hAo/T6hfAtt0bkdgmQu3za/NwKJ409
MNxMKUEU9HG96Oh4SqNFBeMR6pweMLqeW04WD6fT98ElDQtsntj9fPr8Bm4NOQbdFKhpjqYLyAEK
zz7pUHMT5S7jp/LOtI48Pacy9ZOXVN93XkS2eiD1mNL2ipYoXrN9FfVqCXH+sE8O1UoFdSANvaBO
Kd7TKvpSHkkn3l18q3s7N7Ku2+6gBfn/YRjX1q0TLVOGsF6OsEOik4QwnwPNEUsmNdVXaSZO+aX/
657HjtvIy0d2co8AZPnIqXty4USNRfXtO186IvYFgFCJ5ecaQuxoQ+DyGwQAGvGXk7tPgkqfZwPL
roI5IjpqHgPBtHvN+E8MseTJMNpaPBX7sys9rnhgsS8Ojb+iOM20mIJD6rV7owftgJ5ktEdWmkH6
dJZqphAFtZ1CXHhs8OutgQd+BIZB1YmVd6246YzRwLLaYF/pKWkuV5+CzNHTKtsdv50UCPzAe0pg
0UGuCgafGFzSgdeAjGHP7rI42QoNbY2pUCd4L0oMjWKw4mnJW2BmD6Q/jYFU+vsYivqGUUK3518B
zQohhMydEyv0X9+uOJt5Pp3vX5sCcleiOUJjUx868dZYBP2imLITN1Vm7VFvZQcexwCS6l66SCi6
Lc07fqB2MLcz2aRts5UoISe2ZWL3dx2xS9f3HiRVfKNvz24u1YmEnZ5/9aWiKcVTmTPENQeGUwNg
1KGhqCxjdc2GW/z3V43PYHO1Cb+uWGFZDq7KN67ZmDCb376l4HkUG9hgPXlkFPLsklbNTbo+54CD
r/XvGt8CUWuHPj8aDiYs6QF989z90IRKDxrkGuYBsdgLNlnxcBCqh0a35YkMJy1rcQVz1VELqFIz
2oF5aFgPu47uFoJcicNP679CPxUGkwxud1nfwW6UCuhvaG2dW+UCPEAFoJt0yAVHZW7exgEQ7bu7
8eJZZ4AqDo5cWfMwjhVeN6xer4zNtxgxbsLKP05TC+cNbIiBBuidX6BsDfpzI2qP40Wa0LnPtTDt
e4S0rH1chAGLa6oV1plbPxZ72ZrA4AMlJP9Y9cewx4TxF5ldkFacCNYOLC/KQSgOZDZj7TuNBbfK
RtEQP7jUlL7xncuhNq2axrqBNWXJ3yy6xOdj86Yr1uXiNfWIQRPV6/U6rYlWFa20YTyAve2hLUuM
HxuQVSJOSoCCEMvUG1zh7zph2/5BFEpGJYotp0Hw5JZWrJldZWXMbqF71KtYu4JbC2KDxTMeeLCt
4X35tsjU1OyDblnu6NaAhQ6O/4Okr8OuuWPHDL/gfhRU4nhHDe3LtT7dTBF6JtMifjRxUNAkmprQ
JZNdZy5nrarIdxGfTMcXAZSKq/Zdqi9h/FAOBJwFqaT8JoSPBBgbPVouJuX9AuhnmsMXRNSgo7z8
N7qzMoWMpxVI5EkumA93w2pFVSDz977Mh1u3E/fRH/kSnjsnUSwxH2XjnDXpLvhmzwS+GPX0J4cs
894DDqH1554DylCtwD8d8Yr99H++QhwDHa1iil/TvYcdA4lVvFH3W7NRDutfkIOyo25yc9vs0ZSG
bT28kvWSI/5YRdi8czaQGVhX+eTdLQ21uvWc6SyFtPp1CzwAiLHgna+NwlljFBH5NsozSSccdU+z
9MHpkL65JmfjQGEjZmb8P6mMU0LKRVl800D88q83goKjaMWkKzTNFk5AgGpjgVxcehQPbtYWHrgb
PDZgk/ojEi8SOgCh9kmXbh0QxKPEq+AiU/lm4jo+gfgKR8L/4u99Q2Ra4MPaXYJEnbocpS8R/n/K
TFV5ASwiX291rwwSMTfDM0LquRECIgulJQUS+7gwkncTtSRIacQjsZ+DyeWcKtsefn3QnsWEGU2U
k4wKWZETDXf0JNbF02mXKOCtdlBKpeRMojBVAk0hxJpeCrdTFoEz2xrvjXfPB8jtHLx38E5KGv33
NoNG2wGsNnTnINqQXXe3Qq+rvIj33Lihvls2gaFmUR59mOi5c1qgKZqrY5b20u94Nc7MVjgriS68
mvsFzu5NdGiuJjxIDyHSSMtO1ud1ZGwlwODmuJhsAYVEDAtUJgkfZ5OzUGlMms2Op10M03RcC0MT
b+UBu9uihL6bWtbavu0kCuI6xy44g+R3+unIkgUACJlNnI9tqrZwzmImwY2Zex12e4eE06M89Sba
3EXN
`protect end_protected
