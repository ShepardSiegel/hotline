`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Mh5GJfDoRZ/7SICeu7NZbaflgmOeat65GJetjA+YAokZgcqMkA2voMgVCMQwM6kfoHvFr9aUlRw4
966ock9SDw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CD3ojpGsRUMLFUYMiHa97DMGBZXrwPiVV0tjPoiM9asNf2YjvSTP/IetbQuVRkpA7PvSbjKKKBgR
M6BKBYUz6p9O+NeW37lYVn8nbqG5DT/87V7Hh5bcYaFf/lWSnJg9rp778IbkdZnVF0CEqBLl16BG
FVqL40DhxPVV6Bi9Q/I=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CSaXKxvNBdPOrjtNBKpeTelIvMotvaRUREBwj4iBovMpl97tkC7VFmzwmHznSNAGk+O9C/g0m4qU
KbNR8YPYF3eSI+PSvXzUSq8dS5FLH+Ye4QG0/X9dyNtAyoCuStzj+tLcRD3Rd9svWsbZjtXLvf7h
3T1NaF5WAKpUlhG1dbNAvBBkZLo5tO+gHbg/lO++mSEySOmiUrd+bQu68Iq/a7XkIOpp5EABywrk
aZ8AeM0l4HAClWSUZGP+XGFnsIWodFOjG2WOBe7vC7pByvO38OEygFCV9uWwURi+f+VoMeAudMnP
Yp7FEw8h20hHUNjA92XH1WiILNdeEoL5llla5Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Oi3GrTiavEMq5wQhyJs+G7KHiLKVjpuISfdAdp93/Z+V6UkrFkEM1QsENI42K2aBSf4QAhkLIQg6
frFcETpG73oQKwSO8Rd5aebeolUwMBnW2HWHlxRl7Aik0Hxm59jZWbGK75oyo0haF6FSj3/M7t4R
TtXsiMXw3sqQgu56uSI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hG/N9MUK92Mgn7TJCbG69DwYWuSWVthUXLJR+WXOj4I3nwaJ5DCfbZWsPkaeI7+qTLyc3EzadZ8Y
PHVR5nPWqKCnI6qBQFqx80MmA5TGhYpXyXkyq+yIHOVhsmo0Jf2BNvNMCKYF5ybbMRMEWVAJdyoL
eBk63miKw9iyhoMZl+g+QmqQrnOb2D6wjvpd8hgkqzcIT0wR2TrZrTsffKovA0R6UFWz2plxtw5T
I90+lNQnK4xtyNfp8/SuEQN4bFxQNcEkbFPmM7zpFu6+YnTB73ZDTkwKCSXUMa3yOSPWn6cMPVW1
KS70rn7RNWauSvLEOW/R5ssTAqk4sWPZWgAIzQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4848)
`protect data_block
7OxtGgm5imbzqppVdBTj/EF35HNsOD/NgZQyfax6IMu9DlKnVBOg1XkD4FdzL3cuo4X/mw0yy2GS
oJ4hZ/sHGe5a8AUY4rOod5h2gh0qMMLGyedDccmO5rYW2u2jlwzGH1Q7P3e7AdeMfp9s+pDKX0H6
tYEv13/aaxphfHL4Id/pWBvSkk5rCY0uq7Bxfw/KfU3yEhjezJ3CGUVoGnfFhTLyHyLIROVkIQ7J
c258tpJaWfdKl7XBZoEXt+dhnO3XFJQOo01VN2mNuAtcP9yGxn50G/dPvS3YpDufRnoj93fByJ7S
b7/UWa8ED/dAgqeWHBSdUJ5pgDCNygZzEwbV9v7Glq/uu8A6FNzXcqXtBh3YY8F5joCpLNbVdm1A
yNG98JxkgOwYC2TwwfwcZrvJb3w1PCnPk7PKFBSR1pzX3y4rL/RcOV6ISKM+q9NqLtMzkCt7TafN
ztI9tYZ/rdtVs1w0FeEv2lJkghZHja8kjgG8zEey+qLShsB6ZOXBKwdve9CoRKbDpgPKqfxZAw3J
Hn4K9Uw3DPZxVOzpAOe+MP/lznqbrRxNOy/1rS4FK4h58dlcJJ740zQIiRgSafJ+rFhSPbXNgFiD
Q6sf5ilmQSeEXf/umLpuVPxEEVlCqpDV/jLeWMQm2U76kLhhaqe9D6rh8RdrEHU6ojn9cAzDUgyX
41r5udQ/K1MlbrrwB+f3paxFbXN2KQ5UM3VDKhsmxS0OCvanTz7fz0eF8ifzMcg8lkWBEL6kOfBz
Qrl+o3FylkDUf7E2tLxVzfdI5CXZdhw2mJDF1vNuoY7IMPHRVHPlGJppGOKRYshtlE/9FZ0A9oeq
jPwTO7b20EsZbDdlETpo4oMzeXsQXSRc2he58K9fOviRN6ayj1T6f/SXWL5WJ5Ehe64+wEuTNXao
IxChK1sroPg1kazDv+SkOyolPHvlPaET9LrKvci2LDxxm12SevB2wJ8cq2Q1Ambc96AsTI6Tx2SJ
WcjmNPAm2yj57ssEjatbMpNwyZQbFnc0oErssIF/gRyLkA5X6f7u9AOMGTKzStES7O3CFaogXnoQ
Nw4TOWJC1mxFYFQBcZWYHUnpUfJrRthXzMThmJzbZKoA+s5LLRJo9hzTv4gfmwM6hGwrMk3mkbtq
h3kq4RR7AxFwRT0ADkLCqvwoQ143UsDW/7sCGnvC6vj2VxMku7JqmH6BLCtrhZthixeOnpfXbjB7
8uEfgVELP1B+4JtNnOv/Da/i9YRBQ7Uj99dk3OyKJ1VntR7UQC8qJRfVelJT9IJBjJzFsP/WdUhK
9qlr7aJnQu2RCjmT/kQm1rMT03Gofy9J5bBrNRy8d65ts8DjxsJ4Wsv1ZFFIccYVI71M6TUs9lbm
sk+36O8lQmBgltjiOW8yXNzckHnv7mqWq9R95Nsj2bkhpimHRmXIJw8Yp4nEKxhLXxqk67DQs9GH
6wEA0J6bT70Y1bNT5Di9dNfDuXWPZ8inJolyX36oPdrgsTQh+xT3cYQUBMwEmQZzX2eqMcqC/APe
elKY0XBq0pSEd4C2NMBiCYkm6RnpcOGMfbf67CpkFBqElwDHDQ2rJFjYOYUJod16WQ2DfCYqeTZo
jOA25Df2VyJdE2kiSy8RJo6CAPKFdeJa20jQJRf+ZioH11tqYN/ziZpwpCWxTmejoeD+HVgkVDrI
Qi4EFO0Fa51Ywq9P1MnX92DavLnilCaSsgLuv/CfSwJ8fpHOeRWwz+ULjPPHyVE6eajfr5EIkH85
6tMDrenHVRqfQWyFZFKKwXKJtXiA8044rGnrqUHYDMuRxSf5QQA7HeftZGz4v0Q55oGyCZil4wB5
36gNyrnzEbRwgy7JZV55K7mOorrfef71/KWJGKeuk4pNuHwpzaB+bT9BksCm58n0ANg2cazPlpK+
tZ5rllE15KbqyZYuxZYF3tFp3RpUKeqvBs96ckTCiYc4MxXIDy4PKMJ8eXGu3tmVAPuOvAC9o6+b
5rDriwz/Lm3rnbnJwBKxsEvx4vpQhPHFAayjtsIzgfEpqKTw1kK9LRBRRGMvTggG3oM0dfAA6mtB
KEMR1j+tCQTbpnZniXzw/XKgBepd/gk2gpruNipCf82qeKs+VQofzmGh3b9muPa4BUlwscNrgjT/
aYMD8e4ZSfEfsz96RxNnPY84XAc0O+QJucIs0cIRBW377kwQVXiStyi/6emh9ExQqu1IceXS3+9H
tc4cUp6Jyk4jJg5lYSaeRmJuYi9v0jtF+6HcdIGT1OIPq+8a3s9djZEMN+RCdfdtHc5twnxav0UO
NxHpdAU7gH743kssDw4TwS+iaJxynvi01zG6ez2i4vNvj8ELAqpplNz9hICPNrFlDLYQMVIhVQ9V
AD+7eq6aPsgb8ZYDq7P+C2eSgq9ZMiSSwcl119kh73GaD0rNt+Eb1qAsCgqiZzNORWNceotNsJnh
iC70ARsojMtI7pBWRXp7rpeOUuk0WhP35FWYeQyLFWHH2G+e2Rvh98x/B4XB86NF1NxOe0+Em+0o
T7l/TjRH4hV7xg1b6cZrdlem2zNT9lg99CJhhd4WkcnYMNLhLU8Un8rNTJIQTbNjXTFzeD53Snrc
RYxKc0Qovsj3gM+UBPO3mLInsjLW/Xv71ObVH6YLCMC7QFDhe02fz8r90DEXgQToKEt/NFyG+LiC
8iVgQM/fmbXOkQx5u4ecHgpF5NPoHAa+NypHWpKx6kFsuu5y1lNuYkV6O7kiMyKyMyRJkOcoQhFO
F2vVroh+vqvn02wjmMm95kyp6uk8ylnWDekfTxoXXhQx7Ka5x9CpBeF+WFRygCsTqqonfB/P8nuz
jExsw3tvg8V3jybGDr3DXCjQgY4vGodKJ3VEf/A+xQf5V7YGXqDtNGRWZrw+AxQjP++Kbm1e8O91
CG3rcR9UY/VeEozAJ4+6mTEJ2A0SR0+Egda60FE5ANhr4nDzggXyngjvl63OE9oGpCTZ9cac7aDm
awUm0OygbhErza8NKHMDzi+w4BvssvBiuYD6kSxDStWhf5I7+KQHxv1NyiWlgwuiauaYdzzGLw5r
eheBRohZH9R1fg84zlxKyNBLszbgDJPAZCU1bhFqRV1SpVq/p5XLIgVKHz909IPZYApZmV0jF307
59C32aHWk4x6dVOr8CjVuF0dviOMViBvXOJ02ANw3zCngYYitSLfTG1QA6p36jWfrH2sWK+IyLaj
lglkwOkDlXeEjNujXkRm2lJr3T0yErxeouZo2aPREtATolFtPwkv9GlfM4r9eRkLcuqPG86K0SMx
sCReKFQbtiMDUedqLF/DdoxsQtcLTez5z3JfXyQBL1MO0EnPX9tQhdkfYCuPjPpS4sn3ZAEWvEGS
2inL/3B4ojDE36Q50o3Wtf6PVV5OGyULKOjIzjOpQE8b6BXEsAX85d9afNAgox2yYxViSJ+QYGGy
ZM6WNu755REMzPCmQnMB3mjc9ArIwFk1K4vy8K1AqscKh0rHZ8jgPS/o4xFTyfaf3Awv4SOHxVHH
9pB39dffhrdUdwhk6TQhzxdRtdLRkiXFZSW2hPowXMgqacK4g0balWxQS49Qks6XIc2GDiiEkdfg
coVASFbJOOmP3dHxJHQ06+Co4uG+K54B1wfc2vIfOu4LxmUU1xlPCfKWtoXtrqehl45rr569rssT
MSVJE35ShvaDLRLBc6cnyGQefxAOPXy4fywdnlqg7TEM9sbwTqyp7A8miytCOvEbJpXmXP4Q2RTo
X9GwFA+LDi9mrGRe+GkGCkJSHl4UVd+jd5vdJvaGBqcgpZ6pY1odyB1ded/NXC3F5M7InE9EfAU8
nSy9bnoMD7BVLfaWPs681aI0zLZ7Qvoy82dBtJaWfhuNJwaTox1icSjkTlqYzV0P4dh/9Z6+2tX8
lJocVCDWSo1rat6LhqgLY1hh+jkkdfRvK0g1gY71QaeV1sMyK8xwDY5VxGCaI4wg+iqbaeW8y7OL
AdcOtJgyYWNIi50eRn3l3yJacFY4hATVgmJQ8s5N0gXzNIFoabEGHnJGBNcqUGh1HIdBbrMBRyoy
FFSB50C/nYEFuP+riTgwgmoI+5wUGPRfAIrGFOKC8fO6PLKst2I6iVybKnsPXpOoxk3ECBRasJl+
tMolJeqPDB+9YViCXeg5uS/fNGx4rEin3fbhFDreRdAQq6gXHCgXm+fDh2VFPAOm1+LLjhZtuZu4
AdEBWWpcA/r/P3IEqAXkxOxZguH5QOaLR+f6lBekk21Aagz82FD3P8/36hCvUsdSLVUdUJvPblTS
Ebg3Jza003Zc4uJcaaE03Zg5esssjCqGNTYXPPOLNCsbhoDskzDDKmTXnx2RL3hNit81/BO4SFpk
bOtFIR0sO35RbB8jrnbI2H+afq5Krt1huTGpIHmI4ZFmPaYYoB0BJGMMQvlsOu6Hf67R1IXRh3Hg
pWxG7iX6VDLcU2V0cjafpCIsFuC0iuGWUsIkDSKq1+QFb1SJZUD54lZjO3JFFw/j/B+Tq0vZq+kH
eYpJs9Z1FqvvOnsFUs0hQ3u2qsxpFJ6Np1eiENOXwAGr2oiV7MfP1vAiI8mhhOfMzFK5PTuiHYjY
Ht03YnsxYWHyv9UkUcG543FxKXMuqu85eigqo1CTyuWR/r43Jyx4xrHQ37pKEQRL/cWBHtyxrRql
6WZhO9fLysjqIlL1KqFVci+uJB0yG8cAj0GfPmS4jvRlvmbBpfFgze2K4FlJAgasw7rZqUyb+Szb
UARIDZR3JSEWJwa3i0F5KPMrLe3bul0Iwj47XYFrxIcUS4yCXbLpMUmvx4YLckruWQ7evW+RuZSM
JvYrDjc6SMMMX+1B1PIS+xsL8nikhNi5sYPFbNXiVFYSOf3TbAh5N63mFpgMiEHwhxP9ai1zTMXF
ruQQNXNUYG74C9HxVGO/qnqr5JgL5iEF7TQsYt71geWBRnBiDEDsjtgfw52iz1kZBdPtDebCh7Hy
8CF08WLzizkMhTk64Oj1Rv79GTYHAeZxTKOT9yrdGJeF85J2xdD9xKCd87lQBo8siGM/k6xMASJe
WMLC9xgDe//raqEOhqo2bModojvuDj5SEeiqjr6b2veSnVqujzhnoKzckODIYLc9qxu7gEtUKvmY
tvbQ6nbMhQ0zYO/YC/5ARZh6fCtlgZK0vj762M/Bq2O8l/6oXpaZ6EFGeC3MYDA2afGgdRjKZZCj
QBkTdwnzMuVkxDKZPPKypzYjcS6VhWKvNpBFNrYtAYQ6LIhmx6OhD6GdMM8Q9O+SJMWhe6MwLg8E
xUaU+vAHDMWY+FtKcBE0DHMb0RHCkhe+EybMn2r1WHC2Isv6HB3ag2nQVD5VBFBbHpmjKS8qCKS2
6erq7B1AtUbQ6rsSDV14I5CuJaETJsMp3Uxxt77hzgCIYnt8eP+S3aIO8ZDyMxltJtQ6R6TBeZrJ
Iu1efzlFKFXYPGGft3IgUwbhtig2JUHuupAi4BhoBIO19KjkvDCAnHYr8GuMB23J3CxvWXAgmaYw
ghMvhp38ZokCwyWdKOuwuUGwv/YMmSppCKHZmiK9KGdJkMC5iVx/lQc5p5R7TcZlVltOd4fvTY3P
OkFsE7MbU6+/1rPM16v4lzIrLSpfZfsh9VJkha3FALuF4C2uIJl0jrGgbMFUivPzRGdJ0LtOhqTt
ARD7zVAwMyfY+mS0Lj0hDs54Q6ZKx1/iIER14ELp3m3j6XEfrBNbmHdb7wkGD33thnD7KQnmRL19
YkTo13so4ADs85i3/A1Owyhx6c9TQIesLnbEacsX1RwlIz1HdY4qStjDL2tkJd5LHa1JTq91TyNu
ztyF5QvgFepUYsJum7TUg+c2mFiF2dqqqZJIlx5wW5C8qNl05kzbFuy/ZnISudnkvxVMSZ9Dilq2
zwk0GUiZ2lDs2lVC3/ZBpWjEOuDKmh8CjOLIm/sLbAP8wN1zIyzsjKasVytRJhDbNI/VaMT5/ex3
pRoU9dSUffiV2n8aAeRND9apQMFFAUngra/190fnvoJhNSiy4CEm6wELJVJMek64/4TTPJpwmHYl
XeZpyVN8y7kp4jc07l6gT+yDW4z3yHbY89deI3oldA/NctaLNwgA7Qe20V3X5GL81KUQ79Xy2GSJ
riSyxJedqmHP5w+KsG58Jl19/5tuSflySEba0oVQHArYRDSla8ikLBj6oZS/iNoAi0o9p/chorZC
5C6BACB/dfiOlvC9kYoTHFAPDc3q0omROD6cOE+DLwObrG/G7MA9A9jwtEh9nmykr3N115rmtrEB
sQJx/4Tl5qU33beOPDz99PKUmxDVG3v08mRyuBktj65R1ZS7UDt8hxsYv8neReuYnUM1okJAzgwM
J/W2VOz0IVPq6URMgDvMNfOoaQFlyHyNma5qzQGGkxPodtquoF8aUK1zALzfl13hFFNDWYrMzyDz
p5rZbbu0SUyLbt4CfsOABR9d3jt+IndXNR/9Oy748mquNr5maY1tNiJBbt5Nyz9u27yqo7C50NpS
Sf0r
`protect end_protected
