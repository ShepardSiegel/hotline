`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pf7AqHMU7soHjlgZl/8EHyXl6SlqF8iBxfHraRTjI4hRUWv8B18bxumhF/nGEJwXC8adUNKRCmZF
mCAfG4FvIw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SG1/TnZn/IomAyGMOvSFM7D/YlltZatwZBypiYYScEQLxfh+6nlX152KB+ylByTZQCiWOFWio5E/
Mt6BhPZIHbsQPl0Wa9oYkzw/iJOdP1sNTC2Y6VV+voC9JHX0eJ2vPByJAkwMwcKj55Vc2kJ/SJ3P
9qKcMJ+2FIRE4XqIrsk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bhmgBiuDTdgMQz9ZzFcUBPzZfRnVTvOetUpQ6VxgWyuPLspOo0nj708Hz1q3dsQ1+f/1byG6hKE2
/jvRZDgT4kas7BebxOpQENLavzDrsBrOyD3JOKpaOfE+vsqUpVWTOLACpZ9Ll0jKIipGN2eFM1EG
eZT5LWJBgCx/EzIx/UQgujdc0djb7TMA+mCVT1eGdyTcT/JfppmWMvhe2nTmHKc+rssO5kLFrJAm
esulV/D5TC6piJhgw3UH4bNImu2wFK4WmUUTSTechHqhoVsQ6RNl0AE/ZWKVukzoSRmQuXTAPpWu
OpAhH+MguoUS3HvKgW4EMM8lm/jhyIRnzgycyQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kAtHj8oFtREwo06CRqikoKOPEePjQrng0CQQO4bqfNMIqADu1EgItLfjW6fHzLQYPRUbEd2WMBDa
GHCr931/Jp9gER68ClIvXW7rGTd9y6Ty/ITKOUQwxa9gTQPd2EYWbrv73rI1x9j3bsnA4ITL1Awu
MEUtjIQbnKDbx9Dmh9w=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KrBm+tTXqQj7nC82qxbFMPD+BMYbhGTQSRZ36eCBHXbxkcieoY7pxzJhnES4YMqqsDZy0A2ZMg+p
xPtitUkI8x3tKBkhZZ5jUCIGLye4xxUH4AlR2sNPsAyCMhFyoZDezH9Nss/v2xucWsyVRlBkd3zy
Wn26SEnj4sKbCFGMLL96BCt53IayNzRkIwF9KHzeK2UbK1tAVuX8e1wuYMVIQmCxy0o8z2Ag6je2
4NxWraPE65fP0BPoTGaeJoDG4pc79FjWeFcQT+JnJ9F2oKfyykz5I5qjBpoqEQINLD9DTrMKjSYT
YuNfPeX2OTb7g1LWe5KTrMwgQlt5r1cCJpGL1Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9968)
`protect data_block
UQEmxd4s8uM4tMmGg5v0DtFyjEwCMlRBKVQ+SIArBy2qF9RC/fpM7mMK6cEpqi3yFPGLw9OAvYQR
hHI+EPxypIUIEV4bXepYFaZAhGIMcV0CRo0XJLlEE96VeX6DqGVxTo+QKepe3SPkCnht2nFNXDRf
AFP8gp+uyed1wnKvDf0QBSlWiIPzuk/SVFYGqFqQXo34y2ljKMGsB7Q/U1SCX3XH7k4R6VcCpjFV
dhzR0GmT/eaQ4sYLXLT8aZ2mOagfXhbrods1jEFUnvfPi7yTnIFKt2BYzMGKk+BZfPys/i/sSBEg
rjWGJNGCCxCmqwV7qWRnMwkJtCy0ffAquLVaTyZ3vAo0mwp9eJk1IldUukl9MAjfrU5+OJsxZbuM
WeYyalYjdmFX90vhiamdqgHJ9TMS05VqI7XuBX8J95ttQgunIIaPnYJizt7SlcWhO1UYpmfhDqzA
FG0rpmHm9eIX0/qrB/fBwE24VdIOLc3qBHyswZcXhuMuYuciJL9zHvgRva5ZBWisrgt8hXmT2j7i
2fJbLN9ZF9sPzbaYXlT++NcwD9l26e0ec9khDkUDdaWqdS9Wp0QtbRFdubuYkd5YsOJoVVTABh3e
8tqT9C0DNHNrSR16UFJTJ7+DHKn8v0UQtzMppxU8fldVLfKk+wkgg3S+KlIjTBaWLtf578oO+QZQ
Xrgi9QVpzfZMfzL6kTE0Pr44z/+4OHrKyqgFoXLt4YEW+gA9BMgH/qP5mfOfout2JCFGizAXqxWt
CsuOS4vtAPHm8CaAeyTPhg58vUntq/Nt1rBoWQi2mDCen1RfJIo8wYFkg0Q/GV0Jen1uaj/qmUt+
dCZ/GixV9tSxl59EaYErvQYFdEH/mfr+o+smkyNBIKMc6fFkr+solCHU8VrYx3IEnieVox0/RKjE
C1kVGzRSiKXG9Unq5a0A4KV6yaX/nCIfzBD4df8NRbudJUQlj4BNdZo0eYI3dmUTnN/ECV8ufBJi
ZVh0oYC8RH8gPwNRpxfuzlgVkRIhL0SUo0LeAxXo9vyppErL4xHqHbmll8rmSkoEa/Ru5yRvPNdH
4YSuk5QYEV5DZZa77ANUdBKBhVh4tYjcRCHWfHRMvEpwi1vd2WhxwIuNEZI9xJHwpS6M3W960+Wk
sSSMJwUNUSCk+xlwm3DnFuf6tDtxCX9TTPNZq1/dvFRJEe8IrMZXnZFltEfzo0b/rXcPx8G0had/
/0JpbBQg7A+3wH1NSPSevf51iX5xGIi0+vFaELzSGrtvXEkTbjFqyp/VQ73nezzjqVGlVKMqAFhA
lxnn45G08PUHzbIievjHoDDXbFbHgt44ILTLtl6Luc+2Eh0OXjDcB8/3yHMaMBkRe2CNgtkB5eZk
0L9mFqM2xGXoZ95fIbXWKuG6WYovJPMKR04LQz346DBl1jtcbT4AakpAMccpYHEaRQu7lGgmOgWK
5D1zqWx/EOTGgOqwjvC+jcdrCTNYdvT9kdhgiOLAfk8a51v/1qeMPKM1KTDKrdwMFj5CfB5t9hUz
EpXOqKbvZ1q9Xr5x2cqFfOmovAs58h7J6IGQFpcdEuWg93PLZFTN8wI/eDikUAXRO7Zylu7MGo5G
8wp0gq5XX8rNh4ZPGe3tl56ytzPF9WS9x0L95X0yJMbHMg7YwOOV7mHXvo4vmzuT8rxwlQw80t/5
zjCOHmEVjgbwOu1f+XFCUD9n3Qf3gaU331a03k1TWakoBsyBLFIfcIhdf0MCsxVyywAItftFiPHt
UycFawrX6s+Thwb3ftgUIzLddK8iWPVSQpvXzfhB4VY7mnON0fct2/GmJH8rw1IIIpHlM6CKkE59
C/qE4OYlJG47NJNRbgwhNSmgAQlf2uwR1T39aoHrcPNrp+ILqappZgdevrwTKE4Qdb6KI51uI9iB
c++oTlUHDXWjMOiVumIpEN+v2Yp7VwRSUA+Ie67DRW6bh2Y2z6AwPNWxgRm4Js+uoykKlVnbwm1/
Zeus6NjWSISRgn/g8CEhMJfcl9QNsnvOy/xCDm6CDX6BAMmD+WXBcQ7ZNv2p5rKRCubUM3sFEd/D
SPA/0LQ34ZhLwE26CM/j4C2halVXkTm4viedF5l6l30p8uRodEdHFmHKiKSQf6O3Yc5piJr+D972
1Dae8/oay+qO3S5b0/+0+F9SEFwdqlXRQAO5n4XIo5dqy1Gz69sk6TOrL4bR8oM8rImJJSjsDoY8
6tHLcx+XxjtI35sjdDuuQAcEfEBl2GNYWBdfSOjti4TU1r1DoEtTvVR32scYjfuMZMrsp72pKTP5
8dGtxhnvusUugAT9OfoBlw4/Le4b1i+VR2oS9PcXvSDd4QdeJDB2juGBRLWxKLH7UL/Uc7Hqi5pW
R7jbrvIKf+rzCXl+B1Egzt9a9c0xRE/zsosc4czCCSS9taXSrxCwWVo2enp2+ABh/HWtShwkDPaH
aVieJX2Cyw1P1PvIM/+anfeisSd11wup3PLRj+scZBMDtJZ/6n2keBleuySuS9xJH3PJ8v0oMgcU
x3uISTlKH3s8oupFmZkvgbyD56AMmSy3YzgSeJpkzR58K+ppU3OeK0+eKMAMP06T9XhBRU+CzAeQ
aRrWkU2M4LgIEL6VarCEeyVTALhtZpXqCOgGi/b2micNYX0cKPQxeQRrE2t7IBkzcKPRKiAn8UOo
wY7zNBQJm4fj1JMgXEIUo5wMK0mCqnclvHBGgQZ1xIfViJgTLkq5wef6fIDyMoY3b6Ws0M/LCsQE
FjX+WEd2YW5fSJZLmFQ5ilqC0D1dh5kyLPjFqiWCGVxGSnETyxZT2VrJe3m4zW2BnfRXl7cOsanc
5aAk0M0fY0UT0PadcT6z3P4Bb8yledjiQS5yhzYjq03HZadfIgvQCG6pg2UZDoZcnr6hdKKNwY9t
wKKKzoRHTsIHyPbCx/MoZ/qib9bWq/4wXL58+BYNbfF9OohaJ4mLqFlEQamWRbH2O1aX7eSBwMjK
1dFGOcSzo6CqQOEafCjsFPAzAQ4clQCP2S3IEn8j3VUqx0J27pxkvbYBL49j7d5u4w+Jw4g8C0O1
N1ldjQuS/vFdjp2kH2Z+J5kdOyX38+gQ2kU66qLdkYxfUxxmmc1uL1i7yqoYqRoVsdJ16J4Y4TRB
EMoveiG59CY58maZYslVvO3/eOkSJyudbOB/0QUZ4zVfQJoulA8HjajCImFjREo07iNT/+WK2myJ
UP2+9Yfmsa0lJ+hkYvmZG1ZdpiT5UhrZHd72pXsZmYU576bYkUyxLMzaCRejk6uT8JMbTWzyD381
jSAPUjH6IzNqiZ3VxEP22XmNXk7I4t8TAUxXg+hMR8+inLmNy9U3RU22xnnD2nUV7RReCo8h4/J0
CMDnM5zbOcR2aMgZg5B81lNnzw1pW+s6iS+V0MYdT3TbQm6yddsymNdH53KfzMGIUCJo6b9lwGPH
i/ekwShqzUchIoIWt4pNKbTlnLxAZBcbgF3oOGQu1655GXYzS5rfW+loTIrtAe7Ug2I32DSSvmyB
XwkxVhSy+220ISMd2+2HvJo7m/C0PINwECNlH6C4GYLlC/1dUdQNeig9k23uki+s/yGiQb9Uf9I2
GK4Bq2G+mZ3ONLpNAbA8OoDxOJnKfFACNYxX+/N41wvSL9qEnVIq2xhB0eYo/BZup2HaGUrlQ7M2
R36bY60AHOit1WcXpdISLKVdiqBJvOGEzx3zDp1Cr3JptxkYJ9xFzJAghecJCysZzO996B+BTkZO
CzV4zTDAXH4B0QsSgzpIY14no7Y+i/r3R8Vw+Dz7sdgV9wS4rW/WlxJV1fZ6cCTe7Fbi0XqPArYp
zRcNFTcnKq/FtwB/tIbfci72ai9pTKE5+/SRtON6W1ss3ergYFnKF/Zto5GJF6SuePL9yVQ/O/WP
6HfHcJAyES/vWVczd8pHzgLEl2mD/AGtHpkDRi9ATcudt4fDm+ZS8Ku2XRoVLEw8cFlbukjeVmD1
Syl2g6Du1lCNuZAXPJXDEKuZKQTaeGNrf1Vm8wU8/KC/f/1lMVSL1I0NMokCumc1LrhJurEf5KZF
ZFOTSPgnkoPa0i1oAuqV0rRx8VEOwPvRE4m9H2ekF7CoJU8iRpK9PyyYzGTxcDKyZxQel10AH1jK
xpV3O2qS/qpSwCWmNM8JEv3HbmVkDkEYSvo/WiCllqHsKtvBRMo+vS7aWQKcox9+HDrInpWD+tXb
mRUIReXnV4pcUQMhMNGJ1W983TK3ejcdLFskNW8Be15uBGwDaDrvVjfyDBhnD3miiIXyAJBzdtmn
qOwa6mPZqBjCbaKt4w40Yzu/dA8BQ7S529C/hLdHxbun2Kkr9jtFu25ChmbnOSOQ/o4LKf7V0APq
XMW4wd3/u1u3P9+PxGVfeBxFVl6NmxKy76ephbkGbbHoUy4HSgLXiRh9uZ5wG+N12A2Dpz9Bz/VZ
pkwxubZsFv+/KN00dWwcqyaOk32pM0X4xuLg4TFsMC7k4L8wwPbx1C3qs2FJelddXWw+pSJ2pZc6
dJ9O79o3G2+tkUlc/5dhNreZyQhpGtlRbYLS68INaeRFWEWLbTUK97UN5E0wvEO7B4KioSLmfnp5
/tfhEwE4Kuh6Zf4ZHlb1XOnGJE/osb50dqz2cXCmqCEZ4Qn5NsFWWX1npLoZ/LSh7cSFm8MMLyze
R1IFRAkFScE4d6uV6KygRu15LG9IbCJyBjg/U7+9MhShb+g7aSwgwct6on0KH9v7R+3XDYEylVUM
TwC0Ym7ZDtaSGavb1av89iYjkW6P5T9noyyKzozUInJc6dB9X6HtDCSU4k68WSlhrDGKOoU1lNHW
oNgE5QbcNax00pI8oA4KiTQT2EPBR7Ji1Mn/kq51+e0LBYZAXkgUkZynsDTINBb9EB32UWOEIFU1
5QF6Yw2yVWo1lvyHLN3/alAyCvRS48QwWBgIRA8AStXVJnyM6KGIsC3kZJm/m4JqykWx5pIjg20b
RS8SKVXe23ZRtRBvKWDj9Z7ff7s52mqFAjYA7/Sx5L3TiJ0bwYgp6by+/HbUzQ/ImeRpeXeuG9Yc
BxU4MEP2DPi8hb6IoxGDHPBB1EhJ+Fbgz7hfVrjAPXrO6w9qR2QHz2QIMk9srOsfE1LFzPwbPP13
IDPzx0t0HTohgnoR4/IWIpfNFyQZ7fOSvolesTgF2xUc/uBueLF+Ie1XWCwyddx553QTJbl/SW03
yjcBHW9wG37ob6puqYEl74wuDcqIhzmO7m/GViCzSZ5bHTQCT0uHEAWJB/pIC5HIQ2c2FYJh9NP9
6ZLAQJf7mnWFbbEcP7PJ4wxyoIsu1awEDCkxmQbdFiZ74jELJbWBBCnC1u5y3PiD6uhcfYTxL6r5
XxtsSTYcL6Psy6p+5nFMei89bg4bwE3wmnVavRd/samcbzJpM8ADG4dX323h/AotS5+6+bRsaHlI
oqMeZQPc3zoFnHyMju2vYBfmo+EZC83qQiO0M0f4DzZ1/be6EFWQnRvAZxZ277MzH6xYNTkY/8/8
zTdkSjuR8UzsOJZpV5eoggcIiY26Qr+gnHkGowI3ARgHJ6i0ZnI3Xv5UHpv9hxxABH+XaFMAucao
onfVdK0PP7y8p8o7mBQmx2AFPAoF2a8idmhq+MNN/3M9M11mDKvWYgh62NWJZ9Q2xziDvYKRwQQZ
6Sn2+PVIEduTqGpOXrAyvGujLCDigQZDM27nOYGZJFKj0xn4zBLgfYt5jMQo4mh9C9C2D5n5RM1R
cyEmWD+W5bvaS1lHOVdj1l+AzjdSP3PbWYvSQos/7QmGPVW/ncs4bInohZ/+gBq4Gv9DVtyzJ1uA
gXH75ssDbN6HCCDaGcUFTG6kz37u8/Qp69CPtmVZO1WUJ6a+SWsKysyCv6SSfchyH7/Q+MQu4pbb
tOrpG/SSnqigvm5pc7vlxeSAAd98e/ZXxJWohPlB0ZB9NxILyl8PRs9sM+zb3F3o1746H20Qw874
ZSisjZSXppRrOl/nusrmQSs3UsLzJ7iZjVckEnNYu5k1uM5XgTvW2LPBuhkIwRq9Dl67MilTyanx
GRRpYpvf3pYa7ukOXuxcxrvPtaIhJMy0s5aosOPP1s6yXREs9etCGaQNzrePwr8F7S+soIK4IzhY
P9+WCowllvquk8KGhuGXzKKPpjfYG2BUtRBd3C0cSs7j5MJXJAJONMlFkStSGcENQVuKKXd0kiqp
cGQuewg3Pyt9FI9ApSDLZtn7pIE/cFnTLay6YrxUHqcttlPI258T2ZsRYSp+5a3uxFD11lDgk3lz
PbFG3I2xaF70lpmN3P9z/+4BNSnLeGWSmB2glNgFXgWlXc04VGhAL3umePOvPXdL5CUEWktxPpU8
sm8CtYiaoa2YAinpZGeuoqFaEPNfuf6JesOzv2HQfgLkZj7IOljIv5Fax3AExoDw94BbDcerWrx3
e+OCgu5Tn33s1QTuAtHkoZ5yvqhfA1KuE/s0Pd4++8n2BRVCh08BKK4nludDAuwGk6OkF2PtdTN+
PqQXgmteLINf50sI56+fbnLkfVNlX7q8yBHKnyXxVDfwlHMKDG4EclggNWdDg8PL/XJ9qRl0GD4i
4zQNJVx7qt0cH5qxsP8FMV/ZwqAu1OY/5xch5wG9UFXepLgMEPih7JH4oFziuWGpuWm9fEqlz6C7
vz7zh1Vs8//QV0Aj25FfxLmqvtuJphrqGqZGLTd1Sd83N0IhCuJExOQQzSOkd+B52S4feYeUebmn
P0kjjFyuFSMcWvNWkJ4XOA2OtjYngEHsJHtASmhAHtvh6agl8QTZyIIzAcKxsICewaI9UaPyI/nD
yFgJZY1yiHjX34Tk0ulxEGIvOEnmzjtm9a0fMuevxtkYtjl9G6tTSm3ldngEbFxG4VBnhoHkTivC
u9IJKFJCC2jR3NEFO+EaL4zU0zYKpvK4ghj9UaA9UpY+bqsuAg8VVUBch3gZd1QwrlYr5p1NDqRp
8IjB5ioImJBh7ecdPekKoT2Kzy9KHpBOZBu3Li0f41Q9G8W9mJ1/9jYGJd22zWLl04XS4mY84Z8q
aD3v+fK4U5vD1aXkn7AKurf0PdchuP30yWkNJ9fBDlRTBSGqUZv0AtapfGJMrRdZtDbDeIIdL+EU
vG+kJyGTnbh0Ozl6h9zIJFwiMh8h9EtnyB23XGi+qAgeHSm2/SZ4aFufDE7p6JtiIiq73DGrPVNt
XVg/TJMONCkql+eLYJJku1OTMJpDprOX5l7jq2L6aWnovWACyFsjgT5RMbidMKko/b+fahXhpHce
NyljwWJWjdv1DkjJB2meGhRhz1i06AQRgXuKojvx9ZTYcIPonQrfPZt6/kHts9tcEgeewcBV8uvb
jlsYVKqJLM8VxpmXw81AGO0tUiuXP6ISZwLqLF7ZvQGcZ1DL6Jo1WIZduzcOQNiUBeUEEqAB8Su/
wrIprDRlT2S4UenPr/HAx2b1asuyAI7VCu582Bw6jlLQ9RLJd/yJHWB2gaASIdUozcH5KY51FM87
lQAatP7lIcfYeW3N/6MVZ9cVtI4oJXEgM+8xP2fjUrQzwLwmQechobWRESkY2iV4Zf44Y8hQiFHp
ibRPjiUBsGaBx8XQx/q4CJJLyiopz6j/gAhC0gY23ZCJn46Md8QZmTHxrvVMEt893274AA5FIuRE
QhB7KCiJbl6B+6RSkW9ww0ZxqoXRf0BnyIhUy5oXXA/ptxZjWWU6fq0woJg6fDddxdK7BwztQL2s
4x+iso6zxY815e4t8jhI7Bgc9D6bo6phWdt5ZhuqqO/dfZHFdXHEWYQV4jcxhXdgGSJ6ZcM2xDR8
vdoEaV7fl78LWttIqlDPQ/kjuB9FXUl34xxVVP8uO8QIyRJbUXPKBoFlIXTCgu7qw8pq/dkvXPeU
Kk3o1MI8HHryH49ZcGo+1RoUn1/gg2m4P+hVnlb7+xQECbPI3EonrGJ4Sr+5q4yjUBOGTSxpEXPy
p75rGwvsoDULOz5NHoGiNONJ+tVJnPwrBHVaxbTEZRWeDdaUInk3UnGlm63TKVNe1xx2+dzuoV7b
cDIeY/t/QnWR0eERgLmuPgwWVRjc0H+WYtrIuHLmBQq3o3Q+d3xYjB4pgvTPB3IM8hlxO9gqu2Is
K8pxY8aTfd46GNJUecAnwOtLW4P/KhMp/UABdvEY2UQPxAECUUCR5VCOHNUQ80OvRuKC+lNqONnx
V4K+h08rB3iGcCzjiCyH68eaNQLPOR6Sl3N16U5UFZq6nmbwgoWRdEO4CBe1exh5jfBVkgRP+Yjj
fET3AjGrFT2j0urMPXsbo29u9p8CaWi7pvPTPwxwwW6O6kPno/JNe1IXVMHMdNMeqNyhWAbddkAm
3noybN11ba3u93weAbAge9Y8v0scja6al3rMr8ox29BGwjxpIRiHbUWijt9OMnHb/vp1dHvahT/k
vMxqhgHXkeNGrQejQYNBJyFIA3uOK09Fiy51Qk+EH5ZKKBYNVB8+d683up8xus/kyPgErLWxQyBZ
FZdpuZJr44IETR+vMvQTMWlwBu2AVhF1uWyvvL23ikpNVvMP0CAi9kwUwhFJbf6AdECLRW9Dfz8k
C0pI0i7W7f2TDsz5OWiBegteJ+6HwazwqdBwIhMni4UMSutHFKHLrTpAkdnhuhkw/U2Up328o89h
2LqY2mPhuETUMaIJcAi4cOCgCJ9UlmOKjZbIiiGuiXobF56xgVm1njA02Uml7xxWycD/kHZvyFgp
LXCyST2i3qzZ3V9PhGtvDk1ld822QoiZkJkOUHtP6UURPNdq+6wsGnTSz+fQkMvdqsD7aYLQhF3Q
ScrCG3orHERB5YpDWY5eqhCqlCsQCEJbNP7Tvxyqnw3q0HV2DOIMIZo3UxsN1b/CYZhx6/VRFu4D
1TgQY7fEz4588ZELWwSjPdI10S+gTVVCpukulwwTpscn9noPPcGa/mtKt29JCYEHTNLJV/e6GKTm
UlNJfut1ZtqjQpO/fHttKxJsi5i710NpKSfV0NPNcx0MmKzbeeATl/d1ksczviAGGiAhrFVZZ0jy
EMrvmu7XlBuLtxrEHClwgt38J3prykuuWuSU4Pp0qUUNRdFSpRch0iXI+L7gTO9aPH5vgevbmjrn
zSpAgxJXg5tFbN64GZ0O9qRnn+1MvoCVpOo33QSqpj+ThpJl3LgsN4bm6BW4WPsy2ByDdvqwi/hs
bwdtZ9GfN0+Em3aY+4reemCSMN+p48qHvJW/0Qd6TW/SxrYh+5/AZr0kl6IIuraAD9qW5DPqt7Kv
JC3/N7VKOQClj5Cbdgpyib9XDg9lVDb9cUEai3TZbUBtvFj/abpIUtY5+ZCQTPv/yn+FNb8ypArC
XqrXzp4VuF5HufIqOD+U5uTdkoxkUGP3hg6LJ3+WoRbc6MwsFeStz5QFqEj22rNPpbWlIntyD4Ye
01kavmhfBT/Ofnzuz5dryklk6Xph96T2N06U2qFHIvrmC45OmzzF4U0DgJotTF9qtx/lSSkB8XH3
1A33rAvJT2ZSJog+NKeGpqWlTsFuPZ1ijtk8KuPqigd8Dxqq7olake4imTVMn/fvL/Qb1Mp/TQDw
2UBpuz0PpJ0mjLvLEI+KyReADZxvqkL2FGNSl07whJUgY0iZsa7HwxjBEDG801aapZieIMFAxXYk
laTSCrmn2U9MB6j1pVDpJe1cYD4qieX6SLZQeSJwYu5FwD6WK7McdBhpGLmyr9D/dPHzEfaTRRXK
5LN3vn8e52ULK87o2ePf9Xmt6PfGoz4KN4/WvTREQRaMrJOpf0vxGQV/fFaaIQfB7Qwth7U8I/Rn
FlGdgYwMNZhjxzMyIwW6VdGuYI8WT7a1vU4zu+48F0P8wFdTfBYZfAD0TIl6qLBnG+4ZCsTdH2Es
JXKf00mwQRU+/O1fY1MBQKjIdYomrWsF4vL4u04PbvhHt1/DijI78osb5PAG6H/zUJJO7Z02LRUh
znioTeGBMKcOqeC1P/rkL4KQnbqVDuNSbWpWqBCsXmIh6020lKGlcnSDb5TtPcUZ6e9WgkD18YqN
zJ+wtNUNhk4sK0u2XpR9u5W2xYYoCXWtMSPvi5WEx+RclN4KY5+GfwXBA1Al+TC45eil2X2E2gzw
PQJBe/6zVVpR7NtMBzlheKQJzJJPeR2GqhAVPibtt+ty1D6pty6qusRD2k8JdYjktyuYDRVfz91W
6McWrKtdSCE2HsrPFwKsleCeaRCORMGr8AQWx6xcEGPoUsjFPLjyeQzRaURzT+/nsgL9J+dg6/EB
hhQJ1IypleYRo6X9Rp/dTDChNXIJgfomPRl5BZCNaqgp4PhpsOqaztCXxENXBW8aLwCQl2ohmw+R
QrVMtZl0hJ5EDItt1HY5CigHv/jUBf5RE5GvPpC249ld4ZNssaxBnhWRnXb5pjCdcto3hKzZeQmO
rF9Q9nbIayMnXRvayugzp04sajFQDdoVhFBMOCvrWvb1Y8lT1x2EzR3S/kBx4sYsqACJfLELnHUC
7r2luo1Qpbf82Eh4woifGkAimWqPWRbyGMBqRWjAoDROuXa52BStyPUvxDjEO73wzFcOTPbNa+Ua
oUuFgzP/NTzaE5FiKI0/DtHqBe8iC9dOyCKCLlDl2xbeF0E36TOxq4OIlDhg7/KJZIYrTdQQucnd
uZbIKsoKX6oCmMhehQ8FBEe+RG0KYcipWI/FM4XDTPzqbO8BnnOFPH0jifK4JYS8UDZZQcpJkiTN
51BMwDxJkCOmo75NVo85OT0kGfFiZJk6hAOYaq3wkiF6EIwn7Cn99Q8TnPlaf/bMQpFZq0eL7uCM
hq77lshJRiCGkGid1oN3pTg/yJIKWbkiGBd2Wa49Pmn4HT2xxRrell0agMHIq3mzBRTq8W9HadAH
JE9Kf+WsKxAhghqGvr3OxUnN/at1VOnXDd1SnENSKqnn4ietm5pGfR1veUglNc6BQBQ8I7AuGY+7
picXcjFwBt6gPTmv/rHlUvrl3MAJEPe3LR6vCt+cOe6cxWswTKJ5RGC7u7t/0xMQHWP9gHjlaJdv
vbc9KPOjpO65ikpMN6RIPrmWqyN6eAgOYpYW8/la2lRiERYrZk94XA1zsZMla7SOCnclf3j/6BGT
DBHtexdN7FNuF/IPunbiulWTCXWG/5r01lqLmmm3mNV2CEoLivIdaohsTMtB6SeR3Ea9tM+a/C3z
Srm1oEFWIEFpPFSueT04izjXcyQujVYY/zxcWfOd73o+pGWjVHS9lTWugZCMULI7l48KSlPuoBIX
o12gYEX/gosmlWx/Ts9GA0JQ/Dyol1dJWSS/2uMFJwMxkwWYAWt7Mu7uxd9keUCeB9XdKzg9j+YA
IYN0RvHzCqQl8QLEQ6Bc5xX5RkrTpMEhaj3QjHufPYR2LwcjRQKINknFYoyI44A1o/B++RPDp9N/
oaFRtpLcyQcTQOxMQ5lPSB6PQnQV4p0ZCv9RQl3PyaY1QCqqZlZqJqcIksFdurvpnVOT6t5Hw6XO
WUieO3EkGjauuj/9iiOcVrF8VR6rsOw3crc4wwZFqjjSLq0t1+y01jb50/TrTg6I7VjXOZhbexfm
SLBwN1eIeEExu2EP5ZNgFWF6Aa9nJaL3szMeZcntOeBxsyCLvHuVBkgiAzrPbyeBxSEZMH/OhqBm
jv8MXNDBINOO8JiZDIS3yFFX30wB9watoVcKvcS7rSV+m7eS1l+4hRQl2zkw19Nlg2wsBnTOe/Xw
g1iDXe9mhbSr8OhAC1Q9Cq6CbM65Jm22aWRanmCrB6LmYqoAyJuAhay1r816GHvDBo7EecW6QSQB
Go0mcYMV0Qo2azwkP879q+V7S8BerxNuIX18/luZzAn/V/wdpQH28FBUs6molnOov3VrYYOomqve
IFYHPkVVZQI6Kxv01HIH9ydwAGxODC/Gi7dEoSX0aBDhTXtpG6UUb38BmvvppMDLH+Z5+539fNi9
chFSL3uHBxBIibzcHcj9hlt3Ja10ey+OJOQQRRnHWQENdl4P8jIyH+JUKWqphK3Z0vIXReaxPkto
/IfDzS4L3N8yWz6fNEkW1EwrGlsTiRY5330QxhGEbi7dlxHj3VwE1IJnm9pouJDB795y4CVj4P9H
6YhWWpUkWPlFW/mmTXtsMDsdEKDzktbIRKe/uskBv7BO9i+2yzdz/pXekB9CbksN5PeYKvudif6q
0ODVp3apWDwYluKbTGmoahmkc9/dJpwyWx7m/o7t216YLDv1S5Ted3NAtJYGyQjpCWGdM8C2JmCX
JXT2robUPkY4Ji+4ncorGSTO6FEj5gOlNTEGbAf3+Z/rzdPirJMTvZD6Wd10lxUTuw9I0Oy6hRUF
h0wSqer21+glj4yQCTXxomhBkrpKZF265/JP2UVs+jFfnAnVpa0KRpp/w7oA6AmprDAISKYLCp4J
QRNVtU8CKTDYF2z4Xxf3+NPvKKLEVHMNkmwlXiZUNI9iOWsU/qY0wqA04pXIJNjg0VOYutIyz6/b
jLj2UQnJWsiUAyNQicNbvsUFUdl5joQ25BDJP8oerPcyvjF++DfN08g2KvaFfBhhO21fjjhg5cQO
2ZSg2Nq//6JJl3d8G+8t2ySpVH/f6a72SxOi+Wp3LBjNR5nQbQYEV7V7+sv+YnuEI2IOF3IJTlwz
aSzMltaGh+8JiliLfgN7O5QRI34Gmtae3U8xbCEtCSzgw+jcc4jGsdLVVmrnka2V5YIB9MoDYfVY
1nIwVBC6TjTDXA+un+g3P7vHepARp1KUNb712+mO+NNeCpA9U2McGlQvYwSoV56vBV5gJoUVMdmo
ujXNO5PUDKhlCaLFa0FQPIjxBEaPkQAZiu/+3DhwcGiadTrUbfNHnFQQ1nLr+ZGrt7zOHBES+QBI
s2XJQWG0ZS8jVJuVV88sGHl5Cv+BjjPwXl4kfHsiTZo6AXHBY9fJyokujctyYgRsq5RVJZ/EVfCA
q8XnRfAztql/up9BTpaYo/4rQVpc5XkS61D28szCHLv14YM82yQiGHihyfI1/omshgNOqbpD5Huo
vpOs09RRAjGg6cL2q+UYaK9t5mtpWqVV+ewX0lSkX/qIigr6jYeMVEC4xBPAPgSSgOOKaSXr/OZW
mSQ1lg0p5Pou7Ir1BfSmlic70tfVD8DOyoZfr+8/jOnfpQ11tFi6G8Z9/p9mE+7U6ILU2JApu1o1
2sLYT6BOpr6KFrwgMunjIXNsltvlOhNCvyFmGxNhN5NSUmdEFbW5TaKJsX5Oc5i/SBtGJ5VxQdez
4FsRwjVZ67X7J9M4VKGaGxXGHW3JeSTc/GgCsHQT7kDyTSiD9CPrgdiMojb3jIfCHhmADrO4m/GX
hjkruvBSnPDBKXzZpYLpQ8Gq70guT2aG+36GKFvWnSpyJw/0EqwL5UsddIlaNhIBrPc=
`protect end_protected
