`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZSnYNuWNSDFBUV7PdNQKzuqqVOd9MOcBFLY2C1DW8vFM5VOV/rgrzxMRdN8KfJjnLf1NE3ik1DY3
Am62El05+A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OuOJDKjBWRbReIaicI0eAK8ZSCoGB0N+jFyCYWPMHNg6wTaij5IEKvSuqyOjVXcAP8o+2QioiuXI
e65Hn6DSKS/cF2+iV4qm+fXmYs9440yCMb5eJxcr/kQJhUB0+5qhVwQ4qQXSv5ch4MietC/vlatq
gM/KDAwO+faxBj8WPLY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PuSR+rK68YXKTaVPZ38FM0nsnWn+tTm69tB8WsFJ9DG8c0oWlTrK2TghGNtxZzz8YEmT/SDfe546
p/W8S1YSJTxH3CgT6Vf6KNS7yyqwL7PujKb7HFXrC9tBcYaCtniPfNXpG1LAR8ULQ3WqouESbF0V
80/8uO1zJsFk8HcTRAEeH63tO0BBdpyu4ApSwixHKr9sAdIjUbsKIX2IGuPsg3gg8Nm2LQT3MYmD
zNCeOyYxLw7T306vZP5rrLyhKEf54y1K7APlwT52oFGkTQTnh4Z3Gr6boFK2JMNugVkxc8MXfbcr
jXEwT9J73ZZ6MO6DPAST7/FIfOHqiQzLGVchig==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sFU3RvToAxDNZKcpbE7cKq10BzIiHQNeyGnMu7YaXhMAC88i+T85nefjd3YfhiTL3fPON11uttNB
v9lL+dIduu8nJMv9tCK3+Dr5FXxjPPJABPBjUdPPvZ5J4Spm/hdxOGE6RC7XE/OENPonA6yc8HX/
P5HpqA5qc+9IEMFDWew=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TJ/CK4BPPuZfICnjkSogIt4hdnB6btFldZVZnb8KH+mysoBHs6eNHNgrY6/D+XJw824P45JeUx5r
T2SnUVvU20i7ciw9YIf2WDjDCSaVl0o9uH3rzfFNb1/UUK4jz7MM2DgVsnnAr754z3S96Ad5xUCm
ka51AgIdoGLZYWWV5RyaIgoVv8d3OfydX7+0EKevOlJIAVb5HJLOWkHpZNA/Vk2Wv+DhkzmJtGIA
X7Xg9hfN837g+JKHlx8jQZrMq+q4e2VPSgQJhukHI2n5gH3bEHWalH1Ir6Jxckxi2mb7w+2nuKYl
hTkBHhLZKyRp1W/jcsA6NSOZ/AA9E4e1x0RR5g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18240)
`protect data_block
dOVYarHKI/Ve1f8SwwS6PpM/wn5yivcPR6cLDkdptPbVLFrc9VXKvt8BWx9qotXKyhJq230lvnOp
dF6juXA9yp2kKWTZcca2EQvGbaesYVc06p8nOZSrN7ddvRKNtklhxdI4tlXWZ1/dC7UZs3dH3Tk8
/7dwkzgtYwfA31r0G2cZR2Sdfoi/LYtOOQKQw3t9PGG7RochWG/yY60bc/r+sKxSAmbgL+KzeWAH
eurqBlU/syEJ+0ju8pRlfv2r98J2UaYndGNPgkYSzMw/w9CxpDrJYy1HQsRfAdjwP9ol8FtPfX/g
omS6PwagEiAIZRQY9H9lfp6Xg/Bks5XmXt5vmof0QzDG3wVncnq+7kr9oEXNJXxZTF+T7IZHQFfb
EGnxaJtjWM4KUsYaFYkak4R8OHumEBwpoyVgKqTCbyYvUSZrq/FzWcRpcNHZ/0lyakzFrhQZJi/k
wpf4Dit97XW11ROP4V1npWHR0RYhFp0olM04fB+6DrbbLrstCfrViXYeqTIsu3+KRns2EPt1Vt3q
W1Yrjfv89/f8WMgysNQOeswBSChjLjo+sfKGhqexGXhKukJby+KyJX44cAx51Vdl0q+wnm3deQLU
c+kvRVF4yoDd4VSb0GcBGHTKHFnz0N4DXPX65MvQxydMhYWI2c8jVWBjTFe4arei/eTYmwZJya+Z
nbXiuRaZIUXJIkVvhw5dCVeshFbV4+f6GYO/wEDqD7hE0bJKHcREd5sxNfnTIkQOT+yXE9cGGf/0
9w4QBr6e9tWOERGVcspHtPVXEr5PYaWdNVkxPSiSOQyoJNRjjcuB6zGW9J20sUqUqkaO2W7xiH8Q
M71SfYstSPK4Xn6dyA3sJGx6IgEzb5F2cgz2P5SuPOErtUTcw+R/OUbCHzz4v6GLeR2BXpy84591
GSerqXvQ7E9fyTsOoPsQ2bzpcJ8E4nFnozSuU1KF9+oui4yqNWLCNvY4Mixh0UVwaPYH3qgKoAcz
UobdX7qLL9sUjB0D0B3LCTjHarzLB3eJlX6RtfZgA0xJ4yfu/4WETHMmVk1KnUpUGLgXrs7LKh1g
pIsihMyd4FXI/TFD0YKjri74eRv1p7VRvM5cqxiThLLxIw7QWXm7LZJUA6ttK040WC07gujM+2MR
H+vMVyNRJXC3yt/DIr9AuqPkOmUTsSjsHEhTm3SUGCl0n2Ky/9GFVEINH3UV2nqohP3+OHvXyjRL
C9rAQE9W3+kOAYdxPL0xVgQ6ky1X9gLAXT7TxLdfMxLnZmmkeTE7hMczaOxxgBYEki1qHXYQMaM3
lw14lGM+CIaIZzqO4EtmwBqHBw/YhlxNcxVH6SXN844CEQgNTV8zOMCfVunpowmdq0e/WL0Jebge
KLqyErXfausWfctVSmQWWeOiHsonGXH6M1TLQArkjIzT4gL03+eaKjYQp6mdnHKwbcD9aK80XQeu
lhoHve7G2EQVYSigrhdrAonsVUUKLCUyIEd69++DQoo+OZgFo9bklxf68AyEenDbUfGuwOBTRB3S
4IZSsoLuZ83Eh44JLQhl0TjooqPGkRtqaLobcla3YehKneZH4bUDwdKtrRQ8c0JXBnbOORLJjH5b
7uSC2JWGIF+lvJb7LX9zk2+E8Z70og8TN6MNO52Il37+2pSG6xU8qByaD9rW0bpHqHoAgdH3VlU/
y6kKyJGyW4tNwUJzQEW6QVn0Qr0Hjoxndka/kToWvD4TtxWm4B4txUnwMVcv1pgxfL8zz+C0Pppd
szZrIZj6OOP6d2FmD3/FqR9gwqwru1/p6sn/bKJqQG3aCstaZzKrcu8jjqSBUvVKEK3j26Eso65j
rN3MEwWDc/88aL4AXWIkIROLlA1ZSzEEGe1jyJj/O+DjGf+K0EPW6ERRTcbndE/vrESqAnJQ3jTe
M+zd/gtLVxJRoBLcfxOEd01EusEhFpGf0btMnE3VLkL1aq8FkpP4+ArcLXyo5n5R/obG4Ftlk2oN
TSvwsa1s2yfqitbqYk9ABGa9ceqrkXWfhLno08HtyIqnQLypvM5AQWDy6Q4VXBu1z2F7zBxTOtrT
XHVfRR4utDjfuat8zHi423ZceLzvzj7eAKs8xwiWPzVLxCwHDMviJBXsrG2gLMolYm8xBBXi8UqN
oE53FzqvcIl/Bs/yGE/QNDaV0m2011evKvR848FNzgzflqqGCEil1ajvQEF76oGdnQ8DbgrmVBdu
iZ+JI1DdlQtttdZ4BmcarbthJJM+kyqzfePH96DVdKDZ01JL9YacgS/Ba3mJNHKjjaqERJhyUkbd
qCQrmUcstFN2/v87KVOFWiTohf+hseGe0ddZq/OkUw3wjQ04taRpBPuWd4qyM8Wx8Tb6LLtWGALo
M68pu9SfCnakDN/CL3sqPg2GMb7lmpBFDadnJS4jcOoTlIWk59GsgelJUZsieS3cTmRqnYl9YMiD
F3tBMWQtAsCBh6tr00rqNudJjYLi0kJQTUW9+QCcmcv7QpAREiRZopDcVITSbCe0j5mXGnrLfsMu
u5L5vFFp9sxHnswZejaRcKXozuOvl3VJk0NXD3vuxvb/9M/doQet8nXz+O0gL4My7ysPUSSlBxKK
uvZ5Wsbys28v4m74W6s6NgE0E278eP0G1vYXfOZpJXZEqWEYUXTNVSkJr2m8gv7/Oeb9ndpbG5PP
j3j9j8lame2kxCB7l88hXmO2Ax9RSo2NaWCka8VrHsTVDQpjRMYwuX2ahxO+WeqlvGb3lReQlkDL
UO5NyZYOxlEtlBloEDlH7jmWyN7Wg1zMbZmnrd4virTfs8ACSKG3uu6vRUhg3CXCyWgtJfw4lx6L
wGfMXFCglvYrdl4dNrxiiDx9FPDAkF0R1w8ydiZ8Sn/LRkC5tPxlN9cks2fYIJ0RzdnPZ3IajUds
C3lH+GZPrmZKgs0tx5Jg1QKTqZjUANTVHuKW83qq9nxACVofcz/uYaWKxLFGYv20DAc/WyvzPEzP
f/zbLsAwhvH5+9ZvMzJrIM0rVV8FaUcyQ0aAUqXq/ayWI2Bv6XCVKrpjIi3gSnZRcZ0xOZl0B9TW
nk8ASxk7lWA3YCi15D6nUNg11yvR4iNS3O57EIPlCYm1Jc5FeB50Tz5+p/UGcKGU52Mf/JdwB4h1
OYqde2a+GVx8HrXw4gMhx8lTlPVtuHh6VWAI7/GjQ/6MGogvedTYaaszOG9vNhpbY9CfZ6mL8MPy
zs63Y0xWF/V4Vwbbb3ljHz4nuK15u5Vd6vrvBfU5wJ23JgGbzTTExgXylhRfXcfIo5iUQe4VMfot
sJx86rfb3KJffe0LTFXTxeE6QeoecZRf4uh9TdtYsKBg49N1Cr3v/bwE8/p3YqFt2SLBFC2D8qZe
wDMVLU8jQeT49JYJRvg5PVnrRQND+vkx4TZUa/JCz4ApA3+sArNVlS+L4U1ojcC4lVQy9W5lYG67
7SjvpCsu8PUBsYAjiXYd+kyJa7bE9ITJ3kc7r8X43wDl8e5+RuT3LhOHUp2AttF0InsTSX17tIB1
XkJCdz5kMcCrMeJmauXF6yBIx18VEE42Wekwu9gJ+rxQt6aeouiIBygXZCvDV3EP3qSHck8RjILK
IE8/U3crkwCB3UMImk5LNbXTlCZcqXYWYYcJUvJLMsi+DPn+AMCun15KBnsa4PYAz2pBe9ojBN8J
/NLPm1gl677bFzwkx15sk0wrmLP2TuFkH9m9INdvEjwws5+xUELQWBVvso9c3fFuAdr1d8g/tMGU
4lxRoJ+5hAt1Psfaegfkn2JFrxijW4O/QprhbZmJA5W7T/Hiss5Twj2jthtxanIz22X6jJSzwqtA
P9sFGMajlIW3gfmzgrYB3Sf7YgZ/aTw4zwlS9grzB9rJJAabM4O1W2IsudKIb2oxtYrPZ6j+bA1j
ZwDpuH/lWxFGOAmJlmhM2dnPTj0pz3PpdhacZPD7f73WDaYaxwJprNi0EIneh+2kq27deJQKXtIq
7u9P++XrLXoYJJKSRWpkSBv2Geeq4NcunpyrIOWuojhdzYzdfRdNWAxBxDgzXiMGrMmVpNMTvDDP
r6Q1r5vfn2pPG7OC5c4KdgAtNmbvPdsmur7uSUOJTzzIy90PSNhpdk9dROkFEhU1jcYaQ20dTrLX
bhQoMC1GfiU+VEfVumQZFM8Ylvla8FUo9GZk/tc7HqXvxTP/ZVQ8EtCWf7gA0OUEZvXH6Fws5voq
hc+j8rExpsqD+OsgMGLNdi8ZlxrGwzF4sNo9EzcvZMNd3mXjZB8OZ107q9bEngDEbdya78oxMH85
+BELnRDp1WD98YJOyiJRrPse/00vs5qNsa/TrlEH4A4a5aPmxMHRNMtaTypId2VHVUrg5CkJR7eX
os2nvolGRP+E3ngb/fWN2njGGLaTamZP3PH41JbCr5jMp6OofDY+boRNMUOobqUlFPdvfi+gGzdq
csQvFZyx8hosn8lu5SuK3ycqQB/45ySYpzYuNQBcMrlGQvcHpvssqbGzBxMgGybvJ9nLnVP8Pi91
R7YAYibkHkDHzkAwTcG3GGckVioryA+vu/Q5CpJDsWaLR/Bu3z/8TC+edsYyXKoxbkrmxPSKo+sJ
VBfLcCZo0Vn+f0OEvQ08sOMRJ1EORI23E+a9w9t1tUTfnQ44H61dsX6Bu4fpE3h5/7ofgn8BFdb9
DWyGIU5iBOgG9ACbrX/HlH5WwukC1T8oSnqTlQlGbUBYgv3gL8+3+R7jf4bl1i4lMbqKyeTDuF9l
GHX9f60V9hRx1l6E0Vdsbw1kQye7WrpyaeBweN+zhnuKJcNfgFqUqNjL33FavHPAzZon0WTJ4d8K
ou9IdYRcOXpl8XN6Cd5xwmQMAU7FybFYCYtv83mnJSscaXO/LrvdmH/IxJnQlFKZJos9en4MVqep
q6R3DEb3OomdOACxiaWXHAM4ZRf/4k8EbMr8wTxV2W5lf7FwoSxSk9UG072+TTAVMRtEHUCOhKsy
63+CjjBntnTV/uqGBqzuL+cynBDW5nXalllsg0hojBaUEZ8sy9xkhjwvhh5Wvkte5NnoEoOqswOY
X8mjU9hHrKKB24nC3Phmgj2f2o9qDl1iAC+sJpfI9w4w4nRmyPPDvCN31U9+SZ1Kht6hEaqVdSDv
ZIIaOdq6TtNZ65vUdND+9lTsrivAJk2RNjR/yR8VQJwsrXm6c66reK0YzY2KSAaD8Rprn2mFjkES
PEJFXF285As86zoqtuEYLSr/JkYli8prKXogBcqZYe/QcmDLpyyfkb+qx7kE0UfPZzZDkVRKMjET
JuzVCJ7JGZKsIZVISf42js9cfhLzgvIAuiNiiW9WPC26G47vH7GCgqnHbHI713bBZaz+/YoLK5nY
ADkTTuiMHyALTJHypLnuG8uVCFIsR91tl48n9y4+DbR7CSgLnv1Ryh+aSCkPBDDYUBG9663s6Ziq
HxQPpbhFp2hD4eTVSJ26WVI6PgPBnq0zcDnGI1intzGm8jNm0CoelnwNa9B1iERk2zZtfPju/BI8
/II9XoTMz38fP5DONYvdHSW+/EuGA50MpHS5ZoGjih5mWKRx+2P60A4QL/XnYj0cG+rQ8t+arbdr
epNva5rYBhp1KtzTjLG1yRVg00AFT16L/WpGw17QbPGePYni6SUBVVtDYWqlj+zP9DH+E+r1sxci
tvU896AbcJ2GaAM1WhaEeZOvMV187fevFnCHA0hZc6BXznAJTAG9QKxTI9/gNR8Wbh4FX5VxmbiG
FUIWO+IkznZ2vCpTA+wSqQpyQa5tvEuVcOh6Ih2CbACLq4RPacm/908TKzwyCOw57DKopPPLyRok
Iv5Uf/XsZArP+A0w0nUXJTOytbWrU/g5vALTo7H2XoYd4f41d7t0KAeg3Lb+CWM4AtZNB4b33yG7
h95TkqAFPHMN/oBvDHqfqvE0akqy+j8zT1NuGvemI6s495rPE/gdYAFC0od+rAzOjhLXVMbWDPyI
3vz/KZQ3j15nqGn/CeYN8wMl5s//93xO+P0UWDWC8vYGpYUqkn8GrEcg62DKO6qo6jq3DiIpUjih
U/8W54gtkFGIXtrwh2YDUV86+NFV2KO30h55HkFsYHREs0S5rYRB6Fh39b5qCjnLyutgU7al+PQc
QUjcODCzMv7PM3/R3e//ZayN+LlMe0mtYuSv+rUbFX2yd9sG5DCiGrl0NpY4um9PD/lIq+TRlJ7I
BpOudY8N1F32kO3jIBHTZFafe5Po9I8Bua+lQ49t4elCv0paZHEo4uPBp5xhOt/rypfDTLhtpIxn
rafD6nnczSUf840GY2MFgNbz6mocaQhRcziDKO1Ffy2VCmvYDgROxXv4reorPMUewT9rFAPXxct5
G6Qu9fiBxmLnPrq/VgwhKheupZiD3qAmOizzZU0Wo00J4J/ofeLk/6fPFjGNViZfBHta1gGofJMD
m9pwuMHNnL89lVrYublFyec6gtrsNRDUFdVwuB3lCLXHATT70UO+fE/inwl4uHvHkR+/OZYkroXw
Ns9pUrx/pn4TdVYGpvdqYJID6evmHkeZMCS7SjzXHhQs+rvjNHLTAtbqtsLClTZGjcIR2cZOPsFt
z4PwCVA4Tw4o+bQ+MZfdNEeqDITXT7csnopFPIqjd8NrN2jx+1lhhMzDJyFmMDefwNnPpBneF2Sa
XJMhJPCZUJ2tvp4DBqPWSmFrrZWq/I1nBGS8XKubWuneRPKpW7heKGfLznknztxu76OVClcgJFrH
f2Fd2VGkm5NEENTK/usIaKg6Jj8daGQCVhhC7n3Z1+veKxK3+wLJKqnurVFREJ6LljqhRbn0yaWI
AEZ+kZF2hO3m+L2AIs7kPv0b2vJciSpa593osu7jyR8XLQaEi2QzzV3BACZ0zBnIwEWoO3gVzWD2
ksqFWQjytY5NmO5a6lW/UchAJ5yZf2oz4pxl66hVxg37b4Y8gBP4VB/JKVbB2jJv5y4GKOZWYx6W
wUrsQjRzVWsCy+FIL85glHBsjN+43x7qwRn14cKmP9IgM9wz2CrjzehtTjByF16VDr1LU9moLaOx
14o7EQZzFK/qnGoyx5/1HdTMaIwMiiJwZD1FBjQdebDXK2O1dOQV/slFjN9i0C9WBGMeh2DQ2iqm
bHtQuTxr2B+oEJn5E0gSZNiOGO0KFRjbWEVdO66sYAjQe2e++BDXCgslAlqAB3NV0AjlrAd70NjI
r1IDn7zFIcCpNXs3+fWoPWOOOicx1fmQt329lSUsahmB9ufzBMoKNCWcimm764cz6kYb7zVKkReV
4iYwYyEs4RNK7uveqJbzoN8kBQmoxfcfJUKtwYHPxRtMznIm+mrC1CakUmQB+oJwY9IEvbZyJls9
Bgp4eYbDVsvLVE3gYjcu7U3twFxki2+d4IysToHHNtAeT/vbWWDdZZ86NU/5nnaqdt2DXnmmsH4/
YvkNnC2TX6gsof6UgtuJ7kUQj1iUkKXVCyF3CE9WgUAefpaPjB5ZJr8u3lc0xxq228Kap68/fcDb
NFD47PCMCGm7QLoY+NcIUKwD5O9k0Serx7mx0BTc1VArR2OXNHm7V9OZjsKsBTNPfqsNi99ded9E
Im4kMi2qoP/hT2F1213QSvVduPnp8q7dzGf/goIrzY8qgg2ZXCbl8W8oyEZCxZYCjryACAW6y1yQ
TS5+lmno3rQmzSQrfxA5+NRTKjH2m2Hc6GghAQhSEn7XgeAPaaYwcCiLug5aKuZsHMIz5pScOEwN
+23/1FEADtTLOU7v5zv0sJ4RIjkHKynEGHio0YD4ooiw7ahKRRNtSAsBHpEJtOa/zRt2JJQD94qp
UOxtTv+1nbUeFuenSfMxI6aznL2cn6/2qLjPPwi7vKmUaoXwyh0Nhi7f0rI9JepHpoR40IB32CbT
7YV25+4MGKMBinjO43e28VvOXCBMXjpV9K22Q/7a22s/7ldQjvMgQTXuFdXSKKpMobn6vh3KnEfg
A8BlPf4e4IKliWNb91n2NeEkNLtGVdtq5wjoXK6ExJZamQ9QgaWhXEvUEpwQXRWdOaHyUj3G8E4U
CxsWX6nW/E021f9T35frFAUKaXvVJZK6NBkEF3Wl7VXhWfQb8XgVBdJRrAuP8P58P+3111RwwEri
D0LDyE6t+h3hajkZ+Y38fMU+27q8XOe5PJ8NQv4gXjls2VJtMbhPRpU2CqPYOS3fruHFu8vjQSds
miDMK7+9oJeW7TAliphEkU3RqEHQa/1JYdWBYJj9tysmYKqf4YnzhSYGhkE9+xvkv1njO01mdyxL
rW/V9gBt07z0CfA7p5fEv2hE6ibkNyna/HDCU0tr5M080XD6xJyGumFSNWkbDYGCGieOjNXSHGI6
mxfT/kEKY5W7Ip5zSj1afFrxlSApgo7TTOjJIfRZrosxsOullf1X1Nco1gGxiLVNZBI+PG97e/bd
KDBZFS+cIrwHbAuxteEYriBN1qZu3noz0B3mjSHI3Almk+YKeW87ZMN8XNGr6DBifaNDJUOfPSBm
CDk94KF/PsJPErQfpo1ZEkj6Fohg6796/YNIX5bPOrO2c2pgXEycfWr7vh1oEZPx0e1I6TdusFmJ
RxNqkYx2orktFbulEqqv5NECzChMoEM+HCQa5+6rEyBtzcmKL1fIVVj2aazLOsGadiDhHRutCti5
BeUWIjLw41XDJpGWVRQ+D+faNWBIt/EGJMqoqLRLZoJpRe3fDbG4f0WgVc3ubSGaDy3QCFq31YPD
liURs5ez9x0BKUXIc94H8uaX6ASgWO5fPmBM+NABAHh6ew7SrmoSJE7/EARd4sedTDY84rYDvz54
9Do4M/5N48P+dtaBQFdh91tXGDKxg86mokZI5uVIOwsIJQjN9veyDUPOZEqjTfUU7Wl9dR5bCbik
4jfZh2Uggpv1WkklF2zhSS0cXMJTfTZuNmSTog9w7ZVOQokEoHeFhLQ/O1cltJ02ZwZjoBJ7Q26J
AKSaXQPoC8TYJq7yDju4+cpnMlXwdL+x1bHDH+4WoK0HLNwrlhry9i9ElCAKnuctUQvot3r7ImpU
lqEpW2r5ENuaVoUM+EopT5JKcnuZxNWCSPPnvyP/Wmj7qITGs3w2scsSJ/DkOSCzVbAprjMERD1i
aBtJ+woZViy8xGxIFjGdkH0aNC+FXZdl6b13GJpKJPOjaagjUUt8H+cGqFZn4We0PuMyglmCFuzW
D/Uwn6ojxy075ujnuWWlHr/1PoNzIxFodgNNyX9QO0VBiUkwm/TZXzrFRSbqQm3lB1q9o0ybZ5tj
MqR1Ac4HygOny1UUBfghQtFfdDRUlNSgH+gzBueLE+9JSe0FF4qbCLoANHlghdP1uHgrC9EqEV/B
OtxdECGBgnaGuUYnDQBWL9glRKs2YAJKy2RPTdr/UwnE/+dbkfq1QwvagIfLVOjFjTXn3ymoMunK
MYxsoUpsU9WPXPv+tLTlbMSriVMjq5oRU00IjRoim9C+e1WlwhbgRe2uXxwVFnnp1GoxqZj7QQ3w
27jCqWGBcgjBs47XbAVvPI1v0oLc8KMerArxfV8Ba9qFH2omX5kKczIZzvjeffeTR7cXnpeSAEd9
zejH0bP30LKu9aoRh+qSzgSz1F0IlpTNhZO1GRl009+3eCOSJcQXxC0dma3N04q+wNjWjasDRSlN
pz8CzRhe1el0mJwGGMs4ZPV5lh9EK3mp0kdujjJMSxX5EkBOUvzF5tDd+COmNDpcsZM5nelye3cD
t13OdxjWIiDU6AStvkEZTTAEFpibnnhiEBKaJMeg1xe4Brltoj4z/t6bt4Vim5AtwDyp7VxNV/l2
1ZIk2/YmATNL3WbB8JSK3L30ebrRu003YtFX5B0kt7ZGWsuv6l+ET501B/9/YMJgyhDyCCu0gjc+
ypiOAB/FhY1Nwh337pdjoq3byTemKz7aKghkuHWAM2VKqiZVyFAk5a4LfVmY9C6+fVOK0msV/AXT
uhveO4BJsO9EelA+9UQlZbFmmqP1JXndqbqGRr/NWP23TamWjfUBbfiiyhNzF5DiU1cROU1ro+4t
6AllMNqqOYrFmPKzRL9IXcdyeXRmhYuhGvUHgkHe5tpEC3nyErBbjkxfUxWKEg0y0B9apT7yD4FS
sEhFEH8AyeXHZsjX0RyBy/C0VxZ1yQkRSRELqpkHU4HSmsmAgZDM7KTb5MyEnbIl0K+BPwFOvEgz
Ml4o/ZDtuiHrRMzu8kgsKphH8R8guU0ZLsaRgLeQpBOl2X9B3Yw9nrnBZIRpzc7tMwImZ66149vB
th6en7BbfDycg9RrrV4uzIKRysLl3sZavMZVAn17tTyzBp6LyIs3PNdb63hJvVcbEyWAOr9KnBgI
0jb1lHzKKGaBz0rHRhvGdi5guX47dD/JTzBgDyK4bZA5Nyp6nzMTc5l74tvShHr+4EswqrO+9X2Z
ynwwu8Y7zQoGD43RLYuPXnH68KHSU2jy9U4uoFSRM3mQXoOBJZy8MMFrqykuxYwqB6Pr9dePrba1
RaZcIrr7xCt5ZvuIgAtJskR4j7LfiKs92tqmNDc/2OL/Fu9+qhMWVkl+pjIBUFCFbOORQfCL7vmX
ADCqEO20BV/bGS4Q3gz7VO6fmb6bp0L6Sz6tEW2Hbr6BvE2mrUdNvXlf1KokvKPpvpKZLBTpkKSS
uEIS6IrCKWcDT5ooqWYETd6PGCAUkImVdyl16iOorJXEWsBmmqS5xzbq/c/pRqntz0Akeb9CQhym
C7InNs4cRzEWuDScIq5/jkVXjpbIlgwIaa0YztFTRAEymLvfLx9X4jAG/KkD3Ubz9raQolE4/wF3
nh9up1317N/JRB2D1D1frXeHgvP4VGq/loK/AMdI4DMe1YABx08IX3cNwHhFpxmO/rpNGKwEm454
s832oMdiy9KbXKlUK4FCTvVI3kjCA04eQtOmrtL2oUp+jqSGUmU6gER2LkN7u83petBqoS2PpfWj
W3EeN2AXVEkOHCdMetDgMYv6iEWUxF+RJ4JHE3tq2EXwnury3tDTQZHadRBvyvzcGPwT7sxr/Mx4
1RrlyrPjcQ62sddO/eDuSQRu1r/RIvnSNoDdJ/2atUXbR/cjxR1c5ewH9pcVqRO3nCq9MjEonObo
oH5/vkpD+q0ZSpAPoggqadhAyukVcRRTUPqUn/gBn3lzUmxxX7psuV2U821b+6ux878Aexf5+HDg
qmBXQw6zcHtIU09mUoMgf41tHvw4bGSqKLjRoARAEGLdy8WLKvilkf3185DZzA3lZWcV7B0i9Yh8
X3UY80kL9p3b8wB/y0/Mlj28q1QfI8YbO7yOEGKt6jP8pLQgN15Gsl6o/FkISgWKQ7YUNKiGVt5S
eR4mBuYg0sjnUKT8zYXca9Dl/V0gTKJjAyDByMlxoQnvp+3ereM8WV8E0++fxbGBHeCcyQejdOBl
5hLTNH39HLuyp2sFE6Ekod8S9EVuO53yG8d5VUwN9N+g8cu4wXfdHngxoulyy1niZL3oW+Nf6qUk
hBCaLg5XmlrlmKgUknmbhTeWcSdAE+TTZUEnDuc6ZSrs7bvfiVDHTDg0h1m2i9g7San2iCYtmBcJ
wgrmtEvjb6GgIq3tl60whcC/GpYlRwOUpMIFYeUgQs+BJvY03zkD1Dro2lmgFOABo5atSOGgMMej
xLbmjuab0y6kHaAA3qzZ+tD2uJeWjmzgvGfwITMY1tWg00LNvFIX3sAee7MHcBxVw8rfKGLNDgXc
rvroFwBJaprPFmDiYp8PjSWFaB/AGs7iWeH7XS1/5gVpEE2HzFkiHmc+zEW8qZWbM4thdE3jC8UL
Y9p/ZkS7cLYmsLTtXlOHUlI08xbYeyJ/WhljW2VWHVjW97+1E/Vx3H5QCr/5cNMje5HMVzhRCvUe
2Qt5DPyWsnoGlzmtaX03jduXMmZv+cO66dBYojuNrPgcmv0Iy7se+P3abxFr5uv6uysqdMZWtw+m
IWrkRoQAttOx8BCE1tTI193/qmWLPYxeMuNsXygrZOyEyo//HA/WgFsh6I1Dw6eS0KgjITMUlVVp
+XiUFi8B1LxGpcTZrEKgeEoUNAKZYZwIr6DV47ioynoAX1jkrJv/Vme/ESEq3gKiAIq/wL/ayHjV
hiIQBEXZGdQBdGimbcVE/f8ln77xdoFf/ADzS5nRzvShzhHGNo2d5ymyauUpm3L25F2GXAiaeTUK
ht05OlYXIEXpVVmeLGweppyOFNkDOHxDWo3EyMMg2SWoiFxuAiTmjL5BB+R+Gi3rvNPyX7GbvhVS
l0in3/zIRO+NKDCVBzWf3PbD1Q89C+DBXuwylkzwZ491IIDrh6Xn9YzWvIUPldZnQvgYgHsBSvdX
252+oHmPIFEOvi89wey2X9ob63EXcJ/DlJF8YtC4oxZaBGMSuRBfOa5Yg8Ho+Aor+imTiyRkQbtX
i+st8IJj/SGoe2e2kM+hFYsj489owW7hrl15FrBsk4SdA172UjDI82CLLpunwJR0oxX3ZRxQNT/T
30MyyxHoevdfNK1WZLXjHF5HwOHKAxdIhlCg/mMv/AST/qm81dmnvENlevW+QWijiPdfb7ISuUOZ
tWWjZiKY92w693c1LBUdlIquK1Q4oU0G0Ft57RRq8BBcfMW/BvUK0Sv4GtvpRW3191wteq8ZunjH
s9H69tIABKYkCdeEvk0Fr/eVmGTbrU97gxeg6WaiIHFXDawoI1zsP3vij/WJjAXfrdKIeR3M1M5g
nt6Fk64VtcegVl/rqyzdo8mvQEPy1Ct8Dx7grzU4GRuXvQ+NOVp4e8CAFps7p9m75OvYYGxNfbVN
cYdH78uTZUJdpus9XOlUiyEGqNHJvpUKzAMj4UsTmD3pI1wibjF4EGhQ9TlNhOpUzTwXbOkkoiK2
LPhWeGm7VENuomqTfLBqR3zaLGJmN252fPHQV7MW8DXXw4GRVhiGGvFIU+YLufX4u3BzlUymP94E
l8+ec9Jl4tXiLlmGkhtwLatVHD+omuT0Mr8FfhV/6dPRv9DofoHks7KfiQw4gZHss1wi3WLc42U0
htlNH5AidkpMPstlOoa5rUIbOI8g8TCYK6JO517tZ3PeyyjTgfueSZOBnf6X2Kke5OxMaJpL1gxC
6vaC6k+v2SuyU5pIs6xuZ+qxPWNF1c+VXliUdNHQ8bODrpBX91oUUmyNu1ArnCE0lnciBDObHfL/
jP94tmxIVx6s9zgrk3ocdsni90xgFhj3P6+gu6ziV1VvWDuYUkf20/BsjoN/Rl07Q1F3BvRGyw7p
TYm8FPgocxHZQOSu92UWK6VaQdy49JC7ST2U+yTD7UnYZ8CjAZIGW0/2UtGsscS53eGZvkjmunEz
aGXgVFlPRuOMECQ0vi+iqGhm7mqF6Vqq7NeEB/8wQkYhpyB2+54/tiNG9VsECdDBiy76bG1qESgg
124Q834B/9db4yQ8h/cUUMlM0Z4CHPYE1G/vUVKc+uLYQD/TMmJ7NHMr6M5irzRef2fD/44nk+TJ
XTCGfDH8t29slBfmo+9mZV6W1fCsGVmTxqKghpctPPgHbWgUUvTgAVugg5s86I6/iSDkfqJi7ykc
IWvkXS4EshQ0yN/bAjP/iGUH+9IXROkIBZ/b7TybBCps0CYLgrRcOSS4C0iIN5+p3lYK9LtpCMmy
6GF4GWFxikr7it9a3NixCgA6tYD1wZ/VybVMmiOVci3ix6ivDwJKeAiPzqwJB2Q7agxfEMAo16kU
yaG1L83++bw7rOD/8aXLPO7cG2U17xp/7YM6WXXVuETkYrsPbmovgbUpElDSspVhSQ17rjgWXAEc
0El/9INWGpbzanDXQ1Dtq0xU7pewiO4kKmtnV9n+WtbiHj8+zTe0EZ+w0FVMUKMpg7uKfHIKZbKG
z8XZQZPpniM7TEOu7pbgfvSqNvQmP5MJk1edSfd8gOVhNic7qOFwImCCcC1G9N1slvoGaecijc0H
l6e1L6TFo9JJri6TqCJ+VCrN5P4AcoPfxdsECZGX9fW72DuwGjVODg7tZSkiJzazxgkaHaqA8OZN
ESg7x6Rjm2xvhHU/tX5YzuVYVMhyAS3WhRdl/JqslbHZxGgJeVUhUBhciiWEWSZWK2UUH+X/y2k2
B5MqDSPxzVHm7LIgHF4p8eA+hvgudn4M02CrA0eB0Vk1FjR5se1NJx7XaA/P0MoaDcr3flx4p5Eu
no0Ptth4jAMveGZqfeaxqgrPYXwZbpz/IQ4MLwZsMyXLdRaA5D/8ECDc+nHMoCPtirJvJ4sfDYgx
LQsSwRpfw+lgiUUGO5TFkxe4XFeiIXBJ1+0fkqqez84vsKc5JX/Q+RBJGgP3Dv8PK4e9JZQwUAFL
pCRZLH/CFVZZOpVni/lQlb2elN9ThJOQRLHrc4/FNQyKL3qXSs6VYNMCMRT3PqgYIt4Qn5u8c4eH
QHle3uaOGXT2X9rwto/myA09MgQ/UqeF3K1asYkCssv3tjE8Xl5P+F9kXzB8Ft0ue/sKE+Owizb/
p7K0GRWucO6Mus5jnfsl9byANhnMk9q7VDrIbudNnoDpUZ+5+Cy9LsMVcpk3lbbUBw9pEVQ5iU4F
J8QhjIWkCgGKnRCxcf9+iM9kEvXwoVLGKF4IlDMrHseTLNpokqMKrw8Pw1xzBifrPugD0v29VjHR
tIaUr8ulBd4vI3csyw1gNRWEI9gmtQVxNoDdlmHne8kifHDMyIkYe3ub6DgiuaxDg6QSeuv9ysBW
zP97hqe3p0UBQ4HGDDfRXuErzBfVHRxjof2Gq0grnj49ooSv4gGTTIpM/mDGfizKxEpyInPVprbQ
P7FcZYMS6OWlv8o9bQZe6RWt59lIBdvsIOQwtMHhx4Eerg/4CBUTxCn0o/LJ/rwJWuJkhkCc+bhn
Hs8ubra71G2d/3A6Fg75QxnB4+ietZcx0NuYH+64gCNgS5AlGvw1ibaU9aFqt7dh+iCru90WAHCC
d5ZRIem3C4mXRHXTq32OLYt2Ikwy1jrP4CFWWr7EA3mWqniLvLsiuT1vGqkoBPLqFFtwOMXL3Iy7
YklTrZma7+0SlKuXHA2WJI/VbylGJfY1gRCxXE73yZCEwyNd/zuTgK9FyAb6wyIItFUHgrpiKDbG
c9DRNZsZSPrsen+zg0pOvTWQvYCq0GYqxlZdpoLOC8DUG+871DsZvqX4Oj+MiPJjkdGji1zvX9Ds
yru98s8qAk/6YTCIWF20Gcx5YhqzbEazlfIg5+9gk4JhiXUhXPLLlzOEhIeS7VFrCgfPfkZFxEnV
S6W+XRQmIp+i0jXNaJeplaoY+bAUfBZU3aiBMvvTS7LL6Fe/P5+Z0yFkSqs8ze5HgQ4SHMVssdA1
xatHXBlABFOS9LiKrirBnv4SR8rtscBK2Ch5JAsGDxt+dTw33mkpT3XhLktgN4TresiXYpU8uJYt
AEz7fwkqmjL6aOVV2KM1xuTty8v1FadWFVllM0Jd8raQqiqT3Cwt1pswV0Pu5m7OBUcUSYNqT7vQ
jwAz9fJEWGE+aYsnT7zfebO6N8043n462g1PDayzM3BdG4QGm7DBNJi9ZOSM9Vk9GYsOWueWEPW/
p1zRqpyU/2UktHuKWaTZoTUw1vEjnWZZEDAzGwTDB2vV86z86r4DyA/4GGbpBsKzEOOXZH+LMizV
0CBQPqeDL/ELF+Q/9COJ0uv37GRFTK5KMC62/4mLvehbLK1UsCbOZJBozXPkR3e6FCoUv8/ImmaC
OJl9i89fOUhfUyEeG5QDO0fCJTe/K2MLi912HrDTsri6I1iIpbIeB/IYP6Oriw/bODetr5sDfVrz
2sL3npPRNUSlM3crk6F+lCbGkn7gtiaGNANQL11ZhkokPiZSiq3Mgf3coiHuANoXDm5BqzGu+Cha
gayLZUf7HugEz4ZD++qrD09ZqYzNYq90tXi9VyceQDgL09XYIRUGfYZmJ4b0eb0v6Y7fyZqf2J7t
pQfnir/vH0nZDv+hPvVeJdkuahPiwCg1N+fCvGTcZ0GUtuu/lVBVdEWRZp2VLhwdWa/jx+uLWlVF
USHq6WIKC49mbys9pfdO8MmvIRD6DNqsM6yJPpAHJz6EpM0fHHynrdHoy7IN0hB3D/lD4cRw5QVj
7U9nFiXngE+ZHmzAlrYKvJCWcYDBZacUEyN6nZ5B6/ueUXK8Gp7cMHYwMWI3sPGiUhIxVG4grifq
1Bd/YceeOl1Hj93DOmbRJUx0Dee++jyGmFUJ5PvCZhJ1PQ2O8byarRS/yfr9rO34jCSKV2jJvuUL
vHHTFaGlO6KxINeMufoMCZb/23zAL8KYmOhxYtg8YdCNpzVAzus3wvPDysy3RjT4cDebtzUaVl9K
Q/Xuk/nyx9dlieZXRRiOkeX9OarnARMWxrHct9X5exOiDVlnS1sUX2eyF86EdiD7uQeQj/dbUvX9
eWDjhU6NhKE135WLV8yAsgNwWywyJwQBJsE5crQop2j91xzBLRRnl4pswKwM3cxtWTPQGuNVhPEv
qakWHPbz7Dm7Wm4bQN/nHu4org7P1SokiaAgeWJY1X9weusdwoP7WfnAQu69hbT0ZipfaniTZJrX
7qd+QClBhxQj2+intd/ngzVOn1rme27n5pJlmRpKfobMSWf90D6amEIcYzQQ84hxITI6LwJGJO3F
DECm6QokO/TBPOjhn4/PwsbTPQyTz63Y9NXvSTymm+4hHPTmLUD9LCT9yoWuRoPTJmQGhpmnuj6L
/ppO2kIUtvEoW7sDBO1kQTvaI3/HXAXEs5FZJbxJxXgzu3bLO0v9NmOqiaUlLD3Y4pzYXdyZOwA7
Ts9IKCTw8d++01Zu2mkdUYKtTHIEPWKHiieckbzyNJQe+vHpfIqrsdWkJ3EmufUBq8gD44332W73
0sOL7Mk9Feuk2kqAomohPVCLEAl/WXibayzqsoACdsMFCwLgwCJSaJXINKcXHu1eUBnYF/KvGC2j
C7M2aSWN23wz4aVhhD5ThN2Q2QjAuUcHtAxL09nyQTF+sISMp4mqUmTFpdTqgDqWdyo0rhcglANc
4Vd/xzeGKH91jGsGKY3s9CckMkbagjH9P5wcbXbyWJBn3S/+9fd7h8UrCmneSCRcmFpUmveYRXQf
8oAMV7Lzj/iUzh/PlNwl1k6bFozMqzpo06YkOvFLZnGlHaeb7UDT7C+QdxmEWeArNhEhDYv/91Ab
l+zzibeXkEUVtCH6zyjEizheu66D4CWZkL/2LT7OzJIgJ27DaS6j3zOB9I8QmtWu/DR4qOY66vbY
he51A0QlLBHuqF/tejZainIoDsHptTSHtHJo73A7sohfJa+3wJficfRtO4DimT5Y6c4ORaai4SbS
2brgAqe+BlYvMUQ6oJijPvXXZfm8MB2U7sRVVP8nW538sXaerNR3/ZyYGactyMjNkSuKJvwDLqXW
eGzJg0yjaviMWhnGHAMMLIGsAXshx3ilHxUfwSyY4T3SM5V2nCRm8n7xvXwCVtZSHX8DBwcbTdtW
Kc0zSKR2shnD1/NWrp7wNroDx0QYoJUBIDaZmiAsQWTD2MY5WTcEABm0zKfO7+nGOflCFnw2UIOt
T8aXSl1b660X8hFZ5EXHElRK9nZIiErzatvRKRgCiM1wpjojCP4bdcsXhi6R3Q9ewgNOTnoXuVfn
STY1SkC7xKINnN2eKlJnJNhFdOQZIZm2Wb3/2/UqQTUFsTt5jYhCMkzAIocBKfLiKMJERApVNHKP
S0t3B7Ld7AM9oH3jXfD6asBZmsGoFT5cnsicFrBDoDfu3ZEHbQoKzvi1lEiZ5arjbZV5FZ5HHZAV
Ab+psjgDtdNkMvDAbSQgmxnHH+r0mel4O/JFsjkUkot0RJf0uCiBX/czVRNMFUVeYSzLkSi7ZDVi
sIkxXk506v67IkqWUc6G4g0o49n1SgRFqo3PEGLKn5WE4SWsjdEDJHNGS7K+8tfknsUuHKZ2FTFB
9v7I6mrsBFyjG/9u/zBjFCGTFVKCGepWI5KecfIwrzCIPFT3lU2FKgzdglq08MlhW7AMcHRBk5LD
jHF0EYIBNN7kflYI/DWrCafqCa085ORpN8l+/eAwHihK2be9oUhEQ8Y+7vxT7tg66RPh6nvotIlm
p6KlbncAfz1xINurbt71ZKohbLQ4S8G2GP1Q6azXNcHzULQTPmKdpXceNLLRCPzB8Rlq8DaPTrlN
7TDRFAIUsMKpVXFwFFJxRZM+FZSQN0kC4Lvx8zTuoNcvVtbVIKuDWWgBJTvCh5P33cEsZdvLtp4d
P5dx8IT38bQ48PTl9ovBSh4vOhmZN1T9BemHjhzQboKD2BYwgqaPTKUj5XJLVw/eVKYgoQJtqulf
eRlEi67NoRs1DCXkzr430/NXVx2X6ZN6Z697mKaebraJmDXhEiodMc6lmMXTQ6zZNSP52u4yACGX
/ffmeiNKGuUSDQ25Hd7FVndfqlTLqzAh9KIgGj5Wr7ToJ76q3Sutay5eHZ2wQ3+5L67vDhAns1kp
cA2Yc2Lq2cFELoH2Ay1Dg+4aaBjFB0a6PtBZgusfEVV09WOcjjiwHtjpnUkxE0upqHlO8gdkNO8z
abrXRPUodpWGwB5L5VY7iCAMNYpsb119OwqIU4WUrBXz7TGlyCtyiv+xwd5O2ea+4vCs78Gzcdaz
y/Cf1HY+OUjB/aRCxqJ50Lyis4N3DSMQtBv0+vYRuMmNROy6F5LEIBrZB488L+F0677hWmnvbeiJ
NCglwlB7LKe6nY+Mmp6RDoZ82WAf6cvuu3FHtbOM9fKaoNKiI5uoHa6YtMicblVMexKJkvCXvSbc
Q6TZLhyZk/04/AMxfHTr5AWRoU+dX0/wshOjE8nBhzC+ybkrST5XzdnYNWjI7yB9pW9gcxm7ue28
PfLHamm7SQg0IbCS8x1pLb89Xwd/Uf4NNqB2tG7rCw7LmiR1BotkO8AgtixfqH+2/bMcpjdaUacO
kTdOTVwrYt1Zyb8R7t3b1Zo04iGPeJOR55rTntuhUsB2X2nm2nnIyO3Zilh7Ormaul4uXE+KJb1Y
uxtnSMskR44aE3kqcHOzoaQC5+JmLIiyD4wYcFZHTixoPZVdduA8tNwQWP90HLbJV47GyYz9je7F
PFFYOL3JDwOVcWg/QmKnyIbE6I4lo2kdz2YSPtj9xG881c+HKuPD+MZg5p05RFHDZ+dALqTK8QmO
M7VLawt4OjfzT38MzwWK1WqVMDzPyjUXar6w9EHKY0F453cyNs6rCb+lwwbW9hO5zPTQ4uWnWprU
0rTUTh0PGkG4tTqujfH97wLPgXcy10rY0kyx6XSebtoBr1oloKPuSggzr5fKE5i7newc7VIGjeAi
ktdDRoSl+sq9NPDgDeR5Zvfs/0IXV+i2OieCNKijnA/N8aeWaCPJljVLaNy4Z4RETJzBYc3Tp1VH
P51IS5j2K5D9+1F83kz22S6TOOSJm9vHPdjG/ZEc98ZoOhgvrN0xkNn5S3nJBw4SPJRzNeorWAIl
cm1b8FK6VkHOrkgYjYzXAF7yrbR9whPIf+shcZE0GHAtTj8kEiiXezzwgd0lGVlLBqcmGYObLz5Q
lC4BvNPFZpql514NBWJAhf4Di/ALxKZjwY9rnHf92OdzPIHoufPWuj0XeUm0ooh1PL2QtgT4OzOl
0513Abo7P1XGvQcnSLe0D7BB4mS9gW6XVrFB0G3IMeRi3pMtsnAUUPYDrsTdp2/GZcmqxSPKP0Gt
M1PAfhnjaEFGX6qiHQtAGBWmD/GltVgGiV0fDoHYL8zXzxXxKCp6IxSBYFQovNNqeBQ+0M9YoVjF
1OJPcBJ4YW3jZp6tHQLDBYmZN2n5JfEda25KmAN0rBcvjvGh+wnSpHAE1Cu51ZihjY9EdzEPWE5n
EsUU2s/JaOoIZX3JNnMnj4AHTdGn+23qTdQqED9Y8HbM9G2zEGzh8nJsI6m8WRasBvkCaVI5rw8/
8vi1p30nCJ6R7nVNLb0ZVAnOtDe2YILO0g2Ja0qE2r7z5OqYRhO6qb7PR6tG5GRpXlcWwzHjESn9
SCrtg+aii9U3ob44nZ3y8WJl5Cc5/913oJoUU5kHtWmAWI9cCPZHNINjDJNGgoQFaYbbHrxcx9TW
XBYjqeBCA4NOaI0LmSPHDPmpJ8rMfKTbiXyuw91YDED0WAc4eg0e2B7xila+P7Y7378rspEmZsIO
Z64wDsaOJxRcdJ3xwDWTZzfQjSP3OsBvlzvbp/2648HW/bK5y3uwWl7Q3q8EFwPfmT4YGS7omVFz
UF1XGnQfNs2yNr1JPAw5sdceaqyo7V7vAA8CbCSzdG99L59SqI2WnvEi/hoMfPurYhyS86YWETFz
vw6hVW36JYb+qR9jLI5D6dTcSxpf3oEGfO9o83TkVFBj4ZldSId3/OyqM3WXFSAL6Lk/B/IH7Iwf
O3XhKYQ3axG55QvfDoZ0ycESOgEx7gOayDUlSIkhc42RXUikyjH4TejBKegVf59MYr/tuNbhRe8C
zM+G3yoHK1hh9TQDJCqouPDgxovTAQ+7idmHXnp2zXFIZoBZlm8T6hFNw5pUtJPD8Zecq4shXhf3
LPSYxy8Dg+fsg1fAobNFlXER0gOqrWDvNuLUCVPBiSTbayEAGbVQ3rCccr3YeGPmu6h3j/rbOo+S
HtrIfoXZt93NWA//c5OG8YD6naS39ZZLY/bujf7Q+Hb014zgVjSo+s2KxdL17jEPmaB9AEA1o9k8
s2d765dU4hTRC9JfINoK/avusj0vI1JCwUN/4CflQXVMr9fAjyTSD5RDcaYbZjZptEcB+680PnIV
eJsYdogOMz6lU3O76SvTkwWvhufaEikkUlsevthOvR1TtoJfRd6cqUjBwqIv6X5uBoKERic9ur70
fsO67Jm5tHu5e+3Ankx/Wyg/gHDcup0fw2WfvFloMQ6Y/t6uq2sfsM5IZmG3mL4ljTItZJqpUAgd
V44gGf6i22ap/VN5wtNRmvzh67gnAXuzkRcLFiOFIKwIMty6ZMXZ1MPoQgt7pK9paMYYKOQ099r9
PNPUA85op1BKKCyaWucdu226cUbwLfMwYvI3uUPGeiYKY9SWUc39PS6Mm2SNMF4dcfQZPBZtnBVq
0pzCSRwipMJhpIauooSx6CWHgA/5JshWjR2d1p6c8Z3Z/VvL6OAHsH/wp77X8FjtCKuPdzm1AbDD
VCWEi0fQ/ADe8NYf1P2H9n526v4AzY04l/Uz/CTopiJkiRAxzJPNcyjKul9G2xItOU/ppIW5IHqy
cBJHL2biCXpRwzHgjcrtY12WEffPengYhlORg+k1gTmX/+nApr7rzahIMODCelNBwZfAOXDxzawB
BRaVs5yw9qWWrqxsTfBPKC1qesxjd+6aPh9KzvAsKVYwqB2E7RfNj/HUkN60ivJJ4RgHw1hJhrhd
He2mP/0BXWqAFxyOUeS/9bkZk0kA7lDBYRaJTlE/TlC9pCq9diJjJkEj4oQgfONXY+50mlFZ3WcC
nLzG3CbXXq+j0Jl31Sza/rAMAtt2P+9ql3fAeBuXNcsyWKUQ2vU65ppb69slqA9dUdIYhG7anr3m
nBYRihzmb5lHuSGuNIhYxoonrBACgvBrJaIaou26xjyZ4v134UVAeUIHS3vXU4x9X8CFMOGNnayG
7y6uIiTuWKkowBoDfFQumhIPhjG0jnmcqvfs5hja/WZl3ODhxE8hxkTSwK6u/H2ikO/HpmsivGnw
p3Ee+zewVeNwFMI/+tRKtH5jZUClPdm45PZpMnVsLvv+fTnyvQFuQWY1W0/NtuHla07tcs/tm/Gw
JLRIuhdW/1IjGm5ebileCdo/sodUa8srUUgv2L42nseXLebaoWYZtTo/Mq3OLn65S6ofggh++3Kv
gyyeS4kWEsuA+W12J3d+N/ff9oZwkYe4f9dTH4SqEt3MTGo0iy6yWCyutxZqHIt3sOPVrXbuIOMt
KWL3zO07XdlIni+ZDuNeY253WaTYSf31dcc6hxVcYuHrLHVhC791ukVcMHKt76JKl885CtSELVe3
+ntxiO7jxICyr5Hh95HerV7OZ07WHiqAtmHSVtM/96l3L8eE/UZqSnxj/yDuIVVEbz4MJ/k/Ftm2
3FSczPEVI8/UfwHE94sBJHDaxDsUi13CIFFZWOeIl1mqmUcjAAsn+jid+LYeoD8oGeFLhNbbR6c7
shC2rVw22+xhzNbO0NTC8WNexgFMPYBG3qqaXpkXJdapKC/xHU5W0rdl8gL4pwX9nqaaBCRxswrO
s/d8ElzX4iz94Ps3PKvwyh2q2QGLFmt2PKxRqDJgN9fdAXIQkClw+Ka+M3nDdCJajbonrC1v1Zrv
s9/wldGBrPF/0OpGtq4sVCPZQ8/J0jO18X1ugTlUaqOIc4D4Ap1f2uYpeWG/ckf1gI3xgd7mya+X
K7QgsveqOxHsS058yhnMS2hzmlDUxPNphZRP+dAN84OLi2yCUbhtlJQjPmot+IqMnIy12xYsWgA0
Nlo/sisSR3x1CibJ4rxfmlP9cybfIoH8xF2AoWMjJ91QipJU3Ah+OEgDncZAgqjt9sCEVcF1VlJM
Iziz7LubMK8gDwi6VXC2/vmH5Ty2U91/jzBmnzg6psjISCCBasyWmrQa3W7+b2XFl0Utbgr18e1u
KzkgqSZ5mtMT9Lm3L66gLSWYxFUc5ejo9//14+5Wvb60FDYzWoZjMmHb99zBh78Sx9KIwnOpsoHD
DmdIvrQWDGNHQpa8qYr2/RvRl2XsHLyi2BbP3KPr5j/TqdvdbLoM9Ln33vg8pYamzbksrE/CW1or
Lt6pYgzE9/6TgH4p/H+RYd9h648S1diH5i/3RLnBvKUTnE43UWqtEBn2s6fsTvSTSxPKW7JCgmNR
YZQv2sgsDleaIF6YcDXrOcLNHbXdPOsvNdp4dxb7iEzmKXX8QkfS3RNjj90235ZJgvrHkuKTCh+w
01QZUL+liEly4b1NulDAS28ss5iI5Jk5amBrZKqiB5gz2BL92eAYzfDhr8JZLd/kUp+BgW106hE+
jTRrq3dqL736emt4RdhJ6zDZ11JafzeeugY9lnzL+ymTw0UirrtAM7DxsZH1AL0fhx1kVWm1rvW6
wCoHnF8jV5aRCv0h1puFeuyB3or7vKSbwAj/oG1fYuWmtM57oF4lEUasyFzlruUWL421pdBROmVb
nBmPSqxCLKk2g3PHGXF71ykKmD8JoKcezfoiVBpg/xatAoJT3emskiAEw5ouxkIthMSGINB7/Q5d
zgx/zY+QXZygEWQbvQCzD5wlvG4EVTNXKTDLsjBR/uwnmV2W349d7HrwEtgO0p+1aQuqgN46YK02
yzkADjSqCHQSH0aLFWxdrdyHWgUAQrWdNgxu7p5T/ZyOR+Bh24S3w/7lpRNfVCSBs/QT27pFXAw2
kYLZnuCEoMkokVZJgD8tP+rJrh4VlJEKaC7NtSUpKAaBjOm6uAzSLMyvEtYJ4WD+Bq6roAQwSMfU
KRlf4tWgfbVvHSIK970tbTbpFiLadkoBJOiz9Bd9WgVLI/ImzLAf1WIgaWjzw6re3+YCrYgPs6a3
AhOYU2CpaSqk8fdv5Pi55FkQtToZySHH0iN994E7a9eEh54DSz5/6OG0fQZZ3qe1PbXwkpoK/OoA
Wxeyp7r8wcr2wiHg7Ouoi2srmaudOgZXtYaUoJ40RXV0ULZR5yas9Ni/jjIpkQi2hh9sW0C57P+t
ZOZwvSjdGAQpCcoSdUXBFohxIfIKBvSj3lDujAaw/4/TYqRN0kg5yMBUXbLjklAdAZHJjlW1XgZh
pHpT5PnqBvUTukl9uxmoZeCH1voLIelWJe9u4XoIVYEB404WVZZYq1YMCKqH8N/kcj1cIaUtVu6b
Md0XY5QtogKL2et13YRoq9bJ1AGA1X1HfwPT3/MGjMifPfqDLvKnGwL7XnWj0Ei5daegfb0lniuh
WN8rnPQsoqT4xaGdCE13TJ7taBkS/S/qRNDpAHmyxVgN9DJEjOu+3vXGBoeyu8VV01qEMG02tT4d
dhu8TEpKy7vqV5MSqMFaxvun/Oxs6TnyrEcHQ6InLI1nERBTNrFHMs/9CKU3GCKqfWVGmrsBkZBu
nDwYiCQO42zq93NiN947IrGIBicj+8c0XiHYeGIlrerYig8qdVlDXKx04Q6Zg4Oz76ZBAJFemsdo
JN0vfEJ1vgpkb+js5RpuZBXyLRhnGmaBt+i5YRSDSxCNG2w0JG32nsg8UloQgHYKsgmJ+ygHBYjF
shc9of4vvChOiQyPllorZFKDlydqwWRTL8um6KyTB5Gi9J/kRGdswI7QVGNXluc+akEf3naSQzl0
eydZMcJ3U+EQiqyuXmF9rKCEpQeaoIy97XTOFzirUcTOiMwEJUKncR1s7KFvtfFd82IryexPfkE+
EwDjoUYKwfqHW6OarfIospAzY66hkZC8zXvdPaqldHAWCzaWspFPuRTmKipo/YS+LCeRjSjJqVwu
oXX6GRXXIeUYL/nNEyrTNngEkqSSKaRJhr/e+QRlJ52YQhutsosJalI+goEzeC42GOGmBe648vEH
`protect end_protected
