`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NYTO8CZzKAUSch+DxElxJz/Ql47gjQi1agXZgFy3+cNqI4mjZxtdiPw3sORZPheu3wlAPli8gICl
HhM0ZstqtA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DMa5ck1CeReBYYYPQRxEdT+4oXC4ZB3zSjVzYeAGhILJ3NSf9CzDETmWsuHqAU/D0VuB+1mliKoB
wuJxcqoQvwZ5oyP7kmbQ/sMjtArR72za3f4oEOFozLdsXXSI98QhHQ4GopzwYFTY9Y70znH/TQYL
+5sCQqCYphd4oGH6TKc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IC8r85Pozx/ukVOPajqTVyW+FohUxTtDaM+dIXa+buOEXHQsupm1NM4OEhYALzwrOs9YfKxyJfj1
PheLdhOAgY7nKVctpNlHlVaqWQkSp/S7wtreCmlScIYjHV98I9sSef8Gdb5o1aIy3xwTKwSXDsOv
Ba3N8sQO1hiTWb00xQ4/z4tzlwoGG2flRRRlrB3iJOe8gJfto00qU7b1fyaiGHLB0+vEKSGjQU02
3JnPqhFOW1tl/ACMKMGEpdvAZoiiioHku8TEHZl7SpFEDhrsEzg1K92wNh49BqVsKz9dpc9Csmvm
2M1M1pNDMp96O9H9pPKUrfHC6/RWMNNEfgG1uw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
u37fM0qAq2HKZVSvxoB7eOvs4MkPkfpFKTlLOnnnDj9NgKy9NTW912cBDnzIK0QDurP3o7dvryxg
lXtSiKcaDgZEDPCzommcHU6q6yMUqFC1KEuen/A8MvvjRsr4ezsdp6gIR9eYb/nETHYOaLko8Vkn
/+xPMJHhNm1w8Rh5xNo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sKfI12dEHTqD+z3XjokmZgsg5A1kf6o/8RvGCrpCdgCsKnDxyg4qVm9KCHvVpFTLHArYEY+IDInC
YbjBBTlLj+Kwal15k/M5wdlCd/TL4x8ocl5RrzlXbtaJK5V7DS9fI53skJcunMAQDfr0SGu9+2QY
VB9t+0Axl8HKbloQq8zOtlE2va8b7gS9DK5UZaj3ozdDN3ysrETlKt7zesO4n+O59a4UOmVou87b
uDopA4fy+NPLZ5cX/chim9PyaHAopmH5Ffkaw2KFpS8RpxlxNUPXV5rVVgoSmAffP9xY1JsFG+5y
R9DxRFLll3mp6A4MjdeUCeAF3QMOqtD45x+oKQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10384)
`protect data_block
OQwX4fyM+c9IhYX1SpXYOs72liBF1uWWRiuO7qhXBfHTc5ZsW4woj0Op5raaPCHbNyBaU+e4h8vj
jTTSZbjdXCr7nvjClzNhwoDLLrU+PEql6/9XQvv7I0RtBY+mr5+fXz0Mxcb24t1C+fvEzyd1tYd6
JJZ6tbpBpaM0A0gSubiXYpXPTon+tKR8uiqoMD2aco0wR+Y8sHxf+o4nBl02zCGvDMNFR1jMrxPZ
WKsV/28RpIHCpokowJGQin28W7xIPCMizIWSyapLS6eLC3vilqzR1SgRA2xTLjhyRNVv1TtKz/ma
Iv8Cqhw190eut04WkVIeEM47iuGrvuiN6wXfg++K9OtSmtO+Ql1yRvaNbSiea8m3cOvQO9V/QOpW
4A+upc3UY2+El2grhuFSB4GEwtAje/ALLKE2QWKY4xl97DZxV8uwXahunmarg9+iEgK4evXpeHDY
OT3SyakN2bR86YD0s+KATwBBFzvP6EnxCM4/kxsk4yUO+Qxl8ZwjF70VNA1gRCkOvi4geU/uffE8
IKQQsuw15YwmUyNhGIO7SqZpLcoczMc608+t5+TcDlO7xwcEDTFczOtlUfhDuJ/xT2CEoLfBPDXm
76HmyjcOlMcNHwgeyd06i8X/RiK14rmNDwl+ds9uznvwZjpp1GC0d3VX2CHp65AkcMDTcBUdEUbv
4EFVY48tZyIUJwKO75AwqoS3PVZkPjCFKo5ZannZDc1CugSYcesR7pJQ1YEUynpiEhFdwfqVFJEh
P3KuDIVsyW7Mv7C7StFuuPjTYXw+mvbk3/0K3DdW0f7QE+iIcGykGEbtUAE8JHnL18JzY9gnokcj
Dg+LeRhTjJPuBTmOixyj7JgkcZcBWSDl7JaPDy3TAfnC72SuqUEpE5+qfEqilQkpWGL+mFjDFor7
5gkU72pJMz0upWXF2BwNHgQS9u1WdS4IkZP3Az/zZ1rM9AJDTKadHojPko3dv6IAKl9rQNjRX/A/
Tr8zQK+iqvMOrTG9T6SZbroJrwIi7cyPttAPkCP1X2VMFWr8tjT84JMfSgDAm14oSPv9083zp7Xv
AFW6VUNVaGo4QVK+TNeDqLiQGgEEtl+764ez3kwhkjp0BfWBP/7y/VNeKf2H3tUYXqlhyqtfDZeL
XgETt2jTrcAwQUgkgsnPAXCYu8PGe47QrpLitXI3X8//pCtMAzHIfwRt+6GFzP2DKTFlAj2FOaZB
wAihkWGOJrvDNE4cOyBIPhxJzGzrVv+aglRFsa1GenwlIVWh34cqPm0mM6rVl0zrlPqLJl//1kf5
jVATLNEFR6xs1AzMasexL9aTkuFWKxB8tefqFtGypW8Ek/4RAix3ePRs/CZbDNLSRw5TvhgsVnon
mXVX4gJFgOswu9VcJ61ElkImY7beuXLeG3oJM660skDbibTAVwDrmhfJif0zN8TfutGdJEHGOWjc
H/g1ORQq5nLNGuYeV1ry/GmIiBewRiPO44T9OnfqB8dsn1nC6maz04DVpjk03X/JIinOl5c1Xb2Y
Q4YoLy/CK35Rdr/asOqrQ6A2VqR15mkqck5h9LpOlzh0wZCxmETpMNZ8Z1mRMtt1r3nk0eDuLuTI
euoNMPMVGu6TsGsRH5wfS+VJWZeL2Zb/5yNNq/vRww0x0KoAV7Yufeid2sXgfq1t+IBXNPyqRhkm
wX3qRjEwiEWQWRH5iyrd5tYo5N/stWH7XB7aFLe0FXBoy3QWWIpWe+qhVl9by1NDlNpLRv7Y3KaH
9AJmIPc3//4xXkn+bE3WJuOP3U30K1wFjC9mgZQTkXLVe+1/qvCicOawlIBa7n1IN4P5nWRLFsyq
C2KM7KYdzWevZr+cs8nw+ALTaDUY5UhJOEFrzmYqgdpyKyxi499NaXAlQJS2xYwIYRNkKhuw6CNF
NTepkDmQYRWN3whjqZcFe4Lb+HCx5plJUTrMSGUyGIwi23mN6D0sKBxjLPqkyjDJaXSdAHd92sKV
mAe5MKKFQ4GJoY4wGlSr3vYIhNSVeRUx2n/mMweaKTQlOM1BwXoT1pEEuysEpbyXmC8QQw/ukVmY
XrchFJ/k4MZjlRnCJZcI4b2kaILi3lu+St0AnrLrmWs0EGelbzV0B2uCsJQ0nOMqYFpehXJbddNx
O6ZEWw8973G4NlMFsVaBUDaFp5GB5tW+FmdsvRlC/2DsAf4o9sYARyooKYTnI7LcU2HNT3FWMzQj
d6DHzGx5quMpokkflWcHMqxVUo+esD+MNdl3r6TnP7pDYGRpH/JHlgdcWdOg8T93iLIwj5iVPE0Y
trwai8yyGvcODYvUggGTWEu1vbNHUf3dof5oAbJYql7e+SsA1D7PcNt6c/V4kZGOt79R6rDyfBUR
NeORFio4wXA75YMUKXqj1OPYwXCcKaURhErJKIafVkk1P1if+cHfhfNDtaI5uaIYjMBOgTTmRfAT
HhgInscUVOec3B7tNvxM98A7mXl1a80E9kQvkoGNl4fUQ5XgVm481Os3d2MX6XxehRAi8Ym4/V1T
lTTFFzLiEXzWrYWu5uCRAjnLL0m6HpTggBw9XNoeZzkvi44wLrrLZzJqK+lndNNKRPH0jNhJbUSi
S4em9/QtiRflgidiV3BTaxogTpeU2hmQJQnZbyhhSPNYIY1AjtbL80F3fNYXoHSPH6YJnwbXBXO+
kAJCMgxoPZCnIu7VRdYblCLBxsSEbCOCbWrFvNEOcPhn409s1Mi7ntLmd5DaYg5RP0T8y8dubfKZ
oYALIBrI3zyvxe+KTu4pnOjGXP9wZ9LGWysYnIrykmua47696kZhZN5fRPQs6EmTQBZUQbht1p5j
XGcQ1dhvwe3bWIFAAAfabZcEJzHO1/JcI3mNxtBqMvYy4VgBFTquxMQ0mihrwgN4xLjcMGjoDWwr
tOFUJHBsyw08QR0ooBmM4lk9VGr9LC001JD/szm+df8YVmR/TfUtggx8UzPSbuT0kCImfpBimCjA
J4fQiIZdhxRE2sLcmZx+xgyavUzVEheTsqVpIRdpCCG7MDrt3vyR030AF3Ok3NPdlU0/94+3Kbzl
WKzJzI/RI3dj3FlUpp8hZaj8xMt98BsCKa8Z+IZH4rHN9YVwLDdT/71brwtW/f2EGoiU50LdRSb2
LcK7bSe/euoZPvDAIKpGDqOtqScODNXeOwJ6krlvX0fzzu8YPtIvlYW9e3RYqmto4bRjTttpEucb
5ydCeh8pWGk+94RaSC2hmWPS6im8KI4941XT/Y9DtYj/QD6c4C0GZmwP0YeDUpMUmwxB5aNV0nKK
D732heuwxpqlFt5fGVuRejedN+MNtYn7hq7o1Kh5JpQr7XFw8XGK+cAgNTUrHk9otP22j7jN5U3f
KlVlw+UYfsPn6Lt93BkbQEDQLbp25JzdXRpG1A4KOnm/zrkQRCBNRYEmAzMZAzl+m7lBJk84o0xs
XLMXomUMn2ej3lEhLyDPDpqr0dEEKH0ADmVy1St0Hf2S78l8UToMRq5+GaDpiHj1umsRhn4eTTWr
tg37tl2tpW1gdcThyXeSeL0IdWp1j5Qv8WiuPLrzx+YPAPqv3roHqKaCnFHfNNca0ofRqHxRMYDd
WjOOJbGVxOetjVQHVmAY+hZ6FbOiCtw+ynNDYfL9Lwlb6fyg1H/R5ZI1H4zgsqGVAhXMKpfeZn6W
SGw5DTs5ohwv34nGPIja2xSBpF0BciIrAXI2R+Mh+86QPwq1ifDADMkgUfSj/pqvvYOPJ0R6bgwY
oJxporpdCV9N7Eo5WJ/sCCxBLmstMKP/pjChiXwaJQOY8/wSFvMlQ5h0orPEQ3Zefnl6nGekcJYj
lVL86+tw8RSNE29fEp7iM1TsSey8ID7A4rixgODDP1jXQUdJdc3tdTz124Y4VBjkeyeVdo4sdWp7
b5FWmRaXh+f4wNoiQrJ3rUsQGBQ6ljR97r6+zAyh6wkv2dVENVQevyiZdjCdV/VQP/bOeyTPAn/X
IjmTC7T/Y9bCnMipJ0m4afqeGKORXOAzjVhpZdX2vZzBDijdWLGdTHFXfDgAViJ/7v+Qna9ud9VK
cY9NjdJmKDwlbjcaknioAob7eY5Elvbv00BdQKvZ0lt6kvEWbn0rGcFlN8vyGlcMK5UNMi01xg7R
8ec0rVa6+bYFOD3Sjzs9aK9fe2dYfEA6GAHX1/tsFdp2tqUMGDMmFLggew7jfJWqiG1SQwOmyRnW
SG9iX14RPHTNq/2lQOsPKbwLE2ikt6MlKYqnJUJc+aQBC5i2avujFXn29cc4xuqSyn7OnJgaDoAj
Vn+TsiIyqFO6Bm85rIGbN1wmXJQIaFKO7RXgiTdpmJThFgnjlfYEb19mBZS39IOLEZbdTL57cqI8
wdcp+dziB1DWlGWlDKpus+qVAOaYNuWsEY1l6Ow3gyY6dKaZn5j0BejC9xtXg44eD0P+AbH/zbLq
FnRJIjTIpNPdtQ51OHgjTZvcB4xR+EPy0a/izMQe5hwy9oWGhy3iZLkR/Vowr8nRPY45NUk3pv+I
MMwxKVVxRTsz2BF6bu7yisN2j3UDlz+i9UWFk5qkea+0GyG3Ji94ELDhsTAO6Oqglpkj/QNiwq10
9hu9lSDw53ia4c/CfZ7PA3VSevaTz34WBVw0gEHzIpbL99XfQEovFHZzMFFMuvHktPRSqy8uPdi+
uYJ2DDG7TScgoyXaFVvYYDdJUj2R+iaDhEXhPFV7qPcrFp7qsz0Hp0V8xRxphwTR0kxsfrK+dU15
2xe2CrTWJypvFZln9pkHS6eI5qebki2Eb7Mqhyhtk/WTLtKL7oVyMz5MF6SzugxZnBA/CefQhfxC
RyRl8Fn4UMueoDhcs80mHJhR02VGyce7tFGlLLQfOT+nXBg6+xdRL+Gnj2CDeRpDgKpCc8120O+o
tINzcewO8sYp6trbPMZpL9Nn0i7TfPVwROb+W1/gdPUxm1by/Z7jHiiESEljOiF9dQkOyHlqw/Wk
wzdxUbwsmKAY1m2RBsFpEU4D9W/Py3WUd+B84SNrLBE2JKNtOu2emzaEqrdZxdzSi1bZKtdBkkCi
3tuvkr/B9/nN6venU8CkFgAruqBbu/NViSWeKgtylL9zF1+5llTPySZ3aaPWRayctO8fYuETtYsu
W2Bm6Wf6a3vkyUEGQS7IkpV6+pyz7Hj78tYn8d/HtIJiKO/JCswwUB+E97hFwXPtHjc9fJMcpTw6
crBrYW7XLBUXJzxvQ2cO4UiBIDepF4ZQ2e4YiV2zpqpaccmeXAs+AQNNS5teRPfU6NHvKN+KHNKR
MlQOoImzEG7z7pHPk29e93cITF6gVjfJnlhcG6iOVhWI03M7UzvTOIzeG14WkhaFnNWhnQUctaWX
7q1RbMgVVj3OJ0xfRLTVZITaU59cpjIRFhEUmhjE1Bsm2VjC2c8xR2Dd9CbIRmVTDgG+pNBmqabZ
af1Sl9yRQvltvBGAt0M1KdBfbGQZAOvGU6Kqpp+GyYZR7CpiWX7qFW/byDc9pVqW5M08sQN43Lgi
vUjrgQ2BM9LUkWSUdA33wUgGLVQafgtaslu4b2Jd0uGoE4X3V6wbbjYfZdvQsq2Iyk6wJbSDmFu8
+MhA7XzH38S8Rwqq2W2sx+KLMfmjZPa6nuguUD92qW4lMQY+G9A0r/g28xFaHPjE0vgjKf3H1luL
GcU6Yk471/5azAzsNpaQJxcVahhqJnhu1ymChHVb2zKASYgVe7GbKqFwJMzrRSlCLAVvI/yRZkZS
wkTAjXNAyxGKQeEmFrYWM0qVxBfbHYv940/iwW8++mwM7VYhXi/vvCJ2OIArpMChHj/ZAuYgVG8w
zz+Pii2qBv297wfHf0WKB7ur/EE3dlRcZXat/FMj956rEvVyXiYvsSBpCa7bD7KyJnl6CU8bAA7j
xXUywj7RhoCH/6f8of+z0g0saWXsw0KaK/essSXuK+NhtBD3vckm2TG7nMhVbr3WwMBkWaZ39+rF
LbV2x2snoTyrWQi9s0D1ZuOfoCImHECAWk8YMfBJRFN1m2W1SsmhDZOk/K7SHaOMJ9zQugGCbZJZ
wl++q9+KzC0kf0tXfo/OUdsjqWLjQ8bYaHOPGRD9+e9WJuj5ncjVfg7M9zdMsn2J22iGTS+miyPV
6rO24rhHEWYxSScmmg13cAV0pBdbeTgFeNbqZGhYqYovVSTqa0KCtzONxVFjm4diEMGea5rOTpDe
zGgV6WwRtpvJ4iogEICk+GAatdssCNwXWj44okdtwRmxFphCLgQRWf/MjB7MCuMqpFp9IPjC0XI/
rmDLOH+Swq2nzDtI+xC6P1KisIw4LYg9ogmQW4j+M6Mo/JJlTRSxvVg5RNAEQaW1Jx4pZj4fhfWl
DLcsP/2CQOb6yQ+pLg+DDhxDHDk2XTqPqafooVnr1WnmhrMUDrjInY+yEq/Ef+iMuWjLew2VsBGL
dsf+ELBL+KUjmISBtq4M1GZNwBMBpJqN5s10sHm3e4nKl9wKnxI3KpqttDRTwWQJ2cvPl8cG6AUC
dLbTZKgYDIfAeZYKNhoE1s2u+4gobuXnWEy/FF/bDJ0Cl85tv23HHVcZQGj4ZZkAMLf4eVvbHxyJ
DCnn/1vY+nJ42oiVMHISlyBeJ6/KoGfE8m4mxry3wtCAodAaY59qDJmRQc92tnz+WgZ0BBl7LXxk
0iaL89Tmj2S0TfZ8swqUwE08m9ux02xgzLHIcpCfFWYCZW4kVZxCcMszE4Z6oN1B194UUpE12GiX
a6h9jAOt674nbsMzWjA19oHgFYKxgXgbNWPjEDK1zIhmcS16hDgFPnOzszAOtnIj2/x5AYuzW9gg
haAoEXga8zsmUfQDMQLJcOYZkgg4Go3gakdCYLFXo3np6daYJ3tWktQ9YpZ4Gm+bK3tvjsuAtBrx
s81c+6g9trZqpX9MZTBYxdO6e2jAgIZNGGmNdthAsKUkvt297g3DkdSVg2E6hCKQVbEjz4Uy1ZHu
9TCcpbjiRE+x8qP9RdyFDkjJ/wu9bmKv9tqEkfTUjx/+X/fF7B8c6nSMghmKJ0y6K7YVmBI0uhfz
laXYm7G/9F7sQ4txxHGApAbL+rf/Tp23aho7Wk0fJKuE4lo+RA8RA9+YbRlbofKrol1urs9N9i1Z
pWEdsCMZyySJvt4w+1OBh5mzsKeQNjr82/hOAyDpBpXeU9FcapqpVOKj+DMKToA9M6FczKa3mKUg
jcoD+KVOpxZwhohz4QrUJZqHGsA6ZtOn00lChBw8Xdek9FYOo5xZ0LDCiU34gs9xVPkgxVGheG6j
5Pit6sfXOZE46oDvKJASmQDaCPYwQUS4WrDmE1EBCFVgzl/CBmqwVUTqx1yV9FJLV0YXfjL+t9gR
HoKLSMeMsUhbX0vvvYxzK6n0FsAZt7pjCHlaY6ARbF22EaDR4G/LHixmNYdElnERzlm0j86pGavV
VKQvqqtEALXrPkeM77g95Fu7GKBFBCQps1zeFYY2vNfqCOwVm5b0dLpS1aGn00VoT/zgO0Th7NOl
FRN6BNBnZFsLU/ah3fgL+qJAshYGTSWD47NzSjHzZz1S9mUNusvg6m/cIPFjkqBQNsdGobYOGy7Y
dKg7rjwefBYOBxxERRbtN4+VgdcMe99vX1AbFmz/7VKZvHJRTrLlJI+oO3R6LAdc9O7GDRep9JRG
sk3bTzKZyc6ZegPGWksYHQ+CVfMsjGf1uvjA/eTeLzN8KznW+f5u9QHxAhuzUd6mjWlf1p++u0DB
jp/XRWUcDtMqej7/Qe748BiDklfL+fRryCFkIiHRNBVOZvTlgU6BHKXFihtkAKm+GAAT7HYZSkwI
j36q2PokV6i6X1gwdYQDYb8Uq9JvkPHRyzllqUGQ5j3+G18d3/JQNRXEKyLXvh3mDjlYWvVe43qg
EWD+HP/cknyvG93hgebwMAlyyo3+OssII1qMBHVBlX7uZCk5bqNyCiW8U7IBmZaXvzBeLOvfjrco
1mvYP89qUlYuKGLnffO3/w6qAHdVu8NjAQTp5Cg/crG3l3gqOt0wqUkgecWdtJ4JskydPT96VhBX
VYSvcQnaWXWrZcM3UnejT95TRLkZwjBNFaxp30qeQpVWqzhClbSCkbuV1IIgLC+nxhHCjcqFz6n+
QpkkSvkm/doHiyceQkS2oKxeJrGS9OOlS+0E6S1qPm2Y58r057K2ntxJCf21AAil5agMkpuLYvCI
sQLxBNHbANrk2mfn1yIfeYwkqRXExaNWHBUdyRqwv4cGAqaK48q8x13roah+FWqjd20JPL0o0lhZ
6PiPCQWgCViwgRVYKp92IZ3e6gq5lZKEPkhBa+Ust46DcayaUSm9+gcVeD+ms/Wa8+bZPL/tAtFj
Ik6XCw+YC7nexgcNwGFT8+pNUsXdtwWVkDy2V/QBFj1BTEc6+llGo5ex+ODD1WZb2svz23mnILIZ
mWKzFBmoUauGcA8AckwjZlm+V2nw/hm/Zi/qfuKMsAy+URKrdghFcar7VhzqHW1dkJKdagUPf5fL
3KfhHvnVkJzK/OnPxMjv3bEuMfkT7mNKIXemuJGLVE5ug95zz5VoEghrUPSFSiEvu64I6taF7KJh
ffPHkD18Pd/Zugt8ps3NoiQ3mQeZxr9kJe6Lm1Pn6IAm2ICVJPeUcHngJIZdC7mLfG7wQvVFe2+3
e9k8eL4lt06UId9dGIMyOWAXeaX1Cy1TK0C3sqMyPbIy6HzhzBOzvZRnKn9pJ0b/Vy367ll2rEmM
HzS6KSCb/WCOAFkLZKcqPgkWyNzQe1raJIpIIM4+3HT4Z22km4Dhr+wVPWntyukMPjZR3Frh+er5
BbtU4ljVUZsnqLNSjI2zmaqd7gH2ZuU42vfxXkMd4UlFYsJsb5qr0QIqDkAqmQC1jxYDYTiFcDB3
VFzb7hIz/129OGKjpRy24rrTIetxysZ3CxD4Gj94Bomjz2wXybTdSVrJnZo4mPZuwPEqMmZAcj7S
F9IgTig1g9YgdRDhj879E7+QhqcVB0b30jIZJEA8dqpj0Vvrq1hpNJm6rnRp6RqsgylpWtm2wqnB
Kl+NYYXo6FQ9c0CpWDbegvHCHqWqxNbza0mYBPhBBcSN3c4iaYnjusxN+fb61btrMFBXmSSL9Mob
cL522s7DPa5BsOuz4t0x6J8uBuMCKp6DcJ1dxZZXQT/sCr5ud6/4EUmYUN/vIi2ncRMINljycAjJ
hPuQd4RK8esLNsXOJWa6nXMb8RCjldyRJ36EdhogW0VlsRrr1ktDHJokwGuwpLB4mYgZWkdAYpIk
PveoJGschS8d+MN6KYFzGToP3buaWaq+7zh53jOdHcp1k8EL7uyiXd+0YLuS9qq+qxYHKpsWiLul
JWi7GYjINw+gb2hNwZD18KGpZloVebWt7ecfW7yTroSswiQgvoHrNgpTXMX4AOeXNfx5MtapglzS
eKu+VM/crqoSf7Up0ZS0gmBeWiigpFm8oH5yVbzTB4stM2dFgaQxihhOSPgdjo5/twZxfScX/ECR
ERqkkmmz+C1wY7aMl7idUDrpgtfFbs5dudceLxG/aoZ4UE41LxH2gSnpEIpQIA6bcWfu3a/5JAGP
FjeadKqY3CZKg+EIsLXIeByiD35fDkIdmjBZ44HoNVS4X5YnUPZDTrOL6eeKkcxTZdkvR5wZP+XF
odDDG9g8AE8k5ca2gEbS6OWCn6UttM3cSVeLwFQAUaAvN02pal/EPkGhp6C10yhPbIGg1NZ2/VEj
XJRrhvgE9zM5Xej4JcbbT7+iunMljLdGka0RU3s+tmBUMOJXwmf0pac58J69DvhKMqZRRAw6se8c
6OlN0ncdYA121ZtI/sLdtz0xBGumG1AwoOwUH+0jsjaziY9XFBdBn+XdrboYXzIgEP0OMDz301gJ
yroIIZTEdYVZkUmoCRl3ind6aMS7gteCsdnssptEFPuBw0CjQ+tITOYMAIhuoGEgbO/IrK4p5qge
K7wuFjXoEuR2adIA4I+RMBZ4DoAqHXJmqzppSgTW7aLByNs1p9Ljq59lIC2drR/xoIRrF0SuXz2g
Mzfx4AIDPZSHG0mlt9wnMRhBypDOoQAtgVG0nMimHGMJ95dOlN0IcM6aiHg6hjdeKGNmK21Aqni/
CX8zaQZ4OQbus3Z0TtNfOurTFsLVaClP9ZYQIuU3jqcbJ78Izz1MLTlo2aEriahZUtuiJSWzw8rH
dJVF7+chYS8F+prloJxc9N7ZpNz5Rvi/I5BtgjBAvKR4dpm5+mj+dw2RCPLj0nk0PduKMJaZQiOg
dm/Huw9ngPXiYYdjUncWjYQZm8DonG8psKbxhsA/soaM+phDhM8PNXeecejBIm7kpJ0t7ynKtJnT
KdiNWA4QFYy9s2SivQtMhxnhcsZbQZILyjB4HZI6gZ4H9icVaJhtzeEcZXWzUl7ogYfWLhSOlC2a
rFNJiHyU58RNmPi6BgINNqbel1xZ2UWIXbUnmpzeUuZ6gisXxj8gdO+7pRSnG3jb2O74RPGOAiE1
uC2jsdhzcPN+Z7NZVNtvYUAqkkyb0YbJxBbPIspKS2aOkJmVOy8up5fr4o5lqQmE77JhZw73MAID
s3nBGbRF2BtydrVhKiNgawndF44hbSCKJ28eY+GgkrkUXqR+NlwcPrJkbFRpq+NDrUkGFQIbN+5k
dsir978AaI1KwKJ8VaB/zlfrq6H4gpGK2gagIl2wuqmC9oJG3YBTdgtLiKuXr/3sEE3zVRC2a66D
fYtIudPtfu44rDThY9xAzfbte7IirJG8GImAFeDiFpMtCVL1iies/8QaHu9DMeHWbLwVCJx2SOFe
W0A7U70ICaBiBMNzqQHLXMqn6Xa2gkThkumDqsnAA+q7RTG9oglMSqQzZUz5OEm/taWKmaW8gIGL
6AeDMmaCLwlAI0KZZ1c6q2VDH6UpcoZxJAYAFwPlpp2VkaUdq+YcmGm8QK41/RyT56q/CroFdMeR
QaQZhIcfin8fQQzkEIBz1oBLDD65DBua62kbaLNN3ZYGAI1cyIvJSUUeIMXsgCk0I5l2tSCyaPOg
kuePjYBhxqBeRvPD/tQn2/8uBgO3Zm2tR1r2zTUExtKbn3i4S+QYOt3gdpKpKXlhyRZTrEJZFQst
zg607UM6HGZYzScWC2FjL6tjak0/tMoYipAp6kB9HVCkTM9Pjl0ZSFbt+zko4D+xcwGCuy2OHW0o
9lK2y5Gt1w1vk2zRzS2XTHRtGdHP3BTeVhc7PNzrXUpXoJD8tm0CQasMzxvdEdL/NlcqzRbh+Ccp
0/TWnIoU7c63qeijEQaDmt2LB5Y6KHdR5yq/jHzLpYxiaI6nChb8AHunJgjdI0afEtBq8AWE/gH9
oAC9BgsWVczs1/oUBRPBqLRLNszILcvsGU2MSFoxnhwaMTtqbExojbiY3dHytBVnVuaN6eFkT29l
2XLAEj9yGULxLj/t/KYrnt9GDcf8CaWcG/kBHP35uViAFVjf2Hsd73z4MdvxntvEfXyR9Msi0iH7
df9Clv/XJjkbNNTQ5ObRylbmEUzOBjSZfRqgWoHo+cTerFzEuk7GiSER6ud5YsaNi/RKAxn076D/
nfoLYX6gX8r6OeD8ouaDVHl5wRhwYhvkVPKOAaB3KhrVtJM8FXzOWFjsGDHt8w62ePJ0KDtD9SlZ
jDDakwfxuPNCaMlAr8RZAUt2+D9Xd8IQhcmHOGE4MsrUiKb70gUYafvQLMZgNzN6IYQjQAsqE47h
hxfLE+goL9n7bC9BUJ+hk2naLvRm67cjTl0wiRI335Rc+hYCIYuAzI48ytTm47Duk7jyvVOHjaUn
wIQVn3voedPRkPZusmEqQdoQMheaJVM+q+xQELMf1KTqabYIXA0dqYStJUL4/kuZ2Ptdm+vP3col
OLPEiYyJinDEMZmIn4NGLEEqDbPA7mObbakFp2iNeh4oYsVknnLvVYscmPUWJFET1UeoeQgCu4gH
VnWm5mQ7CtaVgyAt7QK1hiIi01pftdVyL1454sYdSn3Ds9htilml/voNfrG+cz6bOIaxJUEdqW/p
xeOwVpb1iezrmrQn3KBnNin9OsDTqrusGo5Q59ryfDPj2HgVpDLgE2siLB8OhY412v9UlI6BJDBR
/RPZHcKCuBw86NSnIFGAOhJZGR+uhtOOIx46GW/9yOWg2IzBS9DqnJChBHgwFN6K+fpzHR1fHsD+
FiSQJQhEy+EK3wy1EdeGoDtJUd93+t5+WcmOwhb79nM6e4AUQtm0SuVdqy/62fPhPCHCG+M/fOrR
zfVzWYyxRuLnUVmSFe+QhDWMkNP4po7a/7wZXbya0ZMJwqLvbMCDJ2aeJUmQGRqYOqmfojKnPVYb
gH6XvWEvOX3PWM5tjxLzuIEdNZ4KPHcgPuizdnpPfE0bX3LGc8rOz0evxw8Gx5odUGlpDLYMph6s
VaQldPn2WZVAVsghL3vy2tWtPdIlMNH4FxSeDZcZdZSugcBnYMtODLAqZjNlbHfAarTkFJW2UoXB
QnfJWjbF/dOB2ajsDdsCNn5CR2m4WxNW9dnzE6xQqkfQuX2vaXlQQc4d4JUdqVYrwaMySYa3AP4A
TDAAprbDS07/tCQ4X9vBpaEdTe/s7NzYJTDwrB4MGjhFLo1ym3zXOEecS9pCDVE/rvN5pBH2ewag
qmlMM8DuIo4XgrRkN3kfD/8fdAhsVdvwn55gEbj/jAdSSjVor/BGiXQw53NVTa+uH49CL5J6JaPg
4H6qK4pRS/IfGP+soJeC/Gj+757yhLuKXDWllWY58iwU8AvoulkYy69/ll4Bd+1E5RD4BlLXFhgw
/euumPbecPD9IzsXaL2N68nBJftp2LWN/iA3xZjNtI5UgdKSAW+sXzRhH62NPN2AU/jrtriBwjDk
Qyv1HOurG40rirfuUO+Q3z+X5ttsF87oZUaV5nfUqQ7a1M3RueJXoXyLMEyD7xWQAlYK/7jbr/s+
wtbu1G+LIyI5qGF+Yu0vs9gIzeU+MVoKzRxcClhYJXpd/KHBs+BZvFlRioPxWLt7ytTI7r+4klgs
pHfU7nd8m5hkzVZSwxXLJdkk3kS6Pkf1VGTJkV/ZqA2mDcZr3ST07GwvWy+80GPMuw9H8TidqwXj
3LdXG966ZAnGLjbMLe37jICAc0/X9MBTHuy1Td9XOMUL98tnF3ydn6EAT2y3s0WH+zxACzC/9xrv
T+sxxN+QrblwkI34hLh/Cj67UgxTzOyrGORH9Ji6OTpz0sXkl/0N2Mv8hBE155BthoFc23cWIJhR
cBbxrq4/w7y3p5l228N/8G1zjpSfucnjEdT2ot2SQr4uuUFnUVCr3dr4rwLUhRg5jHbfiEwiu2qz
+hR1R8Cb5TIBBwRMcD3ubunTd20zCz19V/OBoxNFZf1HBbTuMtLVBcx+RbpaUis4jfbrfboUXCL3
xSajMuhxvOQTALsVSxTiKjaTHoQstyl/bLIY/O7TmLyS1CEtduJnbgQ3yjgaI/hEJux4Cx9G8KQp
QBD4Lb/E+OHFfpKnRJDde1+QP5xnWu2jjS4AcYGOIUHDrD+ZTNCd0iGkA0tHzS3una2kvl9adzP0
b6QA9/DDwH41xAb3AR0sqIWYkoIMAGjS8krZEhzDI8vhBHHtsxkOtQsu54ofZv1wpZq1vIaP1PGR
RC+CjA49/USGglKz+jNO7lXYodmFaRWGAt2J1M1SYcJHHfsIw23WTLF5PxSPKdc+g+vCYXYxC72v
jO/oLWZ1tlQfk/JPeSUOBj9/6wKvDGUW5AexP5xG8xa7V1y0i7NePtJrGIghP0NHyV2Hcu9EOHeM
q2r+9ApYW/FszY/ZX7kem93DFdqD3HiHeEHAY9IyXlp5Gz7EjK28/gM3kJgBvum8yYaUCDedL2/M
UeAcggiFZWye8k+rLTq/Gp8L1xRgG41kPzgZJ/c2Oqi7auMlbGo7HMbH8TblecYNwnZ4Hf2Iu1uM
3Mui2azwGGFU0g==
`protect end_protected
