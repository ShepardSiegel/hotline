`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YC9LzGbb9UZi+wp0HAEBk3wT4c/SdXF4j2RE1XRuwc+DAsSFcETPwR6cAW8UBEiQ1WC6VjWMSkxA
kDCrg0zkzw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
n9xexP2bwBdS569EYHSUFSnJmpcNLrMIeApi71Z/mYfGsSaaY6Bmh8GXkbVs7w27g8D6fw12g1HY
cQVsRnIkPCkbzYD/8cYjQ/Ho2gF4mIb0gIUwIpx20YiLxrIqluDe70Q85/5QbrkvkbJsdj6VT4St
SvEIykKs0FCxJ/qQxPA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZnVADHXX2uLgJjt1zDKhRvt1zEFzyvfw7safBILnPu1BTXMhiMfEtzX8xPW8pfaFh0XizN9aexyD
dCGXneWkxIdUNaQ3dLqY7r8ofnZz15tCYQez/drnvleNuvdz6jip6yBFasKtFDiW8QEP3xKapEc3
vicHMV9yUvp04Hzv8qM1ls0dK3FDPN6G5zSE3iWdaRwdM/XkZhUo75LSg8tEfd+sH9a4C61bmyQJ
gW3HEWPkTmTJbemaEDMXx77aw8Ojwu84I+gGtC6lTQCo8SbfdIz2Wsw2aBRHZ6FYcqt7HnZ1csrs
0hP7nWCsokN6dylvpeWmPH0GJp/7BhlmnB/BbA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1I9Qw3a2QXjgtFCNO2zpU/eW7g2WivrCwXCWnr2OeZe7LAfXHp6riu9LLD5fLvkPJZBafGmKA8uW
oQysvFFBQ1/BCcFPJyZQ/n3VsoPPdufwR21XgWaSPcU+2HEY1T7+Q4mfWfV5IDStu4CTuSIBKm/K
JRvOJxxeTv0tSrbXles=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gHlRyCMlCs0mHveUKvTRtqBaX6NTaxgOEwrBebU2mKWB/qBkZb6REG2VgTyaOUzo8BKY9CY3uXz2
Y+WZsn6kFG6tReLnWP5A9DYlFqF7BYLFqI9LGBfjq2brP/oSgggem6vIXlozN+xooi5NNf5VLNng
oa/L5MHaHEBfvzqyo7UT9e0RZyS2kbmhP6SZG330xv1zihNDH9EtgBcFltWdMirxFlsZv5G6YNwu
JL0Oyg5I7LWFiHoKcT1y9iXOBp/XqTaQesWJzo933UmnJmIo2zOpWnJnf4Rr0XV1McmYH7N1+fPo
bx1fW+TksbCSyfQ7TN1jvflyeeVI2KKcYgq82w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18304)
`protect data_block
7ubEeIXaXoZJfKToDzOQf0gzPPVRJBQJym4xmI7bTiaOHXNAO96+tIAibqb4BeUSWm/2h7w5cQRK
zOeWgBIl0gJZhMURE+EhNW8U1VN9eq4CvH2a1oUVME8ZBfI2p2YtmH8cZiqw55IFJlCDJig9ypQZ
aLOfipTeG0AS+nOP3kDnFbNxt7N6+Dr8zVhVMTaBQz5u//T0AUTozd300l6KKcJIaLAytacyh0Yg
aqZhDG/jhyaHvSiyu0IP9xCy9Cxx8rAPDPlbGmFEGWbU8mA89dBFshvhBZMFozAyth0jP2jFUXBT
05PathanKgSaPpx/87dwYJvpl5D6CpZ/1fgccbLQYPg7Wz0ehpWP6NG6HUON/vk2/A7L3W6mVEx5
BeFgry+PAq5zJCmxsAzY7UnhMugP/lmL4f6ENQ3zQIIud4Vy8tcggHgbuc/DQNkKrLvMT6Sus8VQ
AoTKdwpe/PoscrzlHAvRNay1DUAp/VKXiAdJqfN7vAl+ipflQ1Z797pIyCaPmygelzlrCRccNW1l
nq8Q+1HVJb3BYUqeJtLEvxtX/G3c04fN5kIiOZWr4GA/IYoY1p3lqGEgboN4Z805NLTm3XLJ+QGf
Nbo7sMO8zy5CCEUz0J8RwXMLwct/ME7/0yVRR/PJ0i5/bSHFjC4evtdaLdE3AExuGxmFj7uPKSmj
wRCs5GCpl3lyiD5Tuxw2tzawv7H1xEM93TuIqH0FTmboXdj9iMNCUOHCPf39NpWTnb45LwImhziq
hOrQ9iLG/fINeF2caIP4siqtEum9nUFxBUuWP0+4O9w5dQlDCA3w8iQv61hjSIBIXk9AZM0/30W+
M+0cD3FyBB1fzDRJK1S2/AgnKPu4XV2TEGBEdivHqu8y6wRJw69mr1k5c1qzUVdLa2ywE/AkzMcK
4peeVjI+tp6S9vsUk2ptJAbA2O8n0i8Mil8CKc88W6GOnWOP5Qu3MYRSyJY9i14/7C6ZHuyZQN26
wxTFLZsCjDEv9rTqIY2IilcH64SBOWHtprjRPJHk5bxIa8Trs3STu0gvh28xOfGoNUr1RoFJ4RHF
swikqAix32mkKCNWedjPAbi5Vp21pHHBHiRKMvSxSXi2z/XJJ+20sJSDEqAZySR68KxuD322yw8R
Bp8sohtLXxgBR2SmFucT03MMr/INQsWfp0v4UrOltdct58pZZMfZGBIJnGJIBi+t0UUpiBekTjK8
Y4ERibKAukP9k8SQD+drHrXYvvAH7fnC7lm3KM/LpShjMS59m+mJubSieEJ1RLf1FOl85YUTl/D1
ltWR6j/ummAqIIraRjhKgc7Y5JTVyHHLePW89YdnJd1TY4RUBKHSwsiW4MoEgWZt/YeNM4Hg2fQF
ikgi4glleBvMn053KiT0JXy0DYSMgtacunsoUcS3pOU5GaRPovJN5ZuclM/P8yZrU5bHu93Rjakd
Y8zDtvZH7RLLrPC5FWHSARVsIRZHMbdh5lvOSFed5bF92FRb2UHaR4wS5KdvOabrH5Vsu99aLcyd
WzT6wMdbS/YxNbdHFK5AtPsJzZRMxW/NYYxbhNxqAEImF/eKUi4LEvJY6811sgwy2GqqTJ5Couzt
QhTP6JFrI2xpHVdcBhJG8mh5LjrHa7lq/g7bVcqyzk4QUu+VJwx2l/EmiGsF1mt+Why3jD7SyeCg
8Y2n19Q+RAQQauREKcMIie5PK7iEoVawS9o7FyuFK2eq5+QqcqjK+p/kFQip8PZ9K7w0hTtrHj3C
cRIPpUVfN42NIu1KsQALjlWqgwtsoEEy9uVvHMQSpraPp+bgSqsZ2eOe0e21BgJDXwYnw/DeON/Z
3H4JfcO6/QEtj0vSZMury3qKi90nE8nGcP5ev9wkl0NCQiV2BPHF/kDkEE0NzfyqZKozwhHCUPGj
H5DQTJ/o85L/2pASUrXsUv2Z4uBaPouHnZq4d5I0gHyspaFhdqSHrds54vrc9lhac5vIpjXTH4eK
j5pj6A/Jh8aWsiQcqsnbCZJthUR5bm2leCCZeuIY6ipzCYQTzCGEBm2Snr5P2+uNZPf72JvHTZe8
JhGIDp/XlKe5VRLU18frwwvhMk8hfTlgCbVDJwoXp+Kxnhm4zUCG4eQ4vKBA0iQU7Gc2c9aGNQVx
vN4rRzIyHDEjsHKoRhH09awqpkXn1/T/uPVI13y0uRLhRTjIvHcaDoO8y2zPzG7qKysLcVrGfFCs
TIOnRRYO9KUKdpYmY3LLGg4ls/qPUZgGaaBFl+JNq3poQk5qJLLPNAPDLzZEwCClPFUTF5JKeImM
SFxMaGc2hpnauNScYUEDCPdQtk4sP6jBTBdwuVdC8lCTl/MEuqNuKjA9zu9UAJ2g8xvJX9Fjfe+7
8Tr1KNssQjHfKryoq0TmMMWmroyZdlA/Fzv+KiUJjm0IG4xgsPfhLqHCxqEpNJ2P/OB+x0ymdc00
fMMMjodGEUBuBkhk5tlRk42/n9SzqciWCotTgjtNUQXb2xuuf71vOGoOwg+GAb/zOS///BZvl+y6
QKPgKFVfJpjSMniGjwxpTDO5AOLF26e8x+yytpUspw0S0HINXoBeyif0KNFUlMgf3bqQCmjjVPpZ
FCeneLZxkC2h96U8pKxSKrEOrZQgna/3KR6I1ATQdSL+nPx3JKyNJ/nYEWdBcgw3usfzfZ+Fp1jE
LrCEpzR2/f9vt2Bb9cES0XjdyPGlnpI5YO0ij1YKpr6KkyMzBEGqyv4bkDigiOZvOAmZTCi+EqSy
ln8bQED2I/wPFxrcH+4NechSTcrOg+GVZDZtzccibnb7bvQTj33JhtvaX1cb/06gTvPSONdk38AC
S/U3YMy0lMKOxqB/VVPxrMZd3f0aBFq6+1cDPrUifPiCMbqkZAaczKgBlbSHg3GtdjBcKsKwGcP9
2pH3IVR0WD0jkQUhhMoJb9M72bbPLC/3mInAj2djY2lFCMx9GGtt/8YYbfYGSzwBgnBo6kWql4OM
xdJtsm5JkG98EdWQlpDpFMWaTCOj6zkOfEj4EiCG2KhmMJyvoRLhDDFCyilvNPJ1ynnTwlWv7Fgx
8cB5jZeECETCXZ+b0cM1ctj68dw/UzQhvXR/853EiGspu/4ZN4Exlh+MvGtjaavwq5fV2RuJWAfd
SBOaKbJ8yP4imajqoXXd0vnCMDfp2N7A1+CJ/LXZ0t/T9Wn/McfybRjIHkLk1lNXY93pnMkBcRyV
POul1c4sdeTsYOnzchbnqbCE/p9hdpM/Y7/5oF8nwAqnFU974XLddui6Rk2YLcOjY6KUm07VuhoJ
biPqH2kScI1fSmKJkkHbPPtQ4ZAuHHLBjqRCyyK8mapu1X2mXP3/au7elerEK9Uzle7qrLz4FFtJ
zztasL6XaC/l9KQiLGg4lKW7mEYWFS4RkZOm3QPORUxKNy65OrCBKZ+RQYFyvebkQi9EMpM+L9jB
6ABndvcreiV0bYAnHk0cRhLSxP+RtJa7FLpxyu6qLm38tUxOm7w6Yske61VgZQ7lfyJlgD029Q3Q
wkmcZRFs9sq4Hy0UNr5hKBmXyIzG3cCMm7gVXI2bA4cK3M15o1tagCDQGBGaLK0/d6kclDmMdqvb
SAHt2z+AjldpxptXjDPxbtlcsMjyT/HEDPKlCIUErrF3IZwT0M5bKg4kxQBHv3YE7IdUwkoCebKa
o5kOPR+wHe30e48BpfK4Y51MDSHLF+gzfaZgChb9VJzg8eQ+K3MvxwYLuqb80TPJCgcZyNStMRPz
tMDywYnSJdS/uvGP/VW0kdl5enbrlU10a42LbI4Hm0lWGqMXyzvBQq1OeYsDph8R6rMyeerDlfat
FxlMqO428OrPrMhPGkNyDcvv9eyTOiYsXD79ojpgw1WNZt45S3s2VrJTMUxngFB9CBFnSLb5HNeI
29WJsAYOUkyoEev4V3t6C/xefoz38vTETu64eHlZAezXRaHwzmkPWhoJajQRDXxDs0AV7IRSn4wx
RZwk8uIibjsM92p6LPA+5CeHxJzod0nCIlQGgGICmwYQY7Kp+XDaoT6JQh5RmNSRZYQClPICOzgm
xOnyhxu8DNXfyTI5VjJr4M+0WlxZRak5p23LsdrR9CivwEyeTZHYlfcVVaOrDdjIJkmPnaon3Nwy
ICVO2YHaby5HVbZbIiC2XeEXyW8u3r0jDenaeNtxa4xRaAXuqPaYLMzo8hGJ05Pc1U0Mp6gcIo/n
x+pM5xMKYYRIxLIpEGvVOMN6kcoa2ywY+g1B6KBGP/L9be3RDceEcGqSkCJ5R+z41ds4LdPi7/Im
n/uX7l5iUC0KYxYiXl35J/CzNkIzXLuP04Iyu7tttxIsQlRryHNL6hc9yVazMRBkEF/uym6o+28v
Da9qJVMOgzWt9FggbKSGLycA5Lk/mXf46LOdZrWCOTdNUG5TsNWAXi2PWOgGCsFro/uNFMalavep
0aoFoRAhNhhTmtNkV1b4mJbHe4qTGOy/kxow9giTML2SUksj6nnIkGqRDYpo2I1j80ztD2XTFi9f
1cvg1nxxJwRQDDxIbIg6RkXueEDsMwI7A3tKd1w8uAWpVM6oAsdZO8ZqYjPTtBjA5WFgBGN4i6fI
bhY+7lN3X0M5vsmpmrWRC6LluuZFFFmqTvdt/98tdPL7MWo/9Icsbead0eRVzjrTAE1l7GugaAp3
JSzlvvzl4e2m3HQVejHSFolmDP66qKj8uIe7xQbZiEJAY3LDeW9guVpQ7s1I7qOuXWHQtXDVMmSc
rnspW+RdRFVl7po7S7jV0j8h5QvoVKTtakjOA99Gd8vJZBllYZ20Y8E54rcM4b/xDj2U/62bVDzY
Z98BC3aYH9gQjmy4Js6Y3C+YAGZCUTIADYz6XaVuxE5qDBRhcWGajJwNQAr0qRaBSQyHtSyE7baH
HohkuyFOOmqWAGsSB5Q/ziIw5sKnMyBTEykZIcBFZ7njwW1taCY0miI3FkI9ZIeOZn4TNxkRx9+1
xrbDaCpzVQMNP90XXS+ODmYCVj6Qsv5IrOYFzZp5HXxbs7Y33rS4flItG2T+uaaFFUzQqJSptSXR
VTAu+uvVPDkpZRCpKPCaSmuxIAxeMGc0OKS1ARHbyBPWli2Bh0Vfrm5sYqihVL6kSUQ9OwzKOH9a
1/yAVjGqBgdDZiz9pr5tTT7iq30rD+0Tuv/WxnuOWEVGftpaxh2/3iw26G4KS782FNzmmmPRYZIE
wNeLJq+1Y1XfAHy8Ut8shxzpjvBvQJ11F6uHJUDtggJPZBcXtLT9vkkTr8PSymb1Xj5aIosF/E7x
GIOybCjVaNz3QXUhg7+tmd2xGz+UhZWT0EgeuFdijDOTvt1N7YscjNMULWQgNrKWaZ+wWam8dzG3
D2m0hQA1LFRtpGEQBmoJetBCIAougHGlVfBeAZ5BaaMLTBxfsDKXZbEhbX8ezKlSIwmzttLC/06a
gzxdj/YLkdBpyCDj5FID+aw4L++jNryB7tpA97Y/3s1924kYfIjZdiOWXPjwzyulkePuSsrp0yUk
MWCAoIC/zWPVDGOhp7WUBx2/wLbfAjROQWdLX9I94922ucgnEntUymxNNAQFVzPS15pG2j3fzrEU
n4jPx2LomyDGYvE61uhxDNSSNaLr5XQkIuQgmB2BFVYtPiW6v1SxmRJgzWy/bBqtlbBmxEn+5aZf
2urTi+TZa+E91Z3a5+YUoCEEPxp1j0CtajDkIDNKPKkokD5bkyqzl6P5WMDYaldsndWRlJp2MuaJ
rt4pMltAA43GC7M7pn+G6UVR3lCqCReorMpCL+rnw2foYSQFVLtKu9qvt2Kb6yqKuZYcxOEqZ5Wg
NMUqgmib7d14Fw+xlIyM3jvCMquXpRFBwBxDSDgcL0oGypTeXUcB3TCunaHobf8pAPpc0zfTgA2k
zDMEA3zMDohGrt8FtOzhKabOkhFfPDXnlVcc3cywNxB0E7Ul+L66yOagqXZCODBrnocEw2IXVapQ
S0NhuwF8zDuEQbGLHEF5b/PjtK+/JXERZIEuED0cfE55AVBE8ZWuQL2WLGOSGAYv6EjP4gVHmzaZ
rv4s+inps+VtJs2aovOQdnXCr+L3rmdPxq+ks/Lky6GT7MuKKSHvF7W5/5fnCnJHBgqvnnb3yemL
AohliElc7zNQCto+2WH7sVS1PF5GxbTnI5wSWcpkW6dX5wqyrPz0FuiQO6VJQ5/qkmD4oG3TC9lj
fRwORj3DOGuzdZp6I+8Aud0JFjDrq0DImsleAaNK9amD/3j6JOGhSHCbSalBc2QReij7584rIoIg
7YAhnJGQFn311crcnokcpvFhdbTmvuKpYUWwgkRNJDqB1OFEknT1xnSpf7mK4fjP39jpI49A6rd0
Cvlm5lxFcKKtdbq11oDsgjxeqOR65rQhOqElidStXgKcTt7lwxQRoO5ojfLVuFVdjOtns30zE5HR
7K5pouZexxKfX2K5sb2RRqZegxpY/W6YamppnFi1HBlbmXnhBRpppNILV9GsKeefe9fRK24XIGRw
ww//s+26+DLfBD/U2pA4GKifTlqY9fTMq0q5QHBi7xBwxIBeSYYciv9VJPdf35hrOh+AAlO2rVdP
N6jAFQEjX8efOgYnDaAgsT7c3TfkeQZVsu6AlON0Vy1yI/taeoCVYTXpAza6XcrxX7Icmsi/a+n9
zfPtO4av00h4Clc4iCsj6Z2K1ezGItzn4dBCpy2BN31N3j1H7yv/37eFpoea2xyiUmCw73Hmcrk6
wmj9ec3l2KgMbtaTJ8ItOlSyrzzSlzMhIpoGYOQgBl4ZlOG8LjM2ypqqrptRDxqn9UDy5EDXInY0
h2Vu0M7VaBrzqcziILBloJb/iw+aDj+LHEVQ2PP/HEzkFk2zn4ipVe8sHwYjk9mxYrDaBqFoxfev
TkixZN7zitNKVuwVMvClXgDlrJZLcCt2vSIUD4SjVI8dnijqhGdkY4/cpJfxqvBeDXNBFffgplKd
gLhSqWjm0PJ1AHy/m7qgTbf9azaXHKqkoASmM1OUIO7U+Ik2vCmNvgWt+hg5rPhjs12l3LnwxQX/
rQ2cQ+mi2uQqARia1rjAy6M9Os8ysDHQMfYDmmWojlLn0/B4ewYJJ3WfmwLJE5qFZRy58jGn1c5m
/fqhhDAmrEQx5oK0/E9tVC4NxTvppcog304h6NnlvQ4MRDUUqZzITeVuTHA8MEUV2p2bTUHAuqmc
Rj8h1AMeFlVfxB+DbK9beKeHyMr6Jl8Zp9JP6ifiYUjDuE1i8uCGsqHdU122kQ1IgzUgRUjbxkJi
3mkmC9xLohsDu0hGc5p2pWvy1cMaCCB8oSayyVusEYZOFJKGa5UzJOb6ULjvJL+fjsHpkI6kWdpe
ZCQhoFp7tUqt8nUunxovMEQpYUEc2osbFl4/CG5V3CQl9Qso/MD6o75Uc4oUvjX/MzNIEGy094gk
rEPlTxbhaMkOUXaq+gN1rbbGjnT/neJaLCJ9illGuvMCgO7j/KFJS+qcJyzs5zxPeoLA2/11nB6U
lw9VBVhX+TugFAba3/5Lo1PYqNOSygDll0/lA1pHdHaBPFVFdnwHRxdj+m1vzJmTt3tvBXrRtA0y
WKTDzb84UYU5tgvHRQSJ3KN15L1SVaTc5d0RQ0yj7L4ytYj9kY5RQ/p5wQG18mPC/E96bH5kfuLo
TgUvwLifTSrYBuPSIzMmNlww/tmuElOrqLQrJ4QVFuVfLpcvWsTaAHMUTTrPJ4mzO+xugL8X9ZaH
Mc6t7gmKmjTH8jET6Li/5rnNljrfm/WdDDCgOWOjC//R9LlV+qkf+t0r/7cZL+kFcs2RhFklM/fQ
SVitiAAKSBoD6oF4dGTn7w1uFYzHuGfs0YXZ5PbfjEYNrPsAkD03mzcFQyF28Nsd7dFcyv/x7g0O
YA82xPjxar1Cuqg/wZPrErDJdavFun5FF7NnQwES4LyYEmDYmhmqiMEvTDKdM5nr9KNzGt/ukTmQ
1FRZ3jt/g0uLMIa9cwuRjOqiGzYxozujN3cEBHL5jw1xYIJRP8KIGV7EL8+0OiJmaX74+u8itZUt
SmR+oG7tRww+lT8oHftXmucHjHA1dkPj2ijBilStmzNeofM8C1V3rNgmUH+mTfBQ9w8TDT3Rg6NQ
4W+ypuqgu2RlK6h93cda6Iv+MJ2ECyPIN2kGWpu4uHCnVObkvqE3abAFQ508pKwAmFYWnSPSeh74
v11I1gu0IROsuLCYCpYPmD580rWpY9oTqEP+AkQxmb/eSfNR72oWANTGgUuycShZ3j5gWoqzZsT3
5iS8dbZ9tC7jlpFTuA/2yE4UHnZpzvxIdnoA978+bdnOZAgvDhU1OBT7MAYdgwFow+nu+ObCxU8h
JIvut9dvWTRj3gVrs8BJpNRXDUb3+ZyfMNPKxxFEXZv4dt2lAhwUKbozXAx9rAtdstgYPvRw4/EY
TFK5w9GIS48eOimFDd9UXgg9iK8pvj0nn87HTkb20aRjJ9LS1jvU5+MTt1Ie9zz9C1K36x3bfQxQ
tp0l5O2THTo6f1EcWbi4DmrjEae/ay98pLSZUZYUU6n9HVlKtwxZkn70EnpRnLu6EWj7Jp8jNavQ
0T4SEo8j4EUwB78FSBqVKyIZthNO7TMm9RPgqzseY5ji4MkAIewwl/ZMwEwGpV774c8qRNZQhvID
HBLTAWIbOMUfi74DPt9wi5da/wEWYfQGfmkzkPEn8TDcNdu9lYPHVp8XFzc0ss6ZMF2TsCn2w+5l
MumCoYJ9/D5Uvkj+nt0wlzq8al2OzomtUBYq9elmRRvCQ9ihhUkMVcP3nn6bMGoLWddX01xdhmDO
yNV1K8k+21d5mKz81MenoEXpyMESdat0riuEXdYMjw50ohWi5wztsTvhxAoLbt3VuCCI1zKlJ9lh
ORRyAnWs9yWLioNNff3u044QiG2d5HI1VTJhPnZTOHkCvbtR/TlfvXUW2DHXrGhg88H+0Qa6SgtJ
kAF9F+5pfCmA5osRJkOnjV/oFb91ftWLPMUce/haCvql3AIJZYHvfZW1jm2gcf0BwkspFBgsfFWT
AXSX6oERD9SuqZ8J0CR4JUHYQgrYAeLYzFcEvjEy5lHdjyDsLOgvVeCAX+4KQoTWUVy6fN/j3zJl
Rlud9+PUk0BCfCgEwkFUnaq4tAhHyU7I8GRD1azQTPuLz4o3ntmnDSDVIiBTSi3rcD4tKnFFTiEg
EqQXLLKnEDsv3I8xti/NUuWxsplnLCL4gxV6HBh2NVvVvXixHsFeC8QHwroEIvojzg8pewJTLANp
a4UJBj7z7QwUsC/FydhtQxzzbEKIkUtTQ3vG+/Y7KMdizhntI/pdpVenPRLSmGNoNmWjfiOpWdlo
d9hZEuI48PDdSDQo+Q9KQvvohQEOkoY6A+tiXx/TOD8Yne2i2pBZp+RXU0EnG0j8+ZXe1xQ04kSl
gaqZ0yOGVuLiE75ZjlB8CSpr18l1dPTH62dmMLs8UY5CqEx8G0BS05qZ8wTJFwNBc/bZqTs7hcfe
Ch/3hmGProYNK/cK1OxwKywH9VyS3UgkS9mYjWgpRW24/zMpMAEoOlOxSzc17pMtbKTU8oYKd9zL
+JXo7lrP8kT5xDQMuBlaaTuy+FYX8BZTLvBmn3EZr9CHWjnyakgVcOtjfCt4Mb6+ajkrHBByTolT
fHiM+b0auSizjfqxGcjudhgmWfO++MRGsj/z0vT6z8PdjkoMz6Ban7xn9BIkBgPKkkHlZF0T56Df
qE6x8VdZRRbdLdBJsER3phnL7dUi1AkCfCEVagz5BcGNJqEQU3Rn9LrgQb2c0mKDTXCZ3JeLMd7N
ah+gFFJqTCXjMgDSszovrzNT7a6OK8rVM9BCZGrGBrbIswWaQweO4FdalpTCUOka5SUvsjwiSbdt
GIoX031Exg84lhMoSJQm/iB9y+jDsgyhL1eXUJ2ZijzEdnwkGjDH7np/TABdiSMKePewqmh8tEmQ
LRCaTgeWSVYqpAuKGYtPaW5TnqvIQ0onBbdmjO/i10MxVYmO4gBYmACEZs1A5HzgBX5CQeNRXJ7J
NS6GZ5Nd/oBrZ7679P97lUja3QGJfZRO3qyUaW+3Xwc5YiN+Q9UQF8fDA90mpFti36YTZyJC2yH8
nkz2p5H+qCViI89oPSJnIAXRd5QBJFUMEl/7LuAFWBLmHcCNEF5VHlpwhuiA2G4C/PYA0DArmrLZ
gxlc9vEBIdEMIAKCDWVfZiyDO1GPilhzHvTH/BiY1aYnTzhxn7e9N+ss5PpSjqH7XjSXiiJUfHNO
xs43mKBj97m9cRRFiyla6dFUijSg7u8JefVlg8gGquv6jw0Btb39Fetlf2xR1c/6ras40wmr0ixR
iyRipgZt14rDtpu8JGTpvCWMafQMAW3H03J6Zt5lkimNvPZTdTNTVAaGIK3PZFWZ4JwPCHcTHhxL
P2fI0RR4BVP3+76xIHWTqnMC1t6ZU3GJMXo4CfuK6rjrQBN/rNy/No03djzvHIvxRcgQ5ufUjD8M
36pmNjcTb/Wd3/EXXn+lt/ew2ZW06vW4NUVIjQNzBU485ypSGgUMpHBb43YrC8blGgq6uYUgRokY
tv4ocnt2joIJGU39fJbghinE2WXzmmLPQTHClhlAwhC7C2dWjInlvPR+3dEacsoLj7ouaQ7UGgen
GXbaiy7cr9YXGrtc+acar3wMPh8jKWu0JaRphNSMeEtFT1ufRYRz/PRhVT2yp0k/iAxVYlHJuCpr
CjFP7Aym91pdoOGPuwepSiF6WI2rNSx8QRAGSHCQj8/iBmkUkQ7Xn11LDnLS6OvRN0Z9h6FcXP5C
h5Slffy5ERCgLxSw1BLyAJhaJVApoOnj73bxtn7B+MkOyKpYOP7Pap3SKWMZfe5CCDxydJDe8YbS
T/9ol/lttzB+Xe3ROAv9gu/d7osYxlfEjPb3YqS9PuDZ6JYJ476gvv2+tg8hhheWFVqjzxo8QWXO
blY5oq0ms6L/DoyVZxlhb6fIu/NsdQTkLvUGhYcmCJGDzLoYjIcv7mF27Dh/nCljXzx/uCBXNffE
84fZaoqu8zIjlnV0/s3L0zky4831bIp51DGUUtrJobdvRya+C98/AUTl1SIJsAlXRNzhAnQktC+V
599qtToiTcqAZ/ESZWIhEJgZnXYqLKMchsJ0pCcWPAmf5qjCX8p54B/uEmjq59Liug+0+a5KHpOZ
WoKLvg4mrH7IoiIYvC5oz1jTW3wnvyZ1p/PB78sdNrgxxiM6wjb3dcMeqSiy2Cu2lqGFbC2KPHn2
lEZNRfCUVQct7v6xiPmgeAomg80BjGs2ZPZ46xmKAbln6FPeR/++Ww5YeRO/l9bhA3TkPAjo7Hfd
YSAXz65DVkvPTpqink9y4Jw7yubiqQkb3pSOSGlR8Z+wcIpovdn9lg2BQWqN/S+0mL0X3Ldk45tU
ESdKDnbURx1cN7cRRmi2erMdGQkUGHb6G70fdegNrswHmAYCB8ofs86gtgoyNayjQ+ATampvGqur
hLdqCasyXJmt279J0qjuwFBumzSqhnuDkKQrnioklvfM3lM8r5wRwDNeZkbwMKvBaMSLgfWXdAXf
VqndObsj+JMrl9l1p1J7bck1F1enzGvrbZY+xAk2CVeT27oMqCoSTbNvpWNBz6q4o+ckyPSu3G+b
nUILcEFCqsteKbbEMYyZ10YPQ2xvZEUlax2loK9yQEipPG3miq/tNxMyLK1gMAiW1ZPAY4u3UO3j
uyKrXFojGZO6yBHb1ZFTwg7VfXtHQY3lVz3DBS7rxX2LPB7jAjeleCWiUfQli2Nmsb0jltleuwo6
cUF/gOvmxb9Ydf3vh/u0HMtSbc2TIlsf8E0pJtpkQbZMoMHWr9gKP4Dq44jau2mSazFgXAgO9LmG
RIG4WVt5hLJJBVpxkv01u6Y3Pg3WFCVZzqKxGpWMfb9SerfJbb87CJphFCFZw1A9T+Y3JQfdHpBm
kRakRheECMefybpTkrPTXfhH3Jr5Vq8mbp9wgdhj7UfWvlOnpW+HQD68R1KGhDh5K2/K+WgVtmxc
c+puqpevCOlBEyINgDx9RwVc7XBuLrYTgXjASpcG1CvvY49rs4VQ2/+h7ufY3vxpownhjmwjLstL
d9u5oF1VKlr/LmjifDYO3h1+fj/OZUaLDdP81vBRBc7OX79r6SXlukZKP6NWw9T5uWY7mTFnpBwR
9+coFuDWeJYIIgHrAnJ4lhoNGbuLviIT9cTLIbe7FOeuKqj2NnmOW99WLNKKTZ0wWnlVjja4nWyo
KV6k+bvWzJQX0+DFsxIxIxjH+Gkm72WfjyUuQj3n8HUK0pbwm+rf7naXCpVXCVPvqcLNJLxPJOR4
OiGWE3Cl4oJr05GymX0q49VHUQunW9K8YAXL8A7at7yFElnf9rBuJ7gxlg08WFcHK5wuRoGXNNon
ljjEGSIobtl8D8Gzae+Y2xs32MZPTRP9JhHBH/UjWcZr400l06hpXcbUZPk1Vz28c2xX+eswH+0c
h2PBc3NuZcoqIhLTxmbmIeRRbSODgcdTT3S2HrmxU1mrmscHDM+kmdkE+HNus8roXVl41HhhsZZ/
fUYlFCF9OHoSkUJ7KkHrkJSmbxq4z13yAs81yjEmJwEY97CIsH6gfUx8jfnV0ctDJ69eoKUvBXj4
4M12y3RmWrNTXhLOwBNcEDUhPUlZYLejfFm+wVadCytNPPihtcE7yerpTWqwmEDCz39yBBA67RNT
tzg0AXeZhZ2DhwMP8kKNRBYK4MpBgH//j4djuinHXwPxCAl7nqzy4Gh3fVKOIcofmNSo/O0Lg2KW
D/JUQAg8IEC7LyTuxKgldnFIRbF2J6POtNftW7etQ8+1Ka7en9VoEAvQytg0bSo8Ldy1eiXoTful
yqccv3Jc3rxey70mNwx4Blm64Lv5TcG7ItUz5TsvkrM+4GEmyFE1u8pP15muMuH4Cjt6OG/Bxcec
rnuV01OI9oSFO+LcwHpGABDMYQtKn3kiPufL2r6SZQ2AkO3PF4ZIQl4ugHmKtfw/7wMcVtAr0gGc
SnuxgsLYrxaoX/fjVQH4eU/HH71zpctlyxgSff990S3OGyRDlvOg15Kz9ditLkUSCMg8GShqW6A6
ME9PB9WaQdOPIYZS/66t91QO69DEgGheIMUAkCh1gTq5V/SghmB5+Z44ZFeZS27VHlol3Ks/Jbr7
I5ZJZ2dKkZUet/Ge2irGK+Q+0CO9h3RliU7I52uT2I5FqoZWdAC7VSPaghfXv2KK/VBvOr7swlow
muwMdP/C8d9TaSnymJ2aY53tcwY9YDi1Fjf46ydDliNwTWL62SndnU3xsusBAkSrrjz3yOlc0jMW
xOf322v8vkbofRJTI6XdZhopOXEbS5kMfV7Vd4vRpYCYTjanY7ITBzFx7mJTjDvCXuytr/l8NBZW
RToNypqHOWw0gA6W5mmnkVYFB6f950vv/k+oX+sLlxyfvFjaLAgZFiJBcHKSNZUIMocgsW0INJO6
p9LePXlacftO8PyKYx8lmo5X/o5MbgCSL2MwCU6+hcSfGpPYCHddtQzzCtENlr6rzpL2o3vkX4V1
VqivjCzv2jo4shfFmYKhELXKSEpCeVZKiNSX86my7oIwrzM8BQShZL6qNgWT4yNj1KWRKAkn4hSg
IOM7sMdUiwF3Xakj0QnKBXuWJyxxA733fUKB6ZfrEhDpUtY1J62ioRffettMlMNpmZPKcAUtndxN
PjoKrN4BL7v5za8GWGf8zra+jy0XNeujEUi4/MGrv0Zoq2/Nf2EYs37Kh1Fv1jHNSno+ZPvlNQLN
Uy3RFi1Z7E17Gy+PeVKz0p30h4HO11SreyYLL+g+62Hmnkdj84/rJwJ5n8oNQr/DxA2qYDe2nWU8
GjMrjCIItuYkgn8e/5DdGp1oXvVq7liM/bN4xIjp2htuB2lAq+Bb54ub7QgGQf1ED3p7jG8ZW+y9
4C9sLx5Zt7VB0ThH221iSIPuKXtgtTDcIfLawgWCUZ0tDOTwdmIfoybjj7+/3Y5wLNSX/0BQJwfz
qkCxLMAfCIg8xn3YAS01gZozbycLQW3/f1H4dYimagQdueDfil0kM/yA1s7cB0A2r2NG9sh18io7
CsGc9xK4bgYPYJPyO5ZCkt5QJiZiTUdeD254tRAbQLzmM8qbO7Ln/ZQVcaE9T6MIMGFLKazOZlCL
oZqlJ0Mwq3zwzZ3RVbQeneqvN/tKTA91S8OBIif8ML+k+s0e/i20l7GrtHD1f4jlXUOJ1sUQFF74
meMt8MMKJs2spRPKWf/NL90Hq/TotUrFk7MC4TfEzoSCCCE35N2J8knUT8mXbtfeUqVf7Fc0HEnB
GqT2SuM1CkJi4rILoLD3fU8wr8me6cei3LN6xY9c3X9Lcl6JhgaADQyqmmMWggihTXJOjBQG5jqX
TGzbPcpKs5sy5qGyAoybKf9SXosLb9/1xw5PuXEGcmSuNkAdHhVvhWkSsBoOIeFnnuZlN0nIxdro
PAkCDnsYmbsNi1ag6ZBUE3e6L3iii+M3gZMmtZh/NaaDsciBDeCgxLAXJnYQll4X8AkJId2t4+gs
Rvi1kfniE1zNau8uB2f1dRARu5bJDYzmyF7AywmSGXFLC1Vtt0+IIaXMtkUSBtevbW8UZQVm+ova
tex8BbSfJoKLVVZ2i1YM8WOcX5XzILRPTVdLhEIdoYZm0s5WP2rrZbgzdRk1SOJ6J3/E1P62D7FM
EuNcBGxgfcHS+6cuEHuuXgd/cluVvQaLnfdwi8oFL+h/f96t+soc7DbyDl9631Zgh8ZQ+Zfjf7D/
A30qlawRckVmnSdc39GwnHgowwwOA7ANkxSq318HiOOth3Nwq+QkFWdZY6R3dLwOAvs7IkI5sR49
u0KbvXIQ1PmQR0HVdc7gj1dPeCW8Dj1bKSa11+unSX35aMEbmAgosfpe97z401EhmVoggq64X6IW
kMVij45l2yld+dPTM+m0cSgJiwzU1cRqJI0nDwM4GfzTkiVoPhM65HD/h+as2NvX+tnoeJsDlMR1
f0tz5xRRWrC5AB0x6kFvrJ4Y27DDlG/2hWbbFMMxCC8QbsvYOkAeRx3MjljnTSwdJ/Ihs1p+TvQg
HO33yb+Ukvih1O/5PqqJEaY/OABxNGD8Np4IvLH842uFxAVH132FddqGC8xXF7cQiTuu093QP37o
Trd01MhuU/q6T4StWtn3Tundf3bnhrn3g02w32sxnuCM+Lae33H8vkRky3ZDxEtfQpVrOzFP7AhJ
JOxzvm8cu1J5aNvmyNMjPmOFUY8mVqUgaJiPrZr1L5e+G3DHYEjVXzAK15JONPRzcZdFuEj9ErBN
aIS5LdUi8loQAyP3BKd/QH3FzCdAjYsXthKfwehUJIx2apyk9+UhUWkZggHl6F0L9Ml86jwFJDfu
rkt4nX6p58xN0NZRO2dk8RqezhTY7YX8IxShLm4PuZa8Aj0lD94r2XhCPn7Emq29waaz9IfpWBr9
nwS7dv/LoJDVKnJKMnZnaHx7o/4ssMR5cHyOIQOd80gUGu1uwQkFGT6myqR9IdrnlkqVa3gxahua
CZNspJoS2/5P5SJn9+y+oez74UYktXJcWTtm9cDDKN0VFyFDVj1QR5Ywjh6XR+g8G5cKPKgvhpyW
asodkuObcISiGjR6Ofr5/ppeNrZVAJAwHt6DLOGrRBHidBeml3I8sRTpJKLRMBmY11mwiVoRK0Wa
J0lLlldDYj0T1VcrfEv3Wgy7wObkJ76ZO1wUSETvFDbgau7glkXtA6cgStW2TC32rgViXVrhvLmK
AP2e6L9TuUMuwce3gDo6Sh7J3IrD7ovArEkXS8IvOifuxCV12EPHrA/lvYQmIVYOwgJQ7aXaIOI9
Sj/eRsHlRE4beI/zGZ1O+COlZbcwMgAklxvMl3iLvdr/7ava0eGzuI8KcmnFjaQ093r3ibRQcjLF
NvqMXl/Ue9JlZNb9msx/o6MpULvOzcOh9H+LzfbklNyG1gu35VFUG2iP32rBdhWK1XTU0dSKA7g/
KYjzFE1IMg1EhKdUlD/UuUga/xRjINQCt9tpfJld4/pbxVyzXM3ziHo2PPVa8uMuHfGfjvSiGBBl
xIYdQAq3xKI8dv5YWQYYOyZzuX9c/rOSPmzAfDJt3QmnNq/Jji/VTXw+I+GpuCNTRNtQfRRowBKP
7Rofi6tldXZFDSUQzAQnDD56Zs4kM9s4uE7ewi8QoefOsA442TtatVsC8MZE0YlMSlntQqoMtsuK
bnioea4aEt6I5hjE06q+LlRxXSZOMQ69XASUB07FG6dOQDjC8n3saddUFVKy7V/q0zoVOOY3zGm0
R1yg53eXkjM54XWzowfOeDu+LMbw1JOdnifn+DJwWu0slPV74uVd21/nW8w/EEqFTgDoUNcW+3h6
KHIAmQo77IoyshthJqBde2CfRr85EXrw0OsFzRdya1lUyf7PPXNTCf90lx9X3yL13z6SBVrxiyV7
c3ODV9KlWyJ9WZ3VXyQg9vi3fkMSDcxTGMEsvjRq9q2PSfcEA9Gi2CrPPh9OycqmZ31XwOBtsK1O
ow/hXFNcQXvkUGj3bJKk3hURd0n+FAkYSpz6whqZ3Tm2kNjqvSaU6FvDh3ySd872htEclttnFIUD
wsLqjSJKVniKao8ih8xsBmi0Pf3TroweyewU75zNes0mC8cbkoEwNzYJ7oHRiVhEOTKgHnWo7HV8
Bujfqo3XJG1AzQYeVMOfj5fSDw5WxhM3mC08UOT17ItO1KTQSVkifVDIlxWFvbQXDIgWIcWniqsH
FjyAc5nUVMaog4uyFldepVDDHRkhsmQ9Er2M8ViwnBV0BIMChTKPnqClnFU6/0/7mdg8VzwrAE+r
f+jNUxz4dHDy8qF7pFubgZmzd9U3fcrEw8hwfgQfWg4Pa9zd7VBRklBgKflIi8eXfiz+KXiaQxbk
Idx65gpD3DjwnP2tQ1L/Qlf9CBj5/nOsEslaUQjaly93eczqEZxMbp3Z2yeOnxuLvNZhGVbypRrc
wD3z81uAY7nwx5ZkBo19YB70fsxFrQrns/iqFygXwCAIs20a0H/YvkcS8ZLgkk+k71aUgDdWM1mY
4iugn0Fl1Ohn5BvijO+epYL2K6Rs/kA35nKjOZrBdKfW0PtZeSlGhIMyGX55v1jEXXW5uSlU3r0I
0ENGBO2RYI6Jzv9+ACbxkaCgD1JM+JD1dpgcbGNSrTKCrChegsuF8IZOhwQdHk/CNALynuQzy46l
yDkDIzkxx+ShDaLQgxjYToHUhx8MdvVx8yGs4XX9LpokSEk+6qap5QVPciEMpuJkft2Z9LW9fDZ2
5AI2gcyar/QJIa3Ce5lYcB9bjrOka9t8HA5Kc7eGKQphOGuK32A5TTBqUMtV7XAErZiuBJd45k3w
bCsp5fXR8GFJPfnGz/AgC20sii/pDQXepam0JyRCH4LZFAQFIBmcBOOYhHSZWWWgn0KnCWs8e809
2h+ZKfWJFtcKBSfqPxr8sgyddomvamaaeEB1ElP+dvRZdJ+sxLYdZwzV9KmA3opj6D3CE5wPebAH
AkDlszruGbyQ1NXgnVfr88OwgZr8iHGmnXLVoSt5oBY1s6HY6dooG/xTxPa/a2H8DorlOcdU6mbE
Ep2dY6DV2xhZrl7CEA4Y1nujLeiWPUNh1jqlFZL0IKLTRZQcT9WkJ2XFHFVJ4UA1xdCAItNfZQQv
grad3R+erffTbmkaWe0CyqWYd544BxKVe1cVSwMl3lhO8Z7lazBntw6bBClwx9DvrP80oIY8gDKd
kbyww81HGxRAzCW2zg6GDshObFSYxM2Sg5okw8QSnQkoJakboMMW1D+S0dTPFwnmG1rJ9KoN7aoi
8DVKjxDbB8QkBFN0w9XNxznP5+Ld9oDPnc1AsvSmWNCNwR7WxWqMHMCnlYRlj3RS0W/cWEeGqpjP
rIybcS6nXqGOwoIHZg2RrECmy9D9EZHhOk86qT2nJ9vBO3f/PGNmqGBEFRaXTNUIesTvSeCMUEKU
nNql0NmAq7nQUOlvxka4DyacIcOmd95nCX49OwUWN6LQr1+mL81l6BB3ijnJs3KqAmEOCNOPOGli
cpsBSjPBmznI+RCzYirgSGC9v0PbGK+IB0UXxH7wTgVkyPWvMnCc77UslnGGOO0p2ykjJxYSzQkr
oFQwU32/3JSe9ZsnXrn87qWoD6gxOYsfz1BbwETuyQX+XHgks7prFsnqRVHArON7njWaj5k8/Q6T
66qEV62+sVDBUNjthjO32Kr4MzkbDTtJTZ2+qNE02bte1DTE40FKbUjMh8C+IBDDYLVV+mP8n54g
tHo5VYfwnrZ2Y4/kDfxADbDuRihWRT845eyckQUW5do2Y9AUk9sZsDbv0BIxKM1CYEjux3tlrpyr
IUD+UzPVK5wgALT+O8lqLxDwj4G8kp53xHj0JGRb3ey/NXUXuhLJS1jtVBw1H0nXHaykI/E4Iz20
uXzi1Yi3e668NcirPUdDw9VK3qtH+FmITq8s0NKRASx3gy+HMQA2L1KzTRouP1Ap9v8RhTQ0UOcv
JGjEVtXmk6oDRVnZu5/2BpXkPREYZgIzFdRc0/7p5L+fjYv3WkJ/pG6F8vk7QFe+gNIT8h6Px+z2
sZIzHsek+7imweoVs4l4FJKlxAfJl3salY8mqhWVPuVnIxqI4KhdlqfV1TdiwfECEuWseGjHRj3L
tOP/T/Ic8vVsZiI7Mkywx3A7hhywDllm5k5gmnDUEoQSuG9W7YA5L9wAU+2jy8DUSdtZbkrzs/rM
hpEiu4l2zYQjMSGXSdsg7uSpQCt3nTgyrBv4M9fbPPOLpkRZDxlejbVVI6StoCY7anZinL5VHoSt
BUDIRs+Z7vwND4qsJkpw5rCv62cHVZ4guCPGoQ5UXBfDY6momYVih7aR7GLDZL7DOqHY7z2R71KX
L8mKmAlKeTT34CidbzgJETMlEXGH3UUHw+jhQu3c0Poo+QBr7pNWzAaiY31+Un40NbOx0OQL3uT7
x1+lEbx11gYoNHS31U0ebV8/YiyCrK1kNny/P8aLB22IiBblwjFJX3bg+Fz9dxCU/oM7oPQ0vHt0
yPmWNNKzSAbzBimAzYHijypEcjl58uG4eEWjbCD9+5Eva7GpvXkTQW5iSLdAxdvZ5a5Q3uMWHybF
FCxeGM9bK7QZ7YBUFUIV7JGwJJP0CB/fMGvOkvIFBQTpNZsZDM3jGxykwwa8xtBRZ4UXl9yH8OpX
7pGMpuhkushQi6MrgbI7qmcDSol/UOl4qzQnJjdYJpQvvtwUd8QUbgDWZudU9zittu2ULSoRQfi7
VBOLXGEPh126vkuo0J8Ht1KTbML+sUp0DbSD720NInIgjSbwwWVitaiXD2ZLBoL8xggs/yBkcnD3
1bPIJkVsKWkCZv4UmOzYAYjGjbH9bfxxrzU4/xuAcp/8aOqr6fOYpDzrzB1hZ+ppoa2ecNB43V4X
mgvnqQA/vPcfshxBk9VHxZUm7PJGBeppilRIbsYX9myqDLDQSMC77OG/BWZ9LcLQI66gGkVVa5R6
MsKg4QChCjHjneOXAqy3J2al7QrQrxoH+BvIEHnZHF5/Q+gClQyAottWkeELbkt2dKfRtjBhN1At
tkgiDTQyy5D6hcQaXOhIHp9ZqFNqibErKYROkPvuUnhudwNOrS/Q9mDIC6B9tSh2iUgDYkq+bTgl
BssRpVV0lxIKDUGVvM0xDgJ87oFnZoX5wob1Jr3dboMKbgY/g3PL1LXRrOyh21TPoWnBgc3fRw2l
4mLASUKzmtYVIujBysmm8PaWir80w8fbYsHrkl4hGzTgnmHr9m69M8iaegqoMjsE+CpQ+Jd/JfFG
X6IxX/pi3FYsUFv62kMtlviEW7sTs6HIIF553B7q6nNZhtnJMYSu2nzQoz5Oe0RIoWH1drRN4cYo
df0VCOdldYEnXkdyhXQ8Z+baPtVlb4zgFmnzv95QbMv99h5bp6OqefwRH8zPYYQ6oR0qk8aqkVn3
iw5nK1RTjr5xsx8ruiY+XHurU50AV+CK99Dw/0c9wpKP8MtLkMYK8HgyMz/3wFrG3AyKsv9PTd6U
kN+q3BhS4G/jB0OIhGjS3fiT1ImQguaVoeZ6tqHfVKuV7xpAPrPhPCHNt7tPLkQR19WG3hFyNeYY
KZknyqR22If9LYxVJZvjTIoIIY9roMhSzTgpUFsu7C5O9VRu7r84MYtWLevpzXocJ7JuXj35G3L4
pZx1kodZEBsv1JSRFQvDeNH8W/HQ23Vw/Z1mR3zLcyRiSPOtiX4jWp72Qtb/AEAAkRcJ5zDivkt8
+UdmdWYJyW/i0FnWHpGCdN44nk0jgL1vhcj87wm1HuAXgXW67JCpTWLx32RtBtG744L+qtvdBcyP
rFGvCsBBkAlqU28X5jQav05HZRp7XSdfZkKFPi+GxuOvylhi0E3gqUo6hQwO5xiYIeNjOK2CLWMT
lpGB1mUNatPPH22nJyCmNubHeVIHfV2rGXTJNMt8lq9uywqNfGhvSCsQbG/nvIntshxWRI+dwZsX
PSihSk9edEt0ACv9yxZKNTyh9N95LS6k+idlIXzW82pbRMCDg4InvsFH0VcI74WvTipTjyElB8dP
oLdh1dSMkofgniJioGhSULgVtnK5L2hxkTPlKF4NPxsrhnwGwyen0lxQ8B6/RJ1C/4yomkPgiihA
aSIEElYb+PqorQlNFew1iJ8rjHGb9+1QHie4suqJHsbS5yfD/673hraXpDMn050SyugqJJtRYZhZ
ds+ppS9UHPto3ve4qGM/oeh9W1oe0tA8bsmkJC1hScn6WXRkJgN3mne9Aa/xYvj7CYMsWMiEIhAr
R5NRNuECEf/y3c6ywk80ILJGPpaEj2O5qctxTdz4ZeRlMb0nDxfQq8LGf8apLIBu1As0NLw7TsQI
6Q1hxUlUGdYaBbMzvjiEEtOPFNbB73J9JdYh+KYQbAzI/Xy9HApsZ9v+EMugxtLYqq28XDyknBe/
EiSSXR/l0UM1AtyvywiSTX1dtKgS+asJaJQTufgkv0F3HpL4m8dXf/5Mqu2/P/Z+lnshn4JSE4B8
813JohRIbrF8QQXTXjtXsy2UajK/wxjGD81mMJucQ8YThhsZgsFphdYampFuhmvW/8jfnDEDXvhD
58vpbdBCiE6oMDsg+8x6QU1qonBuRppkZ73G7Aigdslv4Sz5U3bfEWarKYC2GkCpW5Bs2YoimLt7
goO9rzHOQ7kC20c0hw2OLwRZQaB4EVTE4M7dDQ1WybKANEw18+Qgumc37XU1HxtivR8S1hM0Ihf+
J5VqC6HPuKnAquWCzTp4ySDfEqU3b+MczT/o8N5tXjO+tf0IoTqq9yfqyl01D4d1i2ND4q7K63K7
ot/hlfS8CXBXNK720jzxgs81D+BNTZuwtx/77qVPMTAGSFvEGyQkdTGqEa4vtb1snoaWJm0OUtiT
Q8rXNflrO6Mgl4ThA+VVAWK3/rHXOXRRR3kCM4q62Wq5cfOqIHKo1oyiburzj5xQ0/tiK56umFDv
35Piqg00dyECqgmIRUklKxFr4fOjooZ2SNlzwLTBY6GINj3tJ4JRnLeY3NHtgxGLC2P1Av29NzRQ
d3kI2S9jxDieGGGdFViAQk9xVLkfU6CVcIbc6Rg1ZlhK24TJpEDRULib3bHb5y/anSAVtu21dz5P
GXIysK7nBTeATbV556jbY6VGfdbBl36LgWMnTe439Ht7CVqo8e9VUj0NUCKWlIAdt2FZn5zuIa1o
ZFCUE35InJ9k3t8G73JwmE2BJFkNI7FrJWk6IxcE52YV8H+mKJTq/WSlcc3ok6sPyJTIcA9S9YNS
+1OF0bR1nNdE/S+MbUEOzALzKBM7FZ6m154S6fDEtiM9QIFt8WWBwp7SDtEYJXzqgLSu8YzfQJC6
I1AjgKcRUM3OURuuIm3bsi/9sv1f8I5eU+/Pap8b5vU6NtFs4ucLucipqp8Ynohu0tapL+K4m8Iv
m8AofvXFsXiRM1UsmSPS32PRFjb7SntzIgxLybnA3h3V/OIVgLXHhBnruQNBDVVcZYVN1b6onFsZ
XaHwJn1LbB8aJ4CCD2EP6l/DKw05DpTZOuaRpSIxOtvMLuWALKSAznT2rKRDs62td6O/n5xoHVeM
54BhGeycjC76n/o/hQrwJHabyaBHYvGBaH7zlUxZCcyFfhcnAuZB2Indf64wditH7s9dGLGnqa3L
7Mi4LBQ5XzJq54JJcc2IKiZH98/LZcTG+E7qNHikqf3/03Mz/ri813VNWlzx3V5Eh8swBFV5kZKp
IqVuM62bqJEEDot/neDJGRbxHKYAYkbmyL7EWDBe/0IkkSCHoC1IzTP8ERQnBk3/Ms7xsKU9VHzN
o+d5wewVfvJFQU/KeGBazSVY1xeLXUQOQfZECvCYY6gDmTPn6Kg1UJUwFmgaHFug6auGeB3tQWKU
5pXC3fNdmGKQgxZE9aa5tXFxNVIQjbaHPTfZa97LxfecjUpoRPG7/INpVOpfTHYEoWNgrSzUBjVK
MR+oRR9E3AK0egCQEbWrwQM6/3A8gnaPAalSh492lrRlNsX9+okTScs69wU+J9yw2LPRcT7rndlf
XxMqZmnJW9Caqt+mayb/XIogwwfo2HIsQYgOz3adD3N1AkpcLPZ2vMotVzIy+vgk0mIcxONH8SCX
MwXiN/s/SppTfmk2z9yBwusmZ6fUnSp2R3DUmUMiWM8E2p+N6sr2nfhnOIQeBm4VSOKxkID///Q9
7Kf0bf9aQ5c8BTNjB7eHt2GKyYRLH5tLRLsY4Dst9sUc/bXnVAR5t7TBUHp909xPOgiIvsAUgW+i
mczP4OwP5Ca9mYlpCw/lLXj5TbY3v93t6p8zuKAh/BZ67F62h1ZKA3yoXRap28uJj+kJBTD4H7dK
7LNgrDlHIPDCDnNmzvsRIAT14S0TKMV+u7LVVNSegThCvkjH4gKOsxbyr1ygCR5Q5EGV5y6NtkFU
jSgxjKqMhR2tuA3WPRboZf1/nbG/bWCWpS+WCp3a5zBec6wh1iVf5G+fu6GAklLOpwHFA6TsFkQ4
o3JdmntJshccFiDdPtdyEHa1BqT50RZSWg5v8wAyUD7SWL/MTMKWo7a62BXNoswWqo21GBJPA8nc
SKdJfiAkUMU1L/bo8F9M+DBFy8dLyRayeKjCy0sF/J7noxAhGqkMEvuCTCgRHdSwY4g44ig+jJpu
OsYTB2aV5j5uMZCfRO82BSKgpKgJbzKhxCgkgn1UR+D02rhfX2vlAXEeNla3UNz5CjaG4VAFwwaq
xmErsuVqvApTeQyNaQ7MxRPh0KyGLcbEpdQZku0lTYFxQLFFl8giLhMXlZPRHzeQIAUIIgKrGhEF
8LNK4dCQM3KnfkfEqfuhxveillR9kPAKUUq3tc6SRN0MpZi7hBfWZWYiVmlW6/CCWsQGyzSdmPQf
wdxF8MRkIMwWe4utY/JwsAOexJhG6iLPAp1P9Tv+lRBkPlj4Qc6dgI/1Twr96jLUpGH3lHgBqV6/
CdMcdw9eo0XuCSASNM02yGIywWDSJcPmTgAFzFNRovK7kpeNFRj0uj/jGgxrAF4qMKUwjcKunWhg
Wkil34FIm3Oki2amg23CoMWP6J5tWQxRIP+itxvp7rI8nixLKSdVpg57JMZePPJPIWSYH1tB4L82
uBsNmMX3MTLpLL8UuMQv7svPpZO4dJ8CimFOt74gSDh/cHBlWPVhsaREQaK8uptDlTIXOSutKuoG
VlBC09V0VZJ04VnenOD77iluXbPRsZFh90zcok+dVejjGRMzJ7Mmqunu4ehDozJTfVcAZC8VaIs7
qUK9glDX9a0Dd4d6j1ny8ZvSMQ+z4KEyijNMTG+hG/qlij9vQFr0OZFIiAhZ+yjGFG2U4WufRiQX
SCIBBjn7Wx3TJ7Dc4MtDWc5tOra8npj4ebOSybBZOfUCsBuCs6bum9DbB8bisHubtC2sjeVC01p9
2SdiXBhFlwcoeBU51WjRc7j9/tJT/hfg7bqSQx2fTUJpv0jqrb7sL7vk7vUvkhwNtiND918fVW8F
1nkLsfvDkHDVLdrnw2HFf6a6+zX1j4uEtl3pNk3f9XrFE5NxSfMIEorDRnCLSHcH7XYZz5LBXyFT
4mGMbZ4r5JxzLmgGv8AVRwdeeyoBX3pQnny4KPnNCvg/aHyidW9Ne2S7LzOSMQXp9V6VnBIIZ3mt
UTdSmmyGn7ZsuvV0tSlDpPPv+oYn9oincFMB6hVJl6dDl6wbibj7j8kbkU/miqdIszhs4je4o+yo
h9sA9+NNaZKB1UF+5WI/HB3fYbu8jRzoDo8ukGhVNiJQ9HlNa9fAc5W3xODNbDc2/kHke/sI8zDw
6TNfnuXbreY47UHtKEdcbD59aHpvhWqvs35MIs4G/R6DLdXb7Z9FOSnHXZwjGCH1E5t51vzCWSBz
0FsJQqOrxSyG8dA6ZysPXbsfXUdkcNtIiyGUD4IVpIcD/auiLUxa7kgaPSWTIh3jpNlNhi8UyE31
+Utb6VKGCk4hGhnD48/khrIShktqb9cIM+c/wMnZ9xPdI5cuoc9zWnO05tbMzDfOL0nlrUeTsp6B
J4qISQv0fA==
`protect end_protected
