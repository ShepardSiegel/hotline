`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Kgn41iYJwdKZmKzk6iQIV0zi8cjn39O06P14Q6xWfd1U8lFfL0zkQfsHYmx7YD41yYpaCzhIyElR
brvA/TaJAQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eQVKZkFssi2td1bH3XVZ2bKFpcBazHF9NnORpFamfp2e2GF31JEZi89UVKqUs1QJiWKpYI8yEu6y
wTXhkqghOWF0KpFPDvqGmVpo5JnViuoveKX3RKzC/EZzdEBBfu2XdlQe41gRCOHROXFMc9SPq0zk
0vgLAsF13ueKCfs8ul8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LEBiQ6zaQgznFtWWzf29oa1D11GDSQPAtlwmijjKbuE+2MeGD52LLis0u5T3J4t+ZXkmBZyFKwE5
8JMJh898VEmrHIIe4iAw1n78Ohf4M6k98oQsfuiNFJkKFWMNe6xLfmQ2+lf2csdeAZ2eEh95YmIU
CjFUgEFLHzfEu14GXMju91igwYA1m6WwAh3eGPZciOFCZtX3qsnH6G6bcatgH2H9JFHGOdGbmOLY
5JLvtidYczfKQdpu0o8M7kcNDPTLog87Pxge8bDAOL0K92sX0BBuqgXZMiVyaBGoZwZsHwKf2pDU
9P8diedqzx1ofL6QJ2N9bp34dg321XzpudsoPQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
R37fjns/pPxFvJRkJaCPsw93+u+Eo1LMPVxUEGwkl/XR0Iy0qPN5sEvFiZWZVBGrAzmhbhz3o8uT
KNm7DbgFuBmeL6hEfhOA+9QaOV+5KfO8/IfiqohG5vaNXUI8xhnCkinBUsrPtcLa+DnP+h827yhK
Z4U6d/jfdI0sT9Ke/Ww=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OlMf3zzqFnhsV7sCCiA7oQfMVnJf6vtXtsceHgowwGDC0p8ScFmQTaVnVFEbrxDOaLOYNCRsPWNU
akvwNxbA/V5xGcjwep6C7CrEMztTZotuhRWLqTD87zuudEzvl+jLBkeS+dcgLh/ROJAN4WU05gth
Cm9q6GI8Mr+b/g0ffMuZuLE+cAS1CeAz27BvaxYPz9TGuAKvnRkCf9OFLDprhE7aQ/vrm1qvzXtZ
KA9KL9ah1d9CcoG+GIcBpLfs/GgiR5XvrgWCR41XfkK7ZsPftMYUbYovsnc/f2YPOR0b30P4M02L
aDmS9dglBTUftSrYu2MmrH+TjtHxRMHD9Kmwnw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12256)
`protect data_block
Zntr/az6RcpGDymm02ZbvkSnoiJAEvl/+GpKcS+lzrA2gqzzu8K4IIxjLK8uVJ+whAcIgzPUPs/5
UEyfGoqlHjxeGWdTIeIP+pAl8lm9WZw7nyYPNxPqWhEJY/WBNiOAkmNc45b/sCZ2UKAqRcXGe+69
/onEQoaloX5poeb7V8XOxnTJRlY+8WUCdVfk6tgHRh9UI461eLjE2/2Xo2tz6lYaqYpAJUCY+0ju
AKtu+gcTZfGeKZI0XTuNFX+hBzrEdW7QFTVoTF0p2SoNNAShNQBgKPL19AX/EvVpakBvHCcgY6aY
aiuwmV2TWs9l2hS/sSDWwk+2650aLQIaLDdYkkDbvyTFX/x8lGF2AojuysR36viOzh7pabqgDAuo
ZYsxnChSEbtouqV8z22TXMHV8dYAKauUth/3DuODNN5IcktNW9hz+O2xtBn4kIVaRZmC6F5JtOsQ
sNEq1LtVe5XRCt4RvLvCVdzKUpONBMsLEH5nL1kWJPqLu4mXT8kXwKlzMgQxGjyOIuE1p7BY3/7d
Clw9xdeIfGu7A27dB1r8dKmqjK0o9tWFIzizxaChlMlFuzFWOdKsVwsni3YW4Qb4aNKstu1VUq7Z
mRbkceMCAE5JZL61Xny/Gepr5iX4UqWjwKsQZ1L9P8/NmX5eEezMxPq3zxKHSe3pHrr9ayg6YMOE
Ay+Oy78gcsfn0GRMa68rUVgU/ME3Frit6w/3LSIS2X/tnpsJekOLd5ZX0GY2CWIkDrcUfKL5+ULO
vchPx3VFrVyaCTlBMGY/xHjhB6/7+DIm8kWXUxylDQ+Wtvr9aVyroE0cEBIrVng8bo7wne2YJHJs
u8groO0NvnnKDi+S1YlQcCXMbn3mP4Kg/ZITTIg21Gc82AZ9lEp0Y4EwYhW3IVQnhmCD3bvGcEkk
FEmlpXI1Yzkt/YS1TK8nEbWJUe01onsATMiOFaBLKme+jjb1OxdkBah4N2/D6BD7bpgP6zC/4n0+
5bf0yAapcYDMG7n0UmND/RMC27RvvADC62LjvVA/+l3oLE+wZYFhkscqVtn45XWLsUS4bBsJEXwJ
Jx9uAcmDZyFCNZ84artVNwutXFPU/dbc3Bv4o1F9txnJOJaVmR1veFQbMj4izutpjsOMjzXOGav9
es8G3i38hADuqyb5go/SZYm1gMC/E9CRIm+0BLX6U7f90Ex7zSd9eBYa3IxHfAky98PAuOPsk7RK
OmAWX8pqry2kRFGVTsSl8KiIumJ1FukUL2VMIm/L+YQW6uExzA3HLFIDNwck2fmyN5Hpg5w78xZB
zcoRwebYTqLQ/MSVMIClvn9AV1Svqv3fWuKo0LwqyewDYEdEIZEc4p+MrcxxneSJMzcFrLRg7kHY
HIVY9t5POA6Ht2n6sy6C3+znz9vKZb4nteLEgrb9E7OkcglNqjxMQYmYWnHRVoyYH+ZZA9V9RjL0
L5mGWqBepiCgk1oBNEiRVFnxQBTe6cEezj//3J3LbolhudJb6Vwzh4vjCCbgSHHEZNDohVJpZECs
MFVLJBdrmcgH630WuZarD4m6+cLnsw1Er5jedFOqyt64qZYXY19OmaTtrWkS3EJEQ2zaEJhP3MDR
WFzsMNscDL5t/NdulqzdlgxTpBchubxt7GrBFe15ukKa/tA0lhzLhbPP9YATsZ0B8GpcFh3z/tLt
0OAv+/8xsWBmwvdX8lOesauRVhp3iAJCU3BO9OjmJkhwSSO1/Ir43xH11IUnVJqqFm5Xkzq9mkqb
9nSUNFHVLlZbGKYBnmOP2dbMEB3mwMPaFEIuFHoh76x5I5NLeFFtRlU3YNazu2DpXlk38CfCdzEc
66av9FtdGXYavIbfz0mL31qUgxqjXiU1o1s+DeN9FMNv7B76zcvvHv3HzAfaz9mkEDkNJHeEGxeV
jzyKbm2YQrPHwCMFjunuIb6T6xQVUD7ahvsPw6pzmdq0ef6xy85/ETI9ZHW9p97V9TbzObT4LrfE
9X6U0G/VrdLvzN4tLcFXWwvwBI38wBR0WXgpErMzBKLp3YeYLrle3MglfXfJW/1Xb2o0IzLyLY0n
GfChEKeJ+fv09AK4ff0cEvxhmMvgug6jUjs4glmDOPXHL5Z7g0pNzHfKlT6VG1ZVwnPOcTgtX0U0
yEdJNitsLuqeHeQGN878qYBjpTuSSJDNrspp+tV3BLugyMExibtiGiotTnJu3sJkylbRXQ2e6X2o
lg5la5UJcKdRa4kH1vO4kYQWIzfhRFQifKTzQVb6aD7VLjP9ZPmjYi+k3PS60iWsC8HYP7uQ5I2r
MYDhKVASJISK3GeZrVZVuTIQxaCb+xhNQir1pH+IvJfsg7kCUsSUHXwHZ+W5JInKtpQxiwMvpe6n
UdGqebkx0xswPn/aJrBtpjlinymRx1iNN4WNs09Q2s08FK5Ko8p9/7o1lOCLA2tcLE1DIGTBJAgb
IFYZ59HA4MuFW5JyZd7dPyFHZcGWkgYikK3RF3UFyUGVOzLD9i+kR8aP4Kxb5xVDh6+z7aeGDK4a
ohhY4ct0zp0zuAAOuRnVZderaJVy1n3Wx0wzqViLDEyujpcJ9CP/OMh4B/NrX5gePYsy1WuRNPRL
NO9Lyz0bZtV57Wvs+S9yBISDyYaIGzcMgTwDBakuYPaB93ymA8QGQVR1CSOOlHoV48AD3wQzAl0d
ZMcurRGQayFbCIOponT8HCAr7LTQqcIUnx0kmGiMxdut8Iq7BHB4844Ftce7a4WWS7bHVnnpNouS
c0qWKP3jPVzpl6QJ0JY9wyz8LrpWWDaRjAdl2mzKIlKWBlY3NBZSMBfGpsagFIW+whYXHb3v4LSM
R8oiG8S4+TkyUdx207jrsCFFcex0K5Iv7ZtJl0328t0DchEbV0WA0hXZf26KFcHIecWcsaUpxweF
jYERw5tZdNMH9E1TcspJWVCb+TYewHwlVZ3Wc3/ZWu2DmEXYc/rdT5NxET7rQdp/bNjQ3ASHQNfI
bovsrXVsUWnp8ZXpD7lYJV29Ui73/33eI6Ht7Nqn+mPtOpQooQ2ckIqpaTnXnynHn2olGNzBEuYw
KMUN652CTc0cMpmCMECAYzmrWAmOIi9fat3TjyoSXhb+CDd4l60NKkQHABzg572oba7lcizx8GjC
WZLYdNWuwQX9zPeVUGMDX/qJ2y1iiudqWTugrbbTHVi6CTX2xK3Eup//smKsRCAKle2pcT28z9Ff
JeTRiXcsZZh+WEaUt93ND3ExLk954qy9Oc7RP423/ad78wzH9sA1+aJ4XcvPS/1piZFOfnfpuCDb
XJ35UqOr3TmTSj92Y9N8SO0veVIOxs//i/fPWX234WqZ+F21PDZuKP3KG/Hpbgm0GdkvKGsDzSbJ
WhDcG6Qxu1xPEGMXeKNlUF+xZL8+19IAT5WqevkAHS+KiMWXik7alHU0e8wtBLkuJ652EftWw611
IpnaofKpL0mHhGCjX/d9GRV+yOFQfm6YZwVJS7q7mC1YBUF6aIft3vXxWadoPKE9/ex34R9eIcif
jSYpBAuTZjM9tvsrQgvI4OSvEVd3o5WriQ1edB8ZLBl/iI0wfiZcHx0WUFmhUgj3Nf3uRO541GPK
uNZ6m7IYBaVotjjAeFFQgsOw1qWeVTc6QNJKrAlzFHHYKUH7p5mE+kJfyrAqaKUTby5+bl8WsPcd
d1h3+Y58vMIF3iVPjzoR800L4jN7Epw3kzGqoiS60LS3MJuVo7OAgwW32XIOWUQT79rsZk5qkYVo
5CwDLAjUyF6GlrkNpnyE1qkYgj7AmcufeTeoAWS5FAZsipQWX0yZMZQ4TzchM1+Rp3UPN7tfL/lo
l/HGADTmKG+EzdylM/axrl5hxalYg+9gt+I3bkMaaqjhzwPEbG30lne3dW2ewUNk9yQjtSDp1Bcp
fWJAlUCz66VruEBE4Rp5cmro5Ko26klVaKcQgWVzoVEidi36GFK6ZJKoJguJFnDZvmIiqnSw7Syg
kjgX7OWwDYG8ysYZNJ3B8BLV2MVCo4EFtuD3ssyTL473tUPXRp0utTjXGLShJbSmY9pqXOJmHcEm
oiwzl1CQYcxGwO/UwodJ8ZCqe3ziu7aav4tj/gOl0qS2SzhpKXB0QwHEBxrQioZbRhRdf5AbnAg8
fBjNZMu2q9K4ESCZVNFQorAfIi7+mGy0PD1+xNFcIkhd0+VW5LQ4eEavkd+Yo7QRzjbsddtN0BBB
FaQJVQu/dqQcbeMAmcGSfD4vfKIyoABNu8EA76UqQQaAfKhTCvtB7WmgyvJwe5F4Ixwm7zu8yNFs
TfiK3P4rKkTgPk4A0NPUZ96lcdnruxqeUFqfwGXN6R3DvPOCIa7gm9/gxMspYMuLhCQtKkJleRb0
MNosljtRixZnYkqCCtpM9ceXNDu6VgcI9j07/EaBPnMQtIEpluxW318rVLR6llRsPq69gamY2GfD
jgbhCt7o+I8kxAdTA+wBGNJy4Anc8VAQNKboRHeeOmlqauZAISSJy8NJe88Sr5JHFwUPmUpJ/psA
7oYXsptSIsGfBqfhX/PK40uPmHhXatEvrvShkJJveHRrWTkJ5wQXRXbtO/+YMnm2pxGYHYfxHbv+
7ifo5usrePuKVfiSMW32Rl6kvE6vCsAcfN0xyiaF7rAa8UyV0MkjfhpdSX/0p5PByGZ+cPaBITEA
pk5JgUFN+280YuaDBNBvjlbbblL8CbUvt0iyXSUT3c4Gj6tYNLVC03x+NqW23EFBKJOVYwrzML0q
JUC+7dM9iGfCBvBoAkvE1REwvtneHMDnzNmtpzg3BUJvQlw8H405FqQ6EiBKkc2vfE62CcM8zqwE
YWHZ1/RVWRbQk7E9mrYpird5+txSuuFeTS3wSklCD5rkWvkLegSMe5IfLauQ878UU4bFtgMP0sW8
g0l3hfAFyq67wLvafSrhcb60GypzrU9cQpJnCoN1p2lk/eJwK/FKcq+LRoyXZT2QHRnLMdbYOP6Z
Eqw+1T2yC60I66opnExq7StEyyv9tkkZNTATVjvqKDhHkAN8H1tnX7ky4JL85qPH9fJYSBM9yryp
xqEdh8Ml8RrlE0N1LoYvc6yoi5BUNgwO+9sL/DqpRahz9qlJ8EiVbIgx79c0W+OZ395fo4KJjzwq
zyEsGmYTK5dCTGO9zyRR0ZLk5qqCpBTYB60NH1KBqLsKm1TY9/TDqjdkg27pSHFnp/gj7jsxuFLA
3M2uyxJvwmIGhTJ10LXe+ltVGTOLUZv3LNWPdmFNRFopGXq3qr6bFQmeOZ5/2nITFjXvRi2g/FdA
4r7MQsDZgCzIo7cM/ZVtkzCpDalPDS6xvFlF89bHbBAtxfKtvW3ekdrCt0sKwNT82pWTH9zTFXHl
Ry6Snum7JEInunqiguOOnTna5O9ZOVgBqJM9QOHiGv+m2u6iTAG9w1FpobpzHc/830HZeKIJg0iO
b8uYozLo1L1RQxuT6mPrA1AHjiEIBDzovEM5FTNvjrL8UGvZEDNRmsKk/kNW8G2ml5CxOW82AhPs
h+5XgNQOCAarHeBJxHkVmxX+MX4wTS3eAhNfyuYuFiHzyqkPNSJnUVgYxva8daYvvmdQWM9uM/oU
aP9P+dVEvNeDHKcr6VSfuq39za+DT0qOcNaKbuuLEMC7+xb4NOEp1lFnCjqjCTRXsnRY6TaQDwsV
fVJMeVOpljz36TJlZASt4dLMhhXGpC0K4v6DayIwVeAqOqcx3ff2Qhvpounuj1plDD4zXxvsiGkk
tmhLv1XlnN5W8LXiRNOm+rfnkEx4bD94U1iwmNcc6jxgQYQuOndyTWUmyaPTe4y8ZTLVIQAlySTN
5PZ8ZVtQjVOsd0eacHjSFWavse8kDCGZHCGZ2FQmXNI3uhtY4JjvttYmypZmTuKr49k14Lz4vuIE
rgl22njdSdaMr60CEbyb+wfR0lMNKFGucs9k52UGtaiFbyZ1U+L9IfR/Ql7ZNxgSY+Ql4dELv/N+
Hd430Hya1SEVEQWSqAQbGauTJaJuaXUwTtyegiygNr5TGLuevgHsC2k5WYjcSplqtl/AIanSwmJe
BEGATuiEcODVDN1/FQsTB0xDceN1qzTIXD5Yxjs0OenIsbfV/qXsCxCwx5L3QjKr0cAHCv1HN+Ds
u7dmaw32xElbWvnxNth+IJq/OHm5Q/wpxFe6ZRsAdX3UHHDtTcd7wo4mjt10ACq/YDTKIkL8FI0Z
+mXeroT/iCZOw5+aKZBp4FqtW0dFE/n4Dc+aG0s1Sa9XKHZ1+Bqo/ogKXkTg3UAChH8ZkfZDR2fE
VmHGUZwFSIU/R3aYPpG/oOLUKjLiPJa5JoWkxAF8dUxqouzId9sWoDxjiJJJPjpbIjTH/5dVf4Hk
tcvtVO9I7Z2vX9rg5pQjXcdmof6feXiHwhyz+H53vUqHSLiQKOCrLhW+I0LBOoaceBGaTu+iqSpa
JcPLTXX5KrAWDnlg/BF/M+hikzx1PcYrz2A8PZiUtufWfc01M9obap/m2x6lsLZtTSLjQhIPfaNY
dh5YeNPtoej/p09/bB0NvrPhYv24BnzxZlqW5Jmp88E9bwqx3tN3YRDjmFK56s6sm9L7qiPbuli4
4AnJStLixrsa9a+/romnCC693fazVFmSsV6z0As0GwilLlAzVFTTeGX4YpojILjaWGvbMqgE9x0W
NPj17DXkxtknSR1dUB48mIlVJKJdA8be5j2u6KwOZh+jPF0Ai/laWTMJBB5NXb7W5kU+ra8Q77i/
WiXDxGBvEeqVEtm4Lwb3J/rpw+1Hzi5QOqWP4K68B8gKRnWIcJOwV6N+va74jsHlcqvvilGaYqui
IPMdShRe9U/GGFOk1L9D/Cqvpdq6SGv6opW66ppJumIwyACPYV06and+OV8od+ny0RfTcOFfV80I
LrVwHoqgn0h1wMVO77myZYdaBzyKGN+6/GdZl3FIFyCLML5BZFQkWsh6NT9dczhYQYi74VxY7gD6
fzxYV/IDSWvf9pJLO0gSO9ee7l66zJiVsNLPATQ2wBMT6tZbyWVbpB/qRGY9u0dH5xDPs6lDBfJL
1JrTed8m5pRem9oWmlGFdzNAfZIRBoZ6DOaieFA+w1gzV7+JOEqdXPdfDF1r21BZnYm949u1XPAX
yVA5gk6BWiNcGVybX7bwt0oJNw8MU3TX4vILjcrgSuIAHWFVE5dtyPU+o/A6YK3iO1d8TOWGZUB8
xS2RaJ4fi21c4POV+WqHwl8wd3UtARGWOtDaPJDvWYK4isYmOFGAYPkTiwbXHsD/U+fbb4g/qW+r
GZ0QZU86CbF/MdI2fnbQba26rNnbVAZNxvndTGchZZGupd7eL5dfYl2fDVphj0taUpONz1by1AGS
YdKhh3RINZftzu1dzqq3wihLcb49DAJSTGRzSsd8cEHezgDOnDRXU4OXknwiAj98SAcRwlQmScNA
GRZsCna4PDiur1EiXOoDDsiMr1aDb7y57f06CeLbhc0UuLTAVtJ2n5S/e/ZF15qWEw6QLGzOvidP
3K1zoEn+ZDZZnMuDzoijUKiF6PJtVs8miy2aDJlMm/OQrBviTQt1mD0i++Gr55kIKqJRQUy169A4
HdjEHgTmUuuYrTfIjqN+3IX9dJOuGabjgvDzXFm2nJ+qH5ezvBJDdcBQPpjnsM+GZv+Ghmy8H0uF
NOSHjGceJ+G6B0NJQ+frSmoA3xsq9KBHrF6HEDZJC3QpjZZl445Xw2R1Am/mfaVPVshQ/hvYsLjZ
xUIc57mqwuoR/5VmfTr/bshqNM1XA6EOE5We0XR/QviE6opeff6y2eEB2XbPi2eShWE2GnlcSAWD
bkftUBPR9Va6J/IeWB3M4tIAUfY+RpBMZo5QTzuzAJP5Wbi7i4H6wwbDQWd3b+X8dxx60rpdR53W
BHkWF7ULMuQOFjG5JdAHVfY9+nk7+ePeWwYQOOZvwfSnHdYTPl9Ve6kEkEpXkxiIw1PhxEEL51w/
DLSAHdySyg33SNy//lDea7P8cecbWle+3L4F4Av5818j7WhkUQ97PCYonO2ZCCbsxTgb5izlWk8K
mQacDCTPKx0LhemhmrXM1WToPOswYEKEQwG7+Ex6lVdAkCHT6DoKV3O4UcV3ZARiVXa1tWqQcu9x
SUW8FsBWhiDo5bAaB+YB5g2zCuRnVZbsGEnBmqZi+MsNw5VcXtM1V/oasNyAGLanTNZxAg71qnvL
wiXpUnqMMdyKsr+oTJ0o2119LVoTGTklYaSeRzimuFfp6p+oybrSNGI1DIrkIhrqdlWdTECYgWyS
6yBBKWIOnfwrXLrosGKsb5yoYl7mqKOnAIiN/+G/haOWnVN8TBDv8CRuoOQFEhTkV3iFrttn8Se8
Bzt12W0IoSgP723sUHkcnqaq8nLmIN5erlui2VfT/p/4a1SoHZ7u7mDtTl+Jd1diPC8Wed6Kg44P
TAeR59+Am2KIFqoK6TiRbZtiDWGXfvqTpK85UEpZC3au0B0JWEzQ2TWAHsD+sNSzxGD5E6b67amx
j80hiFOAnHfoiJA1ktUZWuo5x4J6OlQKR+kbZ+aODoCkI807dJYSn7K/otOhVE0oFsbyKMIYZiC8
WNrSnoKX0wBbboKMTspL6WYA2O5EN3GENiEjQ76NmK4cPyDS5VTSWq8+7LPmtrMvgijyn+FRO23/
dv6knjZMmmB3Q7rYHenRvsB28v62xTmrUE5W5KDiNzsW+ViIo4tzEYX3F2bnM3KsjR8/mc+hlfiI
48+PiHXRn0vR5O3qbWty8CAX6dpP4nT3/CtGKXr4269rm4Giip7R1bZU+ujygEkXnfU0m0DZW6D1
mbwjKJS0Jbl46Byls1ganj+edvbdSDiDW6cSGFWYpTbBwFWu2jWMNIHm0653i+KyF/hOObz2QTVV
x1gwyWjnkqw6+XoLU2Qj/HTO0MaQZVRX/znnatlFG1Fc25xqMhNhF9mj84vOFhDrw63MkA1Lzc9v
ta40t0gVpfDjYBNb/ec45AAA2yLjYA3Nk5NULWcaYftfBD8//WfKu18UmNlpijACeET90FbP0rhU
UOn3SceeFm4wZ7f0c+z/O+hneDHWW+H20t+q+Q6aDWkSuww6aLZcqx4d/DX3ZufBEcCU7ukL/KX4
mEWwooZgcbrJnjI0i1mnMReXjFLJyu/phMy7ahe8Jdm2NXoclFPc3Mg/K4SCXeNY87dV+pC15dfY
AWUenSOue+FZ7Ztp+1UUInlkysDkQfZYQw3QYJVOUvtLbNEaYxQzcx8Tyf0WhqwJnL6TuhUThcGX
713HqMFs/r4G+o7luZw0lIAiu2W0dAOT0IQNdgxnRXkGfblBpz+Z5vFdoLS3uA0vc4isE4dpSszP
5gmsRth3SmViA3015oCkZQI3XTcqHxEiHG6gGRiZl8Awqae7xjVZARfHj+glpIPS1BlFa8ieMWi9
s1QniGYiStfzryejnTWMj2cNqEjShkK5Iqu1+U+G2Q88VbRELr0RnPFQNPW4kDz4mQdLgWmTFUfs
XRIoZjF5I+7TWgdluCrRNMMfFq2z9XhpJfMlbCTEVmw1uJEcRg3raA99LjFXtL0Sq0qTvZllaHQr
gw4V0IwAjmg55Mg0LgLwa2pLKhxWKA01FzlkwsRhApt7KAi11agp0Es6RGu/4YzYsQ4O2bvAOKf8
H2+3EPJMgvzmjmvZl7zkhGBxo1qq6j/TAN3VOAW1UCpFtK2NtuSzEv8bt0SJR51qWFgvZULNyO0r
jUAAXQKUzXMpBzim3zndeA2VhjGB/86D4W2W62tX4KlXeuagGrj+fZ7iYsR+Z8sJsOFp0TZwuZUI
Ht6NiQ7U/Rhf3Yseh8UVKroeL/1YoC7mta8d+Iq+eDRn9gDhYGfddhivyVYOsjZcljz3T4V6zSaf
uI0pwZcp88nDwPIqxYdA+0g1lTLedKH0ENlJifXLctPlaTiq1aRflL/GMbE013CbVobojS1CNAIs
PtA+oTeUpJS0uqX40zdrItGPJ0a1mOOMq9XdxZ3J2rrR389zUbxhdBBTiqG2LUBlGt6hJMvzQKmE
I5tiCh0tmcie9/FmJ+f5xAuK1IO3TWULZn2h/wrCaDGmodrIe0BlCrXfOlcdzHKl2x4vg67VllC1
BfGpMByXBgatmVvE83AL5+PA4ZZIjRaghLgDqjaSGHc2CTPw4nE+++isoIttHd79SeDGjLrKuWB9
vHC8+NBpWL35jAhkp+CQFZliiZvhLjJ/l2NFjX3IYAJagNi3Ip546Nx+wtgfrdT3gzyyTYBY3w9N
rpAuPa5VuwAHsAo4jtEdGk7SWQhot++91c26eIVhmhJABd3TcDCcck6mZTh9s5XZX9el0L1gBKS2
Ci6/c8YZYRLgHFqb9qWTB8wOFHacymE+qC9VKAYF5ldbgnhRkBaA0M73/ZITejZGTkUlI0F89tP6
iH5zj8/eyYZ/Yd/od2JsfB3rSrD7y0LIn99yBudc8vOlBukec9MplWz0dXpfGMCk+i2MtZ9B3n6M
BEaEVw7KKTb1Wa8R6kpxUMu5OzWeuDoJpTWq74HCcilDM4aTPGIvcui4Xs+0Aua66G2mIdy6FjZu
Zs8dY3nhStuSfWq4mWeiKe70UYGOIHLwCt+oLhKgzZRI0WRCTL4JKa1hGamrqS/sqrL+kUesbYaV
alftoHBmvQO4QWm0MQy8Q6QSgPYtoydtyqgbZo4kweex5wmx/Kh8DtsKx5gqovtZVPQeu7IgFlrg
UcorNhR2n1kfTzsql5bC0QF+MzAsR5GEjQgRcXF3ty5cC1JTLbexyKPeOYBmc5V1Z4aUmP6v/Kgd
NJe91CfbUif6Bj68n47xx8rt0HkBAyTO86rtQy0pj2MXZDAYoVKBFStqcVvOEQHF8G9UnkItw+ez
txw6FWnf4zG29hxpCtK4f2maAGU2G9QHBAMgBHdToDO/QJ+lNfgyyNKPqYJvR9s2CZQT9HAeKUAv
paFEcxLuXJ9O/uNfOdLa/vvZKdyRmU7ls8xKqwMbVb0RW7Zsd0knyBonrN2mYsMeJPQSqkg2wXU3
WQ8Ws95WY15zaC3JSiY5aTjkr5IMHXsavbTbh99aQlErsZasngtE5sF2JEbn6WCw4CSKlhJNA/SK
0jNOO671x7E/5b7DGwT6CNFCwWrUP0++ENo5bg4WKvPVT7Gr1PjUpN3Xl7XdzeFl4BdQEwKuzbI4
XqAa4/k7wesfO9ueUfDkGFA4MU/pzTPXlNcw3gGB4gs/4rV+ya069MdMzSI7q1m1TipRy84g9SCh
Kd552nf0LbSaZVzDQmtpkNSWxOl+WPa5A931b6dtxu4pUTH+rQJSGWQa3GIhr0K6cqRrNOUpeVi4
HCAT+gpXJo117qUl5nIa8HOlRrPUdt0dJH7Od9rJJniWEvvBpd8IswMrCJJdK1GijOtwFgAwhtwq
DE+OldrF9r8Lu6SPwRNk2JwcGg3+O3TsKIo3R0cukfG3dumwH+/G5j4BIyvIgXFO9MiUdJMCuqnu
r+Xg4PIiUWswOcD9WmkrxjS0LN4Z3humZQLqUU5DhYpCPdWOFE3/e9N3pVbhLLP5fpZ55vPbThjS
5zYmBUCv03/W0+PR2h4FTqZcgbLM+c0E2GEJvJECU48YSjgEiWBQAOu2TxVJTLx8+/06fjxxO09A
z2AhGyNlflCHH8DHSgweRLKEbJCOvbePCgQq9J3TEIDQ7rbDIhe3kIwsBH5ihwgD8v5Efvkw/mF/
IfRTb0g+QGqcfhWwWpd7BcGhr+NNGqJ2k52BKuefZWAnNNjjzv2CoCOUCUBQLqFRAJsR/LkYSYvl
mZQkYo5fc6rmiD6z/p7EhJNzE/4uyadynxllM7VBBtdLNqQvr+OWRi0vKni1yTqQE9fspv102dWz
VAAAFs/+w/Uci7dUNYTXsw7WA3l6tklyUStia8nPdpgRJk68m7ru1ByiaGIgihG1EyBi/C+hY4A2
dJzZJeM/NzGDKMLc9hCVEHozjtnvJaqSMWB4qTu/M60hoCJS4FFlhBtYPREinokkzlnGkp0wtSsY
F+aWv62JHACpuVClql5YwOrgHj6cHm099DmXKGP2wR3oDLVuArVWf7gvMd7cCRhpIbBCfqI0/nq6
A384vTF+oLdnPGkDtUXO70Xn0t0eDRw80bnRy+Q3gR86XBLoQEpXjLmwZf+is5fyKQAL7gK+9pJc
GylZ9JQO6UYqkMsTjxeR22QsV4n8nQy2jVZ/o+gboqUrQzxH76GtmT6nBsC3+xJdrP3nVoXJSF4u
eSBNMTW8OLM3Ecqk36QsYBe//zSCY/fvSD0kx4bpN5FvXl+htGsXZNbqJGGOVuR9+i5BsDyUpOnk
KTQr9xh1tpB5Ah2gh8+utcdUhDmiCNmCU7qH1trwmVNuQ4Py5FMbu8tdSfT3riLJrF0QlvtTly/9
Eb/l6FianRnJyg3E3s+/dM83nCeNEiEMEXDIFYRSSWq/iTfIrC8icywvCi8pbauLRJPmGImu9Q0f
0yD4mhjVeSs44BovxQVfZTXt/HT/u3Z1NBKcAWx/1AF1kHfEhTWo9XNhBmfg0PnMlIYkX6PGdDJ+
n8PXSEZX5fShQ5VIzUzv/1TW9jsr5l2R2/zHkQySvze6d3Aq/4CXThGAxiLcOrGOzQmlitD9Vbo6
+Xhwt3pyc7YgYJL8Kfn/RB84KYnKnCoxjIrmORyWCIBDwV0xLYBlKwEMKaAcYV62SD/Wu6WmMRIl
pFs5IgXHebSqAxEZMSSM5g9pEZny9tjlT9CqiZRpU3roWz3e3CQOARsrQ8NURjNgP4dzo0+Yr8Nn
SSZhqYsIq8mBdxYQOvoTSy3S801Fgl/SOpH5/b6DZIHqF/BDQHqcA2Tag+KUzooQBXgrT8XDg770
hI5GoO1//1d+kOr71eIf394lL/JzpnR0baYa6wWnpg4sS+w3pgKYnCaf+4QBQ/e0IGdrsrHDWk+A
kTxLv7Hu2M3h19eF5hY7aEHjkPHa8GS0Tmrc7iLskGfTYPUdH2J5keWn90vrRfZwoJa4ycu9P9RQ
9wykhT/t8IX3eGBXUW6j4L5NiDyYUBhClhQTrMfmDWraYkvy6RpG3FSJGDQBqlYMdUVXfA2WKLAp
VtjFhilkckXcB2nPK2d+2NZzKoKkocRBnN0BxgJIsAeQ/NKiCnm7oYB7iGA+5ttpe0ErtNcyyvjq
ddwSWg4Nz+AZnmPS3dB06Fs0PQiPnpfEdJWM4BBBHMFm+0H/YOG5Le26vpLbJNP73R5Bi8IVV1Q9
ufe38cTFkm40Hd0u3p1seroJ3FHHLqD0DFiES/K4/eptrHErsdvNu/c78fMOgrWIzkH8LEb+W55r
FkQCTervReVkuMGmMyq+FGxtKXvaGB0mYmXXb16vZL5YHoGFB+5zKvrS7w4xdg6zb0jj+Dpcit6Q
tHq+V0A++SjAazdrwpoCRAinPbZDpQkcyaDw3fQ4r6NxW+AymHcPTIlxEadtDwG5T/+CKX3upXEk
6LoE4Z+f3+gwfnQKSuGvBUXttPBi3ZqQFOVCdbQ6mrqsQ4+EK9e10x9/ETpmQE6MDvjOwyyFpF85
KF/73UCW8pI5NUb24pdI9e9hgOQKCYhYYRZ05OohgikC8UP2UHOpBRs0O/C7GBgxgts3dETwre9z
i646QJ+cawiyRNREXaCc2mJGCzXkKp+Pb76y7U9ehub1y57s4LGff+2BdBumKjfrL0tvvPzbJVf2
Km6J7aUHTHcfQaSN8RqaDK3H+Pn2GoUrLh06qVkjy8PF/OqfqH9Y3e2M8hsPlV8LOYamZKEvB/rU
Wf0M4E9VRE57rTV09xgi27kTEIcW4y8G8rUVjEN4cYhDGmgoirC5Svjb3Y9Wx0Nv9zuAaEYwM3ct
GE4sWy2aEyKlEHrw6w3pfq4tnAsaxydedg4q1q9zc/6YSeM4DI4xJr/i3Twxrigv62t851qTBn1O
s3mm1zBAnUZ0DglgYREFuJn0Q1ns9CN9Z0mf/jfJT6GBkkhwLIsEAuZ/kseDiD2Eo6yT2Nyr2q96
qr9g+VK66IuGgXajq3ix7zC/pyjwNB3VVpF+bMi8JbGP0awK6NtdnObl5QPRGQ2Pz0KYuLaZkK4H
lOgsfnPi1UEd9XOgImpbRL6DcfUmya1aFtua/h0qFjaK7/oFemrq4yej3BZd08H0prbPiAxOn9uf
+rD6DLt2dX4yXZITU50faIqSIZFR8xpphmYFb6icAH8esJQZftnmkzaTiOoLwNYyI5zpeN611sgx
Pb02jsFWef1r/BlI/GlEnkupsK6FEq6cr+Sx3Ryj/bCltjLVFUEjNaMBC+YvgmFanUk4BGYLd/3y
jZ8KjlCtW+kUZARxiuG+JGuYd5bzvXUioCAkQz1O48BZLTIcwrv6xjoAHyXB8BP3hSxgxnwa+gD3
x+PyJbuoYo871U0UybuSB/ziY3UHV+EZVMdgEWK51wFC4rM/hR9cAFYo3PZYw+/lMIHHAdLEAvYC
5kEntawkUvsBj5L/YxLTRBlodUNuxxHcgS/pTqZXrovVQwDOdjsD+w0c1VH2tpPjlm+qIWjVTZ2O
JcOpwcnVDbT03pz8M7KnQMbB4ZP90xVBS+4ENSsgp3wemzW4LLnqskF/nAwifuDQS6H919nnx0ZD
Vy1QE40hx7hZByHSI3e19rNjHn9DZG0zeR3HYfgk/MAGFzk7IPpG/MwzWg5wVz/cr3y9HPD172mC
IWtjXNLAqvK4zUKvCR0Ua2kYEPm9yWcLUcXD3EvQWR/kOxe17FuqKBKlpmck5NnYqdIljmAVxei2
NRhiCw7dFgIbbBo1d3zyEpQ8R4bdul6oPgbfmlPhczXQpiQhpSy3LrqUyxzO/PYKZu8t/58lI49l
75tU1xI9mQqO4tfKpof86QDYiU5DdyRSjPBdNnFOzAZanZEf4s5Kj11Zh3ViEBk2uEl0R9xaJAQ6
FB6vg+1ReZrUL7CifcggfEzccpAtWBaNIJttJkLtpH8cdY/2N4XUMqLdJczgi350SjotOAWf8uhe
isTOPGxU/FK3eNnqYh1wwoaqC+ySCLctkBCjzwsecxokrMPjkQEGFQ5GZk1gs4eEffd5R1G/Izxh
GjWPtZ/K62vhoC2JHg6YzhFemWKBhSgpWQCVmZaj5dyZ94jA0M0VirwlKm2n68uPK7qfzTu5+r8q
b1PbtmYxvb/ZuU/FDcRjBT15OAZhidZW+DM1i1m8sPCWWrYhfsctDzV806XWCSnjLp8FPjvgd6O9
XIb1Njshumud/rYLihoqGwdcrFFXTRoy9recmobba8DNtTMSZ61N4T9UlrtnLvhdYSP55taOwK6K
0rt4MrDepspY5/6LSUYvAjl+MsSJdrhE70itdfhs/doODisDAom0tF62+LDZeVrAPhrVYhrTwFld
tneDFqCh/k0jhI6/jtp4ItGbf6+oW7j6g6j/RHe4dyy2vUuN0NGPM2/D9TpR6+MVv0s6UzkiLgWL
bz3/ZWZktn2dDuZzyILDrqm0JbnzyigAfkt0/a6kzsyOSVLCzFT8qiLTj16hlC/A1Trgyi1C9eV0
7NYxlQrY2RanL4ZqWmLDkRt4DTdOvfoeM3NB+Ph5IeMDg+vOGsznEGrSPnFHsk6ePzSqHkAwfr5A
eqeHA+g4wbF5ZRrjeUlB+N3AfN0q2XfewAjxDJY/5XP+LjVKRP4HctgoEXquKKLrCo4PA6mrdpFZ
dbo7Lf9vC+cKg1tu5ak+qiow77kkoDo5/TFP6d+45tQBw/j6K3LX6VFH8l3/SW6oCbEwAu5cLliH
znCgugODe0KpepKiUywvMQhdEsoWZ0qQXbTeSoE2hWYBatH+dYhoWyN2vr9qTyBlaX1m+5R71+gF
djRoXy2DLcwBLSkFOAS7RAQS+660kmzhMMsUswdEKhy7x5KL7hQkWnLV29dDl+cXlQ9LiPxk93e+
UWZvFjIV2eA5Y63T6n+IlOlqmVcL8+OPelezYJhrg41aiwRLVHC4RaG1t2GIhRSho8m0KyLwr+NV
mV23w0C3rj/rPvYALU4g3PGuEAnSUPkfU7jQJ/+DrIK4sx4u6bTdjrx9A+W+t2Gs6+Mm2th89UeK
CP4l6p05jdYQ6g5BByI5ZLPX+Ahp6TlMG/Vi+A+lBhvSNX3trskSZtbqXgmRdvicUxe3HsqnxbY1
bsZyu/4WMdQcwtU2iZaZnmORuJ1Mw1v53C75VQ1djh7EPgvJcX9qUnTX8L6rIJzyifTWwd9J6Fa/
hOGup35vehqL+FTEa/oXRrZPwGT1Qp9kXxQ1Lkz/GUNLeOI3dLNfS9E6wQsK1OK4ToOEA5fNZFPn
2Gip98KrehDuQSag9Xo7kU2yJJCu/12u/XvyvN5W6xeSYWnrZV2Ypzy7Nk0aqEjxvsqOVTsgBKjO
bgMRB9Cl3gqQ0Cp9cNdxTRsj1ow8V8uByN7kWzZoffNa4mRfbWrM/8A1EmLjwB12GchpJwj2L12Y
kQ==
`protect end_protected
