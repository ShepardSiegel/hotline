`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fjYXcn5oUZhL/a7JVEiDS3FwGZPQiudlrdVSqCK2s74ccYsrPz3PNiGU8CurF3VB8b75sa2a/SA/
0qAxqly45g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
I5HpeJ/tjlbp8AOM9YXU41vnsOggwvQb6gwO4hVGte5JJKv+iw1kbJM9C1xFVd+bjR3UmAhRX/7A
k/mCSM4SVCht4tekVWjsn36+rQJyLzPNyOYKx1B8ZKfUJ0U0x95oKDU6on3Tt8BJap/qg1/vBE3X
bQ1w6umy3+chTrp/VG8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rTY9ON30Wwa0kg8RgZFexHBERhyetS56hS6Qtslg3mO89FZifoy9RFHeqMck6kouGBOAtAttvGfH
VIULAWmshgE6r2in3HaNOFyizQZLZjw6PqrpbT073WNQYmM7P4wPfpbbPw/2wcic7mGIWyNA42JP
ADyfqqC75BCw7XhjM5F8ovoCgg/F2IIOeAhZ6uglI5IBvJKuCAHq8i8jgDibdAHIxuNVb7ybZpY7
WnJ3FWGEeWUc/RyM/0iIc7SEQfNIJJtt9cCRXqrnKVlMYvR6YL6vrY2BdzW+RV/BoC+KBpCXW23S
g+ljTrl7F8/SL6jAn1PDzL0RPefivYM8eyjPrw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zIfdRUf6GRdfjKobkB9dXSTf7gFp7e5AXv4r9kE2dSSi0wGGpftI/jEhPgnuPtbq7Ityd1ewbW2b
njCXiFLamO4iZNLylkKSsn8kn3J1/tARUN9tg7YOGm35kwv2aUWZIBYVd6K81ZFe5mq/6fJMtF9s
fJ1bDJdpO2JmBo0MEgI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bjFWDoug05sMxZn+0aKEWxfvRCl6lrHudEbGEeJftUI7ShB6h/tfnH0OJ7W1IXmABaGZdiVFkdJz
2OWonS/+agym/AuJwJ/SceKHWW3YyokvVY/xHkEE+IdRtiGCQ8ckbn2a8LMyOw8Y8uwSL+6Laswz
oS2KjzaZX1Sxhe/lSdF0E9/HgPP4aZnBa4UDmvj6iCPLq/8jEk0bGoceed8NxsU1JzcxsFO6LYTc
EJXlvFCM/PU+ZK7NqU8gm2c9K76feuikVKmObqnacP19r+FylhP7LtlNV4j4ir07hssyiEuzRjAO
9/pgcwENOKDOOPVrRI6WkADHlHSR+wB70uZhpg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7040)
`protect data_block
fVyZrIFl8PrbLxcTXOvVUJHyEbg5Lw2LcffDuSd4yjQmjQYdZPMMLuO5eUtZj4oZblu8150VrXMV
UsqWOl3qkWZnfF90w3tvXOK0w+i7zGDqbxvKSuO3sAm5TIZWy/qLxYUAxgLz8i/5w0ebjHUAh3k+
+OZVucrX64duu/lkMmY0Zp9uerHMclkZSTUCGDTt3FVYFZ3k3socXC/kh8sACUjeyYmfXkqKEDBe
R9mYliqg+DuPDFAnjuBHOpqZVOE5udoyDfAKLes0Q1ELsCA0cispyZt6cp+zjLnIoLvPY1yTZB10
A/wclelscOM3WMZGghysUf4rWqywzmTfrl2wHEl5MEpUB4QtT5i0kEelG2GWjXKsyw1umlSbd/IR
o3PbGP0FDLoUTk/9w7HaAoOtMoHHslAfTT4GW0KH6hEGzuONFQDLNDNRCmlmre5+Zks8T4exwGMi
ccPjSxPS/F1S8eem5Oa5bjVpvRRRQeTjpJ/q4ZMS97hSCUUXHJR6H/dv+50xIbGWXl5miNAVBfep
8dNBnUCL8TVzyVjCRrP++HAC8oo/xQqyAPhC7W00ObgcDJi71TZ9PIslEsVhT/pg3NEsxnam+Unt
rof54N60Bms/MJOTUP/+mJs7kBsQuvURP3lsxmmDeBQ+QjKrkdewJO2uU7jO2ljWAa4AGNE4o9E3
sQo5vmuLiPcmfUJDAhS+ioulr2q+cvmznHW3a4uM28RCjD2accLF3i44y9wlPxvbiS+/ex66EeZv
NRvP7vRAVeQhnyOECnCQNg2j+qWWvqmdFG9qdNpDoyXhVyYjQWtUM3g6U08rrgoiX/KDYioebUVS
IWRHYzakNmXGmgv0HhF8ZfdmWRzTOdc97H7mcDOvyYvaxB3kEWsA9loYLxG7q29ACzgsymiH8Ccq
qJumSZpQ6PnpHXH5ualM4Y0PgMO8G4bIfvMnCSRmtoUsjff3Xk4KcVF7H8Sz8dNMt5nZpTdWXbj0
xBYGOC9mTjsiNS+Vr4fFRWYf3qe7u/h/9Wms7S7LSj7AbfEwJvhk0nedJWmm18G48OihUIrdkUJO
nLfMyXK2hFTM19KtJBBw2qGPt/8QHRhsRzC9ThtZuUV+3baZ72kyYNhQCOvTFnte3u014bUGOlif
nTklzJXHONVmkxOoNBL/rU5lfXmUGwR+wxRoap7Y2Om4oYGPVkY6znK2AtJMe75riK3oD9HbtpNu
Y1CbEubnUDr5OuhHNmBZxjZcHF9s+WlAGL1YaWxsOJ1fM0ssb8InlOUGLf3V5uJDZb7FpOPXrEkC
vuguHE8tysXdur09CY7VWoInNlm/fTjEsB/Q46lEMlPW6OJZUYWkmEh4/EeQph3aVn3Dv5sVlXI2
v61jG1ghTXQ4bl/7cn961GChT2W+gUnkNHRXqaEhY1Pml8j7/YjHt2NE32b17fUrbU4pNFy8eM/q
S+3nt4TcQootz49ZEoEO1TLor9kjxcy2T4ZO5f9OD0yL+zzhdA2k6VO8HHMY5iVezFP1V2M8CNQu
3VCvsMCkSLkj4yiec312fql1dyBfN/8FtC9CQx9wNcr0d7ZHFsnWXRQKME79/ZyFFeyMqf+IRZD2
48nQnghBVyZtNJ8s1GFJPkYFRe9rOLi0tzyo4QoaT7mzkK4XnZM5kaTS/g8oa2/I2AXZuAj40yTi
Uasei+Ch2UQqEKLBhQhRXfMKve9wezLsCjkksm+i4HYGWGAtvDxs5vEOT1ry8QmxdK3UmtRogS+B
kiVVnzDhWwiWKj1/JPtxHSTSOhwJItwr9prEbpTbWyG13pFdgkzTnRRbIa4RSi89rmL5UjB79Zj7
3hrLKPwDzjaMS/Y5jcMoRTurNLRcKCAywlvjSdvn77ZC4EgFBGN4xKOz0tbuUdmHhCTQOxOjLuQn
4kRgSlOneH2KzoJp55kzd0Y8BZIhQ8jQfcRqJJD6FArbZuD4aYFeoqMTxFyyIOb8RwSwl5r8M550
NNq4o/QpZT91uQHsuk4pV9H9IppXS+UbHMgCbNJPbtwChKri8nF03YHn16k+u7UaCRCPHi/pfJ44
FPa0TM+9nKoBgtynIH+PLGdBCV9QhAkIr1rsBm/UWVrwRxvu3h509bq6vU+75JUG+WkKTChZyAio
3baxshXD/Hx5tHn5NCB0kWxTwT/TtsQ2eKam0e+buxA43jrPJDPBM2OxIvDJfyd09wo/j+8P5fYh
BipOa1zol32GsTiPgl8w/0NQCK832gy7/U20XaRqF316o931PJMGB8P3dMuZO5B6fRC5nXyoVyRU
zfkcL4qEcYv9qQJrYZJYXxMONJp/G/FeB3D1kgkpzALOUgiNtFYyd9Z8A8IOTfXoKAc2RNG73JhS
4MClOGZoGI66FeqjrF4Bu7sE7hsqSRTXy6piNPD+pet87psmQ8pWalOyA5zCJX9EmTpt3Jl8q+AV
XsHheJ1rJnZuGW6wWqysep6SGuZC2vlwuFUjRBsdCEbQvW6Gi+gL9V5FOkgwopaPbS3I1/w1KRGR
FpETpujftQxcdY9EFianQNDlycLaKYx30e76Mi0NniYxEHNeUHPL53J7hmk3WJMHKq66JvpuMOxy
vE1iZdFOL1VYW9aKj4ylky+2VQgTrAIz5pe9puLIe71JzeC+bd5+T71SPLlVOBmfGZSVzFRufY9S
9bvhS1bn6+HZ6nu6VlZvNub2OEfXiWSjxEtDoD+lgYblQd9IbtoU7dnvJ+aMclAqN7ylSKD0gbwA
ukYm7uzFiYD5fLXKmpsCwqv1BhXQeFkTUuJDB3RdBzMRbkz4p7uYi66d1f/R7AdKp4iz/nNQ6fu+
alSY3Ta56aUvv34ZfeozsFEJOKgDeout/zS5BPGUmxqIBMfhO0ybnOibZp+y/G+JttVCXfALz34i
CdTObSvRu2OjiEbkkA9VTx052iNIyQIwdX2LL3YQjzO9yIibuOrGtE6LCb9pBThZ9CvXQGU4F5MV
J7GTmnvEa0VvXIkOYghpUD50KJCWMHGdp4GhnC8MgtCByA19XPj7Oi7quETcITZU3VwRe7aEDoHl
D9dxyXg1dI1G2/9DIDmoH8BBLtBsqPTGpS4At15byt0o7//xoOSRTm4bOASn47VVgvA2zC7V98RP
ZkaPONJLj8X1tzzk9uMwTYR5ko0ZI7e+Uj3mt5WO/fQRlUCqrFws6PO7+W0kb5VIXf84a7ADHZfx
HSuqP/JcOF0e9Ha9q3sI4MAYU0/ligikTtEpz0A5PYTCZTkU7g4pWPg5nhkElB/zAt6geDMJyGjL
7qO0ikrVvwaE+GPRJzhBnZNVRwFL7PQyzFAaTUsY/9MxaK7lAAVUTZ8rEWJW5/Tcbp7E6voNJOUt
8KwxIcCkys1yr7MQLKJzUU2gCYOvOWZCnW+KWvnT4zbSk0o4EMY7UN8Pmt7gCdS9RZqBiLaCVKQE
tfHh2229EKzwW6eVDbCxhNO0m6EMdPJVLcfZNKpK8suBAgP6V/irYcMlRfUaUWIV2+qHDchS+Q9C
3htPNfBASinGTl6eSBiNEHX12wj/NxGCBse2EC+F/vTtlrhyC1cMKQIfURI90WsFk/T3OOpqte62
sO/204c7HhzEwWsB1EJyt2oIzpRo+8BP9C8gd+tlJphVOfgT9TjuonMEd1T2K7WyEY7jpIQojDns
0W98iVLtJ+/E7zfwFU1IHtNKFa9mo1K3vlQCuHYmhBuITKGtYjQBQJT+aFFh8Ff/FdFogm2aV7+j
j3Fyi7tTcICXk6HrXun0d/fJp4ABbOzfJ37d3sLfnfxB/zEbjGkZrC4YDiDe2C6LMjHhESD+x/1U
KLfPhgoLjuJo8mimG3asoiNN+CGJWKRrdpb5D5BFqMnVjQcJNjf84kjI0WPW/23873PXWjvWfjpP
+py22tPxyNzsKMMo6P9ek1HfHSkx07u7hASWSlwjZ9Rrsmxw+9RMQlf8ZFzn+aOWdP707Vgyf7+T
fIGK96nLa7KSRJ4s2Wo/9G8qZ1d65w30tUSH5M+O9y/x9/984Cn0oLh3WDTC02SQeE4BBRmbxVSm
XQwLDDi5Pbrg3B9HN10p3p+34v5/gUV8vrrcJ+tsNyY2bHqWl03gYf052aKs2xS3XM0BpRcbqsmB
emNvFnYzY+msIWocrKlCXmeMZJ57inPkVfk0NKpma39HddtVHOoEsIldaY4s75rdca9uxRwmqvxt
pqHNm1A5xWvScvVxyl+SwpLPPROrOmcglxiWQXkmH753bhfPD1QgDR+uOxsrPJVHvlhyLt4xx8/e
TZs7V4H2T6UbwQEH9vO3DF6jdD0CfUgDj4iBxSIQWtnESxhQa7IlRy5LYiuMHRn0BO2mXBxG3L/P
7OzrU1HnRtJk0uOKMya1xFQ0/mrTDSKicFCukztE/+pOpZT/YgezDT8NKDqo/xdynXfy/kI0wVIA
a8C619O9/3dTe+sgkVcLjJ3YkAe440xwwZ3qANbHqhYZV/RGyvLLh42jfTDShwCBga2Klw0fMGOq
NPe5p5nk3QDcSJoadsiazHbvS6CinFNrB+GZla1BgGgloWRDOLjA3nDTyY+l/kdL15XkYh7yGi3X
QtWrIn8bfr83QmYj4sVbDiEoQN9yNNBSPf9n178WVbbzRd4nBsJD8NKXQ4hd+jJPrfd5vzsRC3za
uJIswEhnxjXaffJpCCqyCQjgOcpIsTlrfNEzbwFnqZa3sCYjY60q5HGcjZbk2jxCI9G0mTbTypoF
/TJfXgGDAq3KM8bzu/hWol3kMqAiHFqjB8xEsbzHv0peSe0LNps6VE8vDO1nXKx9DikyzHY6uVLp
ffvZcVpXsSCMKVwGvZZS08hcpEx4pmT1GGqGrNSxQPJa4HEE9epn8UjRzlz538SWnAoBLdKicekg
ubBGf8HZuyOqxoSM023GW0EnkW9mwMk97FbRs6+86YKhoPBCyp+qGHdDF8Cmg8Onee4wHeLhygqT
VB9pml5LqQrDGmfqwFgA5GrYNi+OltFezLlQCYuauaD480N4oL+PfgLcn+kPpM/csa+02Ts9XmGK
BTS39d95WdU/TLMp0sqmSGbPj3WL0s+/pPqlFeLQJNme4hnDHtksCysfdBwS3Xc8HP4aEJFkLcBH
Q8nQK0+uDLVPN5sQNE10LN3EcqZ2wLsYW0bo5BuH8cdmmoJ8oUChrdRv2I6BHSFD3heA8A10h6yZ
thi+95hGYqzV4b6mEHf01d9krVT2e1q9TgzP9rOAHDt6nFDAozssiyNIsr2NM7lUjYHCp48vtwJE
z7I5Sc4TOhempQCAO5/4fnoZTp/L6Ifm97VB6WGDE8M58mT9jjWbu9g8nu9oXlizb0GzLeQp3TnC
iruzvu2TzgWxmGLQSNjDhI1kCBpFhTmSiK0I2mw3Rvk4e5m6UqkEgfoCnEDPFTj8VaZePY0LYwLF
DTpengMi+5x3N7XUrKeNhU0tBjrQIhPU7Xd6+S1X1jtOeIA7AAidSLF8y8JbqPkAP1ytC5pGtHMW
yAGQ9Ydjj3xkPzOfhwiKPxxTvmieYUGW5Qx6fdhbfStUPG6h+44SE3+Ye628IyZoQQlLfDVJT1vT
jr9XcO6rsuqmKPHeRjfvqybuQnPvJCamr4UZRzPUXDVdS5BaHyVJ7/VQliHm4DnhhmW61Xex2qrG
t2Px/b/e9a1HZ4721Wv++dxGRcJiByFtFSlnz0Swc4+jHW7Cc3QLTn7Or12OgPjA1CujmW2iju/5
IcmB2z3dVSVnMofide0BH9NuopM6O6JqMvRDqdYv9fUL42YrW0uq6p/51FTeWCxl2GP5SKkyqnh2
nkMUK1YH/V91kuM4b/2kB6oQ+jOhIHxB7ZIghiBr5CKf+9eLUAjSpiLNzknjAzzOuGoAShczVw1f
JKL14kSItmvUpBcf4I5DQ3Ed4PXbs/EfHd6ZiTb71AjBOrWAKNxbE1/BL+jfhud/EOiIC3jbMsnA
LhJVJWzrnd754JEHXX8Or8kWBLwCQXwfLLNvq6Sex33RDtBwFgKUJ4tZ7AJBYKn/mMD3HcGBlBLZ
mKnI1jyTdAR2ui5KULENr/6zEyR/y7XRknmLp4SvIUW9wbVJNtXjdjKJok+GEhI0b4co+KZ6yLqs
74TnRvj2nA6nqhlInJnYFuSzi0gtpIfOmXgbynTxPK36bQGkzncRWqo7rIsdoqGtUceKnpE0ryUx
xeW9b+byMM2it75Pigp8I99SS1gXnELFnQxx/jtWf8j1zMWA0U1a+4diYsH00U2UA6jk4UyWerxP
tt3I1tvC6u6jCwHAhAE8I4j5mcvpGgNMYN9DbGnNyYffsgOXpYCWEkVikB/l2p+BOYahDfjinX9z
Slx282gXvui8lXmuQOkJLxrF7mswMHWK5oVIyu/9iY4LfpnPHvbzsjWejI8QepQN0Tipw9sWQoNM
KN/YTe6C+PVoLsjUij6d6y9U6eirltVKNnfehCwID4G9dMIfIRWg4W34gW5KifPwPzvq/rtrTuob
OQIAMsrC6PtPE4NMtRzcHSKvdUVVufeMlKgITsLDpo6539mKfqKLtwxbTauxlAjdj2JSuTiXrB3/
LEA66Te/Pp+QPJ1iVGqhFtdCxVPeQYueFhxGNuaMOrSuKVe5cuy2jSS/CZYPgP1V1iKv6tWzrks+
kfGHUA0u5THVvcUq1xUqx6/iCXzaAwkRUiksT6SF3NKyj0WGIUqay6ARLQvonoOjvyG9Jzgi9j7i
o0TiluyBPjNSXlDxLgLrS2cvrT++5Zeui65G0qJwDoTeGLJwHMR8PbeDgTIOtQyM6mQOli5lFhKz
mhi7QCmb7JNmr1+JSRhZgCizhnjXAVydCLocyFz+o7I5R5J7tr4gA99B1uTYgV3pbk5aT5FtXZYW
OjMTwWdDYRb0I4uSNwl6aEbG/YLzWXP1igzWQDim/bbh9BiOCNsr2yBKb0GZ1aO5hvikCk4y5v23
YKjsg3pBDY2gTHPDRqbCVbnbZDvzQY0tMYRslyHyrzKMOqPI4ellY5nxOE+KzBaMOddCbgtAV7ce
1OsXubB8eNQUE9Hf3i026yjZDnkYehQDdR/jo9W7Yya1oExtMwmuV3njsNm3xPVwA5aJgAHrI66+
Ur80vjl9aDbaBA/QZq3If4V+qdR0ZnVfpj4E3OyaFUWnFXvCq7eQe+HsZ8q3ZNbuy1Xswjf46fVI
qwzUgM2yBHW1oVHpMhXjKTr/H7SrlA8cc3Vpl08lECrmUP2peWgMUqSq79AYjYLRmZ+NhRESvIKw
Z5K5XHZ9K64F7w8Q6MDp0orIpLffVEb7mcCaqGjrQAfbJDUTz9d6hT0UCHQn5iuDt54uyZGqZmeP
KhdQ3RjiK9dRmP2PLrEo2QBGPJoKUYZXQYLtg9GbYNO/eo5TXWRfWe+oFmWpt0bbDxFlMIe9ss/y
7QI9aNWtmXO8mcAT2dr4Jzumae0Lf6/5/d/7C5ThMIdMlBlOQHWP4DXkRWv9ooLuexixOckpFDft
I2NX4C1K5bD+7qoZwdvohm7+yIWaZjqWNNuxafO6BL8OIsqTwYX9EstEWmUM20UEjA5N66O8MVFd
jeRg99NaeinAb/2HctMLrnnOArQcuB+EBULwM/ouzgZ09irm5CKuQB3yAUFcG5i4PsRSvtcqiT3A
G+91uSyFVBwuzOa3gVHB3xWAVo1CW+sJkPkcQOsEFTwHQenEa9vmEbh8Vn1osqkqaFlPGeXu4dxL
lOGIB/mG4rgeQf4UU2/CAeJX5EO9uODY8MJAQOYkYMX6uVpTJay6RWoXjkHvqzjgWSVpWJB4elWK
4acV7534bi9XbBBro21A5/s5jEMOJ7GGaj0qHIuT46NrEjeaCk5DHikvupVWaBkw6hdEPOXe2svu
gVxH3bCPJkb3gOKk0qwJWw/6G645iyGF4Fl3G9ereXcVwn8TPJLWAWF6xaOPCLHvoWqXBMJWhneB
NrBpMgFB4h4URWYKVvsyeZefL3rG/if0YhQXo1uV4mFNeVdxqu2gBzQTodbMhH0to2sDqsiHj6lH
Y6bdtdz7/AnvT9E9OYZJDkBmmEtlOI6sofL1Mwp41BiwdTnMSx0xrqYoJr4MutHxOrbStA1Rvxqc
jgf6KkKTducEkA+8sV//F0SxzMxFntdiKjBJXiMw//ybOA01b6XkWmafZzzJNtrH20XGfio0XI/D
84ctA9BHJj/AZgHqR6GAJDM0AZk5n8vXKhFgNRi6vFqEplKha4lVG6x/COvK4v4Df/sKG327M7ZP
rBhE9fXIDWojpG/lcgZD279uyG1gAtcWhkuRPmMcLOoOXIiPZkm1s55WDc04lhU0srLNRZPyu/5L
kzVA0yoRRxhigrm7hUkle4vI5SyAcLoNmI0TkErmMY8H9IFf0TRmxz6UVh4XOY/ipTuzm8hpHv1+
yMgdHUJHOpqsA3LDODWh9nEyxZDy7dEOu5timwKXni4mqWGN+WD+il4Ntw1jDB+bAk45w4ZKlraR
8NS/i2UwTrOeaYVyT+uXH/DKzYz8ELL7vDTl2VRKexTJDNc9OfcWFTZ5/eYgbsTBBAGtTVcoFl1/
0NzEbiRIOD8SYQHchb7ZFvNasFLAKvspsH9jRn3Gx2zK0h7bjoyyWpVci9z3kMvRQ/hK7lFFWE5y
4Wj2QgCF50c1xSHDBDIjOiIXf7A/GQnS+YTApuOVwISYS8VaOI8lNPMALP1mZq87yDcAohnHfsUO
NXvZ62dh0UkEQAMwTzWlbg9miVA/2+3XTfoB7mcwb5iH09p2uyqAPqpopZXjFH1FTUVpKW7V2bTf
ew85Gx4rjxU8H3FmXXDGZ+yT8OQsheApssAo0uSj2xvs/9pSzQaFMrz1xhWhYsVrlQCtKAVI8sfY
PhNaQxVwP0ue7D5fUShmhzewPpm2xmh9z9eLNkzxu4FZRHH+YR7VMICHoTAyckwVePSzsQkDRwCQ
5xSVySJGzz8LrYchl8nmurzzjS+izn+Lf3Lzs54Yrm9ZJTmzb2JKtD35Yo8hH0EpS5pKIpv8mKbZ
aOQLvUzr4aiheViSTEy2V+Re5AjfO2i3km6WVdwQbXvQOIHjBM9CkyHnVIGAypvGfi4kRXRxqmLU
3E2pJWC2VdGlmsbaq/w9fbDrkX37FtmhNm3aF7uueTHjcZbJEJPLpfLbnNk81i5wCNn7W9s59+6O
Torv9jL6Aae009QZ3c0Frznaq5QbeWImhcWmdfalfxd6+80RBUDyqScWRcuEEomhX+X74081br1u
832VWtY0YpOUgryYx6cOG31iJLIFSh4aqZd5rhs8EVrcxm/X0JZsLcjoJac000IBYp6Y0YKRTeXw
xt4xWBiJ5l2wkoGHv8eTx/z90BQQ4Y/1wYHD6AAMZ3TvbgVGjimcAJVLuSGdxhX0l/IR3W7z27mR
wH1c0S7CSHKqeCPUMB2ApVH0s91avWWQdpJn/L0=
`protect end_protected
