`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
M7f7g2PWePY/9SKLDpTSYEaU4HbSJPvhDBrf126aObPhq2yLOH9kZ0EdRmbrcrmxtglsJILSn7So
1qoDgWvctA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gRikViRPuapSPJHnjOjqSHnQyrROsapwTuzdTactmPgYPCK/EShJ8MebNUprHsUqhEnEKCBItofW
mBSAXcwWQUe2XN8I8xTe2x4/FT7TPgiGpXunvYEUl11AbvKh/BwVZ6yprAgDkliiFwwlp9jHf+bu
mUL6ZVUUAL5uw3Ll32Q=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rXI6VpvuErA4OJg/cduvdH+XaIzg3z2Rtd6P7iJBouPm32M8dNLEPQRGiIJWYYyC8MXerGybRTzk
ATaperBcmg/gyyoE04596dx/ELvQfJPwFVga8yQoQ/6AXORkuGUXktLU/0JqVFTGL/kzZm/PuqVv
5mbn1Kmai0wiIjUo3vsSCs2FvKBuh6x7CON92Z+I7WTGU+MDJhkM/kiWsm7S1QevdrCm40vp2P2H
vahY1MzIvt1fgl9dxSs4s9nwZx2kbsabGgG5tUVG+ACXguKYwT+6ytUbEspLGcP0gOW+7inDVX7M
tbvO3gFxKxdC6Cyf4CYOSwVBDBACv8ylsrHGrA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zScbT+tTWMgbgMda/zLivJKiKXmhUT+v8GKVdany0IF4BpiNqhIM3nd5XJQy9i56gj4VQ2dEvk4S
quVjleJCkSzX4NE0hl0fm2rDSfh0ta4LsA42dbsxrowui7zp3PPnpyooHh5lvoX8FVhODyBtWTUB
U4VrWDfSlwLIUIR2D+M=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CODuspE19+MMai830MbHt5d+LY32yw/TarND7jq/aR18WsVwiwAYmA6VCZimmL0FiY6X2mkYiyJe
5dGkn02GWd8ijDf06r95/8Orf3c7RVcoQBec9ZCtx9ysVrk/v5q77zHw3uY2x67LyfvDzHdcOlL8
ruAxyJ7/B90T3Oj2ZFGShJFkSZySEaYUyjLK83LkUmXx6/mc9cp7Ssm7Q5mSdC21qRSwbUQPnFQx
ZNbyQK0TOeKucmJCjV2f0Q+NvHqX3Y7o+Q4W0iVxJKwkLTAr4KKdwbwOFwu1k2CRMmzN9UPSymEI
m/WDGSV22e7nTh78N416yQL2FxhtEmiBC9OaVA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12560)
`protect data_block
10Kd4aP9N+TAoMzBxtVgyHL02r2HdSFt3gp62ddyWl/a3wuww19WmXs0N+GVraQTyxS1rRxdVqM7
kyWpCwjAnWv1MGQNnmlH5zEm59fYrL6Y+Yqn9c0ZgNaGZqH/Fxba549ZojXy94T9N2FxnH3Ek9fo
+Gkhh6lHuX1YO6B7/ksypEk9wVKK54wS/mqZWM/v4lwMyVKkKJMx+hqGrX113DEDbcMexq2YdNTQ
4NDI71LixgfvKntD9Ib0rBATRYnbbMLOZz8msmMCNG68pIucUvdck8QaW1DD3cHxhNgyrZKQBWjQ
0KRLKcEEhcqvm4TxDje8lqXrU8P1XdD0XAwV0AMQ4GSeWSXNTP+QG0pa2aN4Z7rnu5WA4nJ/uRga
yMCoOzcxi+dhqcJfOvZW6RetwPqcqR2TWw6Hlo7j32pX5Iqe0zi3se8A6+pOnQY6m5J3Var1d9H2
MGOdpx6WDvOU1Y7YFTpNzClDrKjfQQRbFzy4oNAv/6+BUacsi0+NUrBrwHra5GTzwbgRpXaorZbF
mOizQnA9YEcninEUH5Hl5T9LD7DjlRFRuXKXPdS57xwzeJ1Ivqk1V+/LUXVamyxWAw0ZmgOuKaqA
H6pXE80L/ua523YuESy7tJM5AqAUdNCkEvZH8shDUEhFeAMWfIto5kqmy3R4SQP7oN53OfOM8HwO
KeQcoFBY2bGR5KO3PgjSoC2hI0L5L23Bqv3pAEuvkxZVkWAuiV6akkEc/o+vcdIkD/r2Hh07nID4
U2y3sLpnqXRTvK6kulBJ1v6cLBRILx9U7rpUnTnbw86Y9w1WeAWW84GHXS2A0BbHOug6d3zaXMwg
lO0+ZAxPu7mu5m4tCBQFOI4nPzoWPtk16tBHZbyMOOAbqX9B8z01MvW29gusbX3Uxjpp2IwNcx6v
iBTS2qf7qDKF0G8cdlv6RFpgG/l+7JzioRtE3Xf7sV6f9ehCvQwehNFK3EXX76WmEDChGuwzyB+L
lim2C0hA2LVr+HPYGhYml8WdBXA042fTv0DPf7/VGos65mxr3TfkzfboAYMHBmvbzSACqgvCPCAS
zzLt76+34X/rBN9eSmisW8bHF1tmh7Dx7M0qEEFaRroSIJZ5w87UjvKidEoA4/MMEGDfyBPp1jd0
LViui5+aMbxzYDLz+r8HcXlkKRyUfBZH2LIFlW+izg4hPL6kTjFNy4kyY8ezYuIf0qnJzFnHj7BA
pTcr0fpsWB43xYZy85ocK0Z/t4KkypJfC94djdFF8e1dW3JRhx/4Xq2g9DSSexCePO9geR36ksZs
IMmJO0QzaTKlNOEQxe5L9Y8ItalMYDTGmFcoOwH3Px0Mt0kS7RMMFOd7cUBHBF7VVGoChENRzhU3
BUxezfEBW5DOa8JyxJQbqM2N5jIGQbDDLCmtvS2XUp/ZisBTKWjTqA6cAH6Alc9hsL6Suq9Umkzv
8Xn3LitOVUoY85sqHPSfry0kq6cyPC0WMdXUEUeaDdlNQNEzdp+4Qtm+RNZihkKYT+sPT1TxjAet
kUra2TxMir0Hs7qDDOqAkkOXPwon+esRfyTZ0v4ogLrLE/GEOGKh2sYyUF1uoNVoSu++W/hS+8/i
FLmhy9L1WNB4SCXzurk1SetJu+ZScJ3Jwn8IKzVZNZ8/EwJm0OJSFxFObywHWO+TpVPgdgPepZNc
vkhzQ8wMFyX6L+AWa6hOcCiiCmDvrjxAg9TDsCOomAjx6unqthmrYhX4iQ/Mg0eQKJmnKg4qcjjO
SoNQeQbzNuc+PNF6TR6nfhHByNViXsqemfq35AqXBK6CC3z9vnag4O1eyRIg9wbpGa9XsUK1PcEL
pSe/qFNMjoWu/J4fzegW0K3NH4Z+Fj75jrZTlkqrqIL9sHL1sK0wsVjy/0QxweKClqUfkjlMMDqO
LfC0WgABioi0DNkM58XBtYRqMA20PI6lWEzCjEi1BXallWnLrTMVDn0dm/MUcY1rWzDYFMke3I44
iIEtKkw31KrB05xOqidm89kN0cBfus5tlVtfISbs+ok4CddqgWfj7DYjoIkil7k0Vc9KPd+dX8xS
UoNwmE8Q5FbTDTPmd8waRGaYWYnqVP6/z3UkIYG87kgO14jNlGwHc9gvrbV/hXuLrnnXXUhwTw3l
d5+dsrNKgAX7RNwfhcDD7IyRGDV5dbhoKWS57+WV2q4mi5L1Wy73CnBzA5rvU/Ouj5gB9zdMdXYv
2zMVuZwgeIt/ydu0eePQ/lao9wWlGCmSTW3w7bMmAOwV/4pFBAqaYw33SgxhE1xhGZD3yptrKYDA
pPie5sjJkE8xr6N9fuzaBfGdQDfxUQbmzw665IzowTAbhGpF68FhXSZfieX9pjqZawPHRND1oPcT
gBPcSJgIAlsPiN5nERGBMuIzKW5NiB2yhMu1KkYm0+F7nnhi870FPIEtpOCnbno7ORq4z2dhhtfS
1Tdt3h0jPokWe+OhizqrpxNFsPHSEQ8gtMgKuwu970DM6RKVdnDWNg/t14a68lzwCWwqRjcjxpuE
nUGMbqC/PY/Ij1HW/h8WKAwl3566F9nhTLUSEacHMNRAnTg92LgQdacKcH432KBIgWpH/KFwYh+q
FHKif/9DZtLfnj8Ke0vjGAfdIvPuS5SbPjjSqw0dJT2PjPDZNXuCosO0Xs4elZRZbJKuGj+SdQZy
zJpLaemeNlTj5xJTxRuYo3wd04jSBzT2dKSHWXz65WfgF8U5pR4cKfnv9tmvD9TMVJU7LNZecDtz
r9Jb8327m3rbm2+45f+vTJ6ZaHEYvrUJ3xZ6QfDYtVRIEnx6PaXZCqq4QorQvdaQ/okg2sQpA0QD
yW0YoGiUoVAyoxC+Zvk0v+JgTI95a9GurmBY2Azrud591GO3HvivY8wl4tK1U6axSCsTRrlJLfKh
XWsgKDkSXMkWH8v8/nG0NSYM0FvBXfv3alpKWpEb4w+3N8QmZT0vhi5axwRpFJU6SP0FODeUBLa7
R1t4BQwOjAfA9M4AkKJ2CGKhjqWuN41Q/rpaF4KvDSMsuvwu3ZXQNLaWK4DNUPhdMRaq8UMxZSVN
p3qNoaNri7f7B00lN8YBfB7BC2bCADaU4At6iPNwZYhoeIPNfQrG50O7pFxJf1V0j2Gezf39/e/c
DePyOepvO5OSjLX32w7f1ZQDy8+jG3xb+DjNA5Kl2P3UCSe4ce5C3RvVegeNY2dzLSg2ge6n2SDq
IPIzRad9kIHfWmlB59V32EoNGPEhU/EvPt/JeHT2wrBt6HFAYatiRs/Wv6WiydK+IAaBBXOorjl9
zNsYwRMQjKF3VOaA76D7L0IW6dVk2+KrZM763XbkHymgiP9n5NcEpEHrD5QYSmXZ0cuFsPLdkn1P
ufhN17mUBI8rxuiAHjQsqtLszUD0MpC8/qINJkCsZigFhAcGFvINFjpsBGij5lSApphKvlhlJ3fe
hDUsYrwp1eVhQ1R5qLxVZJipFQQ+qKsnLWliv0AuHZeRTZjyYbuiJoyfIlBzPdCUtm/G3SLpZ0op
SP4WimGydkQ0sBVXuifRCO1afwRMpX9Gqma+MKUwU+G5fpNnaCNotCPVGpnHsueSqi2LFaYvXoLs
pRBDwllFlEZRGSKa+VV8UKd1bM+avWZdx2rmHhkie3tko6jOpmBIlmdWwgvkpgJscdDpY75BU86v
eGD9AVlfitwdTtHXXL4GM5573iiTPGBGrTtC42uX4QHHoSfptYLlTt2LSJgwF5/3/sfUc0mrl5lH
e6yyWav2KDzMURUD1+bBwdjwAFJRxnA2oy2E1LQ95jQeWvUt8OexbZJoyxCBloaFQjCbwulZAzRf
TAx+W1+MiKYZJAvyDpPXjS1jWDKC8aIqQHDolEECMxaGN7ax1aAPLj5Sf8s5la0J33cYpBZCzkGl
mVBMbklOqtmshrTvAnsMab/03uRKRcVIjqCuT9C5u/zOEBQi14YYvygehPah6pV+KIgtclx5Iv9W
C5jCTqoC1uuMU8UJOCLZ7UJlHNntZKgsccLW8nhsCMk9Ioptrdkr5Ch9LDA+N6ddRkMrugYAi5aA
SYOTgE4enz5ynTtCEcGo+2fHmwqVQQb0X09cUEueLVT7jjDjWtVyOSk/HUfZe3depXhAk6SsTnyV
7BFKaeAfkGth/4PViO+AIdAHQJblaaAxZS3pUc1Kg+JZ0rwzE0KbbLfprMK0vlQUBzwT3C1f1xNY
FTysiZOf6mz6TDi5puopcoKCwJDSTyhovT2VXFwaXoDlLXXfyj4Uz3bsR+4PGvOIgl7GfrjFxBfS
rmnoD9p1jSu/AjaNKUnoEpyzbCenaEqrP/q5k7fgIMeJHWMqFvQPb8bLKN/xk6VgsFHkaPtJjOXM
W1MPKOVCQwwrC8DVa2vwqEIkO5PbdNnUVz8DG5WOxyv2JZcQ7Ar4NvlThhIUqdavQgBhL2b/6ynH
IHbeCK8d7Em4Q/KfwGtnhWM/sTaCqKNHqmwaoszmBiZAUVmS7tawQgABxhRodjbF1rNdRR4wdDO4
olvIoVOnmwtlMNEnpRAnfXQ+JXjRs6eMmFWE6PH00+6bCetZdai20virGFRGxZ3e9r2bGJUyzLc8
5q9mDYIYFpvLLJ/v2/dH509Nz52YbIEgglut8SF9FlXGlFtZ6/Km4OQzbbbirqOIm1cDmzSEBbWN
wdtssuCSRyHNu5XCRYZy65J4Yx6rbyiBPDAONJHKDQOO9Lep1qSpNHvTjAphlDw/ttFN9+Afnji5
EoA2ZlvsMfO5CdM6ZGEGTFTyjLM0c3xKZbPN6slAnZaVq56DbiN0baRCnZ+rXNtXnY2vZMyjGCm6
FnDpdo0RViy1aCWQMKbED7RLYSRFnFRBOay4j0zmThD6MMjRJ4dRoh+EKX8oHJaeHqAvmVgNS3Mj
TCOo7NqaAFT4xLoYIRcoKXrySVjjYFJkYItRV25Y1p8Khb9UrU0Dw7DdR3JiEihLBaY4la9n20tB
pStQL0kVudvX7Jb5Y7li0Zrh4Lf8TINtlk7wKHUJL6nuJMDOgf7yQBHV+dA9EjJxusVdeLhjzho2
0lrYgebq05myIYDxdypUGBGAUV9wfntPvl/KhaC03IoH2DHV3miStOSFyyWeGJYTKR0gwbe+qOH1
dvGOKKEbCdZ0yDm1aoEc4P9+WGSyXdYFp4ikC4kAe83x20GDFmWwjkCYRncGVTp6Ueilag0Ixfrg
WsGd5SATwkhJf8T9HVygX+rAIhnvMGCvuU9ev+oUniVy/Azx0aGpce7kALs6Bn4l1+VMSIY67fXW
yye4CKlQ4sf54dYsxrp8/YvWxjeSRq4sQDrgsXNYASjaq12L0UeEErThVFneEdVvJTuLa03eZkBr
c7YPrJymwRnY2y9BHEjJvzULEKdjxaR/1tyU5CApa4PR8sxChrCA4TMDX1l+CqftcQ692dL33KEB
4GSZMqgfcxqofeW4f8e3DH5pKYrybR7bgYGOweDFKW0jy1EUhX5MJFtomi2nOhi+NNaEdTGZOcyc
G6pGhsj4hwdzTY7fVOlrirWEnwkdAhalXRr5wve6Vw9/w7boMewb/jC78ARQL7KUc0GYfScm2tL9
QfT8AdvQGzim3n2iggJvbkX5Ik+KIM847U0eNz2UjhY3QSNl+GQIgOwVSkctqcrbvRgMSCKYBsNL
LrIbAiTJo7bQFnoxkdxjteExws2DcI42ubSrmQsDlzjJlgIWfjoUA8UpZn6N8+M3N2kidk6x3oeE
4MaBSlnoF27XM0iGLikgyhJ53qX5FrdNjQrUuzmGXEWnU1GguIpbMI7bN+ylZHoFLqAKUttYwEj4
OeoizJipwDhp0lOo7pKJ0vF49vhSfkb5csOTRrbA7v0qQoy2pHLv50a2ZHiAVsgmWt6/lXMr3Oy2
Hk+28br92cq5lUszfeaKuALEMZpvfhZsmBOFeb7hSNwMJe9vyFZZ9dCHfrcN6o5113Kq9fCmjfmB
LPfqPQdPs0qee1WtOFCuMowkDkJid4SnF7z3cFcESsZ4h9STrj2jB1YsDuDMseZcVQ+03xVo4MaO
gq6lN3XRwft8/RZd99ohyt3ceQv2Jtbvw/nrsgIieE0arv90maJwX8mC602gCXQb2dotydRamYG0
KsKD2WB+j9v/4jid+kj8+C//8zGVMax8pBq8otbUCNoS8XWWOGkGrmE1gPTFtj3qFNJiD3OaNC9u
fjpf4gY5t/igJPMYDB0UcUsLOl1G8ylBGfKBGObwURJCNDTAQwOCYLIwlANyM55ylIhwAzhtMSAf
0ZItcUNApb51ZiJ6R4aq30WcJZDWtEf1iWA7EGQ2EEpbGHzA3s1W95In8pAhf/tlXG0vBWL8DgwQ
/G+v33ieJwaSU10Ml5FQRsjVsDESKvYh8qWE03m0ii7cu9aXJO4t++oHKCTFvCEPiKr8Yp8aYvQD
0ofW73zF7ofWj8Re9yg3Yo2GFWCQZaVzUoy/ZPmEc7rpB4eu/WkoyrWpQ0cs2Qre3ButOgik9h5N
GQUypSBUFWW/Uk4tppjx0tYVFoIo0DVKJAp9CCvm9ww5b3WEpP1lvWemIKoOjYgyKcD0HcWQ6Jq3
C/P6AwI9F/xJAQhLfAwpllH3yCGmFIiieq+l0ZWXg/hRGQULeDyAlU3ndgICbXWAEUrx5rAC7bOc
cE+24tRtSnuTffkiU15TacgAqOghY6znUv0+tl5cWoXUMrWm8LrEcErjjKUth7c2Eq2bp523XqQP
Kxq2CHG9EgFkH1rfszqbqxF6UocvIRYNpt7TU+MAL/Dh00REQb2aaF5TdWPN29uBEcxKgqGZFvmV
gjWuf84HcXNk8m7HZPhhz1LrvuTc5c0xvG0/R5fm8Y26qlgkbR9fS3e78eEQJELTHOZW950EmwTv
QYg4hVJlXQ1Z+FIA1kAHWUz6aY17rO81lGFRGAELRzsfgZVUSqX3qQm4nf+vlM5IYx1EK+G09aJJ
Nqcq+KPC7eI+4+FiqkoDy8kpb79L31//Zid93+Bg+KZt9uF1jBMokE7ucw22YC+nH1+2wtYcU794
PDKIB/L/BTXassDZJHGZxebkONhcgjYqA2YkX+Vi3SjN12fyOwL6moWTiTroL3VSlfaJXnhToX/F
CEC0DxfWLDbJ2kNDr60yXhw/qQWgeoB6e2jR+T25Gr8avyCMh43aN096a/zdk7au6Bh44+6e+Kcp
0gMbUAwY+Iqkw+B8C1DRApzMtBl9TXd4MNU6Qv4WOTiWeIBz9pow6IqlytkoFxLxICV9CyFgVkdV
+LKafB6HeFU63gB4l2ZSGqhQrERdxEm+kqzjKkAtNJy+0kMZVLDP+DNHhbvYzAJ1fSgQ1CkO7S6y
H0natA5if4i0nBW5tsro1zbbOhJVc1iwrZZMqEfiYD+RxnhjzCx0+Y4ZzCp0u+7rvd/71hMzQP+m
AmvNvrV4uKbI+//PPkY0YzDqEfspjfaVqT1IE6FwJDOjxSVhqeC7olzehB4kwtV+xuaytoz+YgI9
/TMeK4r28xudJtjvuYbftqaYihvKjs/cOp44WQuy4DOuF80euDSzRX4/M+kbH7M/IncOKfylpRzL
8wR/IGvWkmsKQDLFtpATrvIjh891VpLODWMml4T7ZTigWVfZizlPIJyzMh0YfZQXoLT+Vy9FiIW+
sTmpl6oj15S9Ra9amf0lnnei+B7fxeeg0Y7sE2MPRt/XcFfNLnrJFm67B3f5wiECzczUsu8IkhXr
HvuurazeYuSP2rda/Okl4yvf/d8onEGCWxIULsrOmNURH1CyYBpH1dti0EZ+iW9XUmB0N7wvzjHK
bb5eLV8cAvbOx2RxkTn2RDeg95eUCYvW57DXlQT6/HOrPHiM2Z2IquzS/aTUABd0CIrOYzA/QaKD
uC0XxA90aoZ6JIjHXzihq6tfAH+4s4/VNS1mPJs6EUadtiWPIdafQAqxJGEUztt/FT801S5SQn4D
9wzhZ60ujkH27HjqP5+8HdXjVdLg9G+2aRWRnTGwx5oXHkcXuWcxG44V91nEKVrPXFZEhdfWjT0D
VnSJwjXK9+bKhzyMfytSc8XFOKipJUzbADDwArPbnx7fb0FSUkw8WSSkkOuy8srK0JUP6gjCLfem
aQZFXp9zvEbndGBGKfB3WomtfSEodaWtBwuI32qYbQvJXjSJrEPBCqORSMmpH/oJkpB0d74DHvWk
2B3prhla8zLyrGO4LetG0z8nM+1b0wu9vXQBgajMGhpbKw2ocP7mVUbCSYAtPmp0j6lRFAXv2PZS
sQQOu0k5NRbIvzQ4HYsp0xmpl/1o7newSs8UHJt/l5CwM44ExRPcClndwqMMYLtpqXSrsHoYTskS
gEeet0LFDKQVXbVDmcZ+qBsf37MwPgh1khjSbsAbWCP+4Wm5/cKuAZ/7RQ5aOVa8+QqQoZZkA4MQ
elHGK+/XbeQyUPGu0ecChhim9bJ4I1YfanJBT9R+/b6RQawzu9USIAcCOP12iU17a579Qt7vnScz
IFpt/mvPNsO6heaTYYGEulgz71ecaOyo0deiCQC/xq+6U/eN6azCwDKXZ3XUQgiWhEwdcvgfVvNS
PnadB8+yLq9aetytVF67J28OjpcQTngN7ASGFV2cJVu81jCAbyDwq8brk/E38/bvQolRzm2KyDFV
cJrLUq03rYWyKep8kYSNTuDrxUby+epzU1vcYiTsB8QKA0ifYM2Mpx2LCDWSqE0GGmoiz/3iaL1z
VFAVdoFRQ/ipqL+cMcAkoKGClB6kX6VhO+WLNZ63rekEtAMv0iO+dw/YEOkVJQPT4WjKqMlHqrAS
qpPijc24VppY0Y1BlFUjkMHYlJzwCi2Y73WgEX/IX1m0niKd+y52UnEnr1BdW2c3s0mqKSgABYoc
N3nTm417V031mR4kMObop4oPzm+RTtsfrV+QeVsGxBFTp6PEn7080kaMdfHwKzEQInG7tM24FvRZ
7sD/sMkHyz2QxTelPnoqPsLQMaFgm5NG99BWbRLajqP4zbJdDA9yQ0BjH97kGEZoX6tC/3YRyqKD
1hamyill8RaPJJUWELe6O1D/npv1XKmt+S70Bit1dxGgYv61D2STCP6hHcLSJv0au2Stt3d1sQe2
jW/1Pp5gl7l9xxAnRHKmxVk8JqXVXjmvXa8n5RPGk5oKG4bK4VcqmB0dT3Q5xYODxIY1UNrz2+x/
mUbfjNayRXjwV37nDEnyDUrhJKwspq4VPWlXMjSSMZc1IAOM1S96WruU8ivvZXsQmu7yAF4eD1+F
3wsiaj9gsuNxJsM/Isj4m45kTSoFuZ8XZ4hb98OX3YP6oGsIedJgylr8LHCS8+t3Zid/0BAXj123
8AaA+8lNycZTanu1Z84ba6SvQ108VwmmylYTF4/WIStEwjixsmjF8CnIzsOOaIrATPnpR0XuEGsC
6KZMsDy6BGEnjDVcqWzhi3gYItZIjDiLj4Kbo/xequpwudzmQ2D4HwaqzAKmr6tEvjT+KHpnK31M
w5XZhEKv+/5Xi66juPJh2zmQBWCFYVY1eGmhxFk3b9lZLLKohrpqzdOOzexpQZiruP5fnKxzq0V2
EAgzE6aiXDCHluiKsm6OBYn0MIUYuHODSChB09CxrbJ7Q6YkNIHP3GtCQoF7qkpP93YwcQcgL2vx
6/chY9qUr9DK7UyvbgAChDeku7D2uQjYIuKWfYeWnIUEj/sf6NKOwhPAjARFVK3pyMLjnjnyaTh+
QsHz2kOCUgFX1ckOJIUxiSSLc0hfUvEa3sqx7Ru5jLF3LudAKjVIDP5ujeSQnvPOqnL2z6GUzOFF
f0R+EZPaeetL/v+IqE5m2apzGUZqrBZtFZWQ1XR7vylbSNoPE+lD4ErcCP5VCAIHwZ53tUlfP/bG
pb3Royg47e/SRIlaAEMDxlRAIeu2xGd6CW0/6dTlHHicG3SMN3fm6OOrlbmhexhi/BMTWU8evTV1
6Huxo+QIPuJFUuWu+kEzo2ifQiI/ZvZZsW2VhJnNk0s0X9kz97CQrDcKLjflhwDLacBXYOO8yMrx
W15i2Z5SiqoXGK+F8nJpSPct1dyrk2L3nOzzrdjOyr2mAD9qR5hocYYHvqxOLXkRgo3CPwU7t3e9
KLH9VMzrxS0uSrH6A9SyzIlLdXu3p+VaPxnhqdQ4AHP8XGezUAomWRkWGPSjiSyOfAS2gi6q+rpZ
FzksZYDhWBSJQqNjo0ryyxiD3p4d78kLF8cgnW10zb8M89OEmOjEFsmIDbqlBPQIxbwAUynLr8/E
LDVHIyzmuRFRc2fEHcVO/Nb+3Lc+PojoWncpi22VI2XI9r6BV7VGwPRTNelbe2P4Fn+s7mPu8Mrn
mhpy4KAQaYDmCr1R2OBzIP7rOrmbo/igtqqa+KsTCmOUycUPa0Q0Apdo+ZokznTlyt8H4+ICz0F5
H82PNPNXkcLp237VpqZDPuucoxZrjYPUTIvEpIYazeiRPQ+vX1we/YQJ7WrDpOeSEVaiyxzkc2F5
REVJvvuYbZwYTCccPoXLs/JpLMKqEAnNvfHOVOoqoNpeYuk/HCf8zrj97FEZPL/7zmqOpDCte99J
17FOgqrzdaUM9Gjc0AsUxAQMGc2JqJ37kjJoqnKEl35nZZk5FyPiDTzs8FbRd+8a/rNaZyUoNgFO
kja6k8omxpKa8SvK0np1lGjorL73MfBOMSHDafF1rNh2qOvtLYzfI5SPPmB5wlbtINLALQubR7HO
/SID/AqVSOJ7Jxa/ZaeuPkBRQTOXwPZ/yE922EhhYoLAjqKQYAozxhkEkrj4fpw6ai9LByz4+vaj
Y71TZWNCOqzPmKZsBxOVrwMgi3xDs8/iAy62y+BLgV6CBZyxmX2GsPFlmMiYwQ6sayqHdNb3R0ld
cDC4wbgULXAWW8jvL/PCpffkzJ4+lCJz913ANuJj/0b19hhAa5zrJWsydkWDrmG8ITXf263oME4O
h4UVlBJNNeQaYGcebJs/7GTowvpZZyff5uc2ymXM+fHmP0GBHfA5QBcxPTb5VHhfTjYwh/ArlVPa
z7BBTLl5IcDebLNfiQFoCuZgVSgyNLqkY1gUBpOx/DXkP9gCPWQHHtysxgQcnFCgRXnFIRJXzq/+
hKFgYgBIgWnT7FvEEXT4wrMUSUFUUVOM9MMf/mcmvtgrSzJfcl+XdRn/VMJbWh1HnRm+UrpiB9s6
nfFObEAjEuYKMHP9cYXoVTmzYuwpbWPSLYp+fRcLmVdJSFeNqIvEyq2A2/UD50o2I7dWALqNWWCx
EUzJ4eyG0BBAjgzHYXQb71/UHEIQnxKXaXcYq4l2TXi7aRdV3Pe/ZuPxXapUI+zUUP7oy5K4elxc
JqsyI9fsq2EGSS58ZMFs8JwcaXknYjuo6lIs5STW+WYFuWHUsEH0oDB+9PQgmay92dWVOTRQUXiW
UlE7VAa2vGIYCBbd41LCHYu6lfYzJ30HEOy3vK7jaJMUKnEp9MIstwDeKW+f5lqRtO0Yhjqw07IE
Xx6BEWwJq0NcR5fG6o6bs/vRb6kcip1UzOh9jgZNogzNMSwXyjPgR9Yozts2/TUOLjkz8MNoIN5u
/K1iVGCdNgPMzflGz1fFSFd0nMEGpvM6x+OQDiJTlFDtLCvxCvyhiUCRRFacBnop7g2e3q3aUJDs
uWrX7EJniwdOata7eUgtYnd7PsZWQ7pv1uBTb445DCZMDFRmiD+F48PeCV8WLn+Eqn8r0tfyOirP
n/yaBccfC8DSDwg6NTRPULpoaPaF1eZwTAhVeszcICdl2/Q2MFOyZWev3Zj/KOJoAmKRPq/e6ElL
WrSC6BumoRtUt2YPcSTQjX+WDVZxPp8qygjPKMWWJKPCqB0QmHLTAJv7hE08Wkr+W3Y3okOyPzdQ
NhWLTo5B4/TcyzMvRbz+SjgbXHxS5KES9euAo9TPwITDP74D9JjBErKXql8yHYUkH3DU1AYUUxgo
V6LzBnyGLgZoxy3QKvI9m8M4LVaSNk7Uh87WSmlbF8ykJJDhcx4yHup/IG5yzMw2vvAgXVnIwW/Q
dkNhcAQueiXyvcPsaxE+DVlkzsQpWQwHlJ0HTdYeKneQR66379hyj2jLyZWAyolFtEurFEHj23AD
6pWxc86MMiSRDktkNhU5O2t1crSrb4oIMhCvCCfhPC6g1cnxPRyBWSBBUq3mUEzbq/p1+jG80PKP
z21vrGs+G3KxqnHOsWJSHQaYJlYXTpMTFR/vCE1HG0NNfmW4i9l1JLmDFBibTFHz0tXL3OxGJJTZ
+eNYAnfwVZvulcJrI9Co/bYvemQPfPdnyJF3VaCIjxcJG7tBoRPkWj8ORFMyRdyBybR514eP0iks
K6pcvoRA85QcdyeGjTh9IGllx4Mz6Ov7OQFPOEdqwV2GY4MTVrkmK/dFlhhymaOzrP7WzGNk9vxQ
WJbQm+Q2kotyOkcF/QcCD/qRrBUuPFE7WqjmCnFrwXQD7iBTDYxlS+y3KN6ry27e+yQeEcFUXmhw
cQBBO/J+W5B2Z1nPRU8Qp7FRfKJEKoumyESAIV+XJW1HOa6zXX+ewxFH63QftLS2cq8f5kC/YxmO
A1OpAS0jsRx3HCfmo+CeK4PgZCgVemseLh2H9ByuuH+tIoxgh/GqTlFEB4xelxhU6YHJF83/iF84
8TdQMpI1v8zwEAg6qanPwq39GOaZjZC0rg+8Pob87FGOskAgL03/BSdcAP9bjlU+bKyVI71g5eO3
TGB2bzYk82Dzic878ggnicpN4P523lmjsGDy1VRUr9xxG1cxGGhnD42vF9xk6qA5DWxS4vaagTC+
mKZMTfCVPvgNFCfqPEMnQXyXNZC/AC2idRS3DLBulQDv9i+3zwl1J9G9FWjidHVLn3xd0HOI5WeU
I4bFIsLBkFDogkY+l/WJkrBDfw9OPxoYPYgL/0sOV6cNyGVuzbZ3VDVZe6bTGA4utgyrYg7o/GNr
295Nwnpm8pGeRUnVMDJMfof+LFhOkijAkEYRARouQjiBje8XxmyQzQJqOv2HYt6/hvtD11VwjxhY
qisb0rwVpKWpT+fjxOwBuYVNUKtQwyoQcBpTd865bLnnVaqvhipzSqT+qtIeYX+NZvzttVx4OL+q
JJ7CnT19giJOpk5DfcC59yYCgxv/T6uwSePIgi/GK32UkLQ3gLBL+8DTRO4JMYwe+MwokVDWosmV
BCMA8Gl1520uQ7GKqZwHVfpcovAr/GQv8LSHM2s6Jv5psJaU51LDmj1ZWEuyz8DlGffYdKlSjzcW
YiTB9wO8cKBQD8PCDxfl7sKmU0N97VDfCsQ7FbsWBBQomLN2ll/03AuDBLuyn0y/Hl/9Dkq8gtYZ
9kve/PNk0uCzsnNhniw25YzcejMCyq+CdOsxQqn05AHxOhHnxu/mnE2VcG3GlmKC6OzJAhbNi4op
tmH7OuCiBfTVXMWyeIdFD50+mkTWCFvpqxF/D0tseuWDeZvBOiGqc8yBWgeQWTRMHbAzcKGM9LoL
P1lTVU2PS+o6p34yeIsYGRf+eR0I6KlobdoD1/NCiG4h3h8H29KG1MHz3dTajgwVf7v/WGilCNL7
VBSKEHnmhD8Jd89kX8Q8K87+A1v6LRbRzB9l6HhFqW+PEJRCCrXJf/QHMkuqR5rpMAtB+AFB1t0J
1xxGmvpEnKiki8NJ+AEFL4AgaXEuMfFDRvzgs2Gs5TroWr7JStkYYE3V7i6S8McPz5AMN9Ln67+j
pDV/NI0XlZZ7j6k9TbwdDUrm0gPg00Vc9MpjgskKzqzCevf2ZKT/PVedZi4Z1/HHrrI1SLiKHl+S
hvwG6P93PrkPaPm+4bfK9QoaDc0zNJfFjL6DPxAPTR7+pMG1f0Ul/B0JfHEufnzDUP+kpmvJLpJ4
xGoi7D+AsVq2HkOqPe9vE6dQhlRjZH4c6R3czYylCBlwJWmRBfB0t67MgY3aZGeApKKlM9ff1APR
LgpbrtQo+t6W5z7a01xx8nztjNrnBOXkUel8p7v+tgZUMvi6kVXewvR3zJDKbG6ay2K0yfqIsf/y
MlSwmkdEGC5UE1V0lNqzOzzpEaK+NNFIYR++ElS42UJdM3uve3VeiG/mlukq4BlVDyZ5124A177Y
i3hAvWI2frNm9CWkB/fXUO1nyb+lXtEClG4ikeqpds203z0htcSWMS60sw8CSWczFZMW3rYYG8BV
wCBahghbj+agY3vZxn6TgJXolaWpb2g8yiLW9wUDhms2QOFVhn0ZC/o79xjTkXTAz/3V5K2e1ubK
0v3f2RkcS8sPZgKJhlMdeb79uEh7wJZd8Wbk6yQ2Hlq82eVC686IXqFFQDWXwoGC6tXmgMaZyfOA
Z4MKalSg2xcgLPChjeLA/aj7AjQfe8HmEqyOB4d9wxphI8jYedZEv32IzC9p0y6ZnLlgYu+opQPB
zElykOWEaFC9yemqIAC1PqhJHui6IAFObvQq5QaLfynbyxGXAG8dgBI6cmTeSj6uc6hHh/tLm743
Or/RznlIOs7S0ApFQiAIVjZnMrt8il8sIPr5GUn4DVotSuAa7eimNjafBZRLwxMHjh9clpkDBtkC
gwsTwE9NuNgTToEZGvWiJO0Nk58dlmSyWf88pFavUXnb7fdnQSjiryz9OUB2vcKO5sjEeo9iYuEp
9G4HRS5DiSWNzr2oLe4tRzMisadd20P31ydyLC39/iDg9v43oHEVVB38wKerg3bq4h65j4YCeYAv
7cE7p+HjG0GRhOF6P8pa3aB0+g2CcrMzLs9BycB+M8hPFBovvDQloE6Z4MWPGjTWz7y1kGYeiJAt
0fsWtNrxwSMDn875ZKmmMQqW7Q3OweeGtRaoTMtkR7zXBerolYFu65MROGZmuPXOk1LotlnvtAwy
n/zPFcUCqMvYdWXdYw6M6OYtnI1iJkihOWzE5/BgY+J1AHfaDFNqJad7qMfY7haJiWWwL1F3dGNU
48hztGV0r7ANDOvZYYSwbuLsTL12OlOIaLh+0jLIcdUsfKa3CEs3G3dQWHHt03jihL1ACXpuj33j
lC7sHfEJIyXkYSs4klIQCgfcpdZ6HViX5CpyRYLQd7xSpQ+iKr5Efw2PiKE07E4IGF5o+h8TSa8D
UpZLOFQ9BM0shtrMtwnPFzN6UOjH7ukRaPPCs9ZEqNVvvXYDbMvfgXSDHzgPCE5WSMMitIS1ccgW
SkjhQvdCbcH3l9giBH+NGEbKNQA2Y+g2cQJXY6H0k8DNLWXNLY3H2lesGDEyZ/8k0+7kzS/YeZZH
4aSTe5lrhVOvchxpEZebzPwRsXE93VnefsJWU9J7+lEFrOIx9DaZJrU1pPHEXlM5KKmWaoNdR/QN
asHYVxH+WE31s+dYkcr6q3bYHSmTRHwNWr1SXJVRLUDkmA9NoBw8RcVL6RepL8BSeduSfnTxmrBQ
90sEXvopfBKXBVL/HJwGXAO/WGUMUcllArkKeycs5h6aIVT3pD7v0zGUyHg9ghpTwNbqobpkhLFC
S582f61DlhzNKi4GVc8paTWNdF9YjTO936IPOQZy01r0L4+T6DKC8VXJPG8wqSWSGNZXefqW30GU
rFdXlO8sjzQrs1oVZs6wVd7BEHqNoUkt8YaOTcSdhNgkGq+KrhV0YzD3I8MHCjSoBcaGBbBtLSDW
wCxFSeXCbUWdxqpBJBAgg2NgZ+8mO7P4nDUKD9MSKDRypJAKsCMAd4Li6eiCdNtbgTwUz4hLLLym
0zhNWvQ7vJ6QiSGatX5qJy8hCaYedHe9KK+cjvvrnQiTaXTkxfLaEOxM97qBQQIRlZg5SeECUSed
svwGkh398HzL9jtjrOGAU5JZDfq4K8a+5MNqTz1S64JT1X6661Bld6D4KOUSXI1bMpyndjgveVEv
sZJe+ov5lbkiZfBLe+IgVXx9vSIy9pkAbKP4fBlhoc/sQJ1t8AhcbpsB84S5uHirrfwiGUNFUQdQ
V16JKNYoL5YKM1W9wKQNkNPRtK8kDHGpd7/qptNsurzyfeoWKeOjk+2DqaO6blf/v+jAQ4BF5gdC
CtLU+GkZSV4b5ni8RCg6fLSZMRsyli3oF6xPS7x8rtHo8BQ5IeWBridr1kBc9fVIsqSU7cVDY4tK
bH5UyZuqYi1V9bHzM/t2Pi9jhDMNVQFm2VROID2UribF9qSyBoMApdz6uAdCiEKq5gb/16Ro0V68
SOPzIZCHYR3Di31ZBJNZI6LXLD5bAKOxsZrv3yjufcshAvkOwtFmXrvhVincCTESULvKLGx4y1XE
7oB7TcPfkcEtYs6x1DNvyCYp8pOcUVyd+XhSEXmiLDassOYslKhqbOozLm8Fmf3NraNI2EPqbXV2
/z0+6mKSNENJI+Rjj4hagJH01MaDqGdedQqZiyR4zX0d361YUgj5mETxJsE6ag3Kk/y12xhXGSHW
XqZ/0x8A+VhQ7NAMmXBqP/+KIfOI14QGUlZE4/qqfAK9Gu8fBrPREX9NlUr8vS/7+mIS7AMm6U7L
BpK8RVtAM3pgZmdmUBRU54XNvNFx47G8Ib9Bjvq2jI0qYjvhMhzlsqGqVKPrlCmKQtGnOIyBcWbF
AUQy0W8Saa/rvBOxyM7Dc2Fnzd/b3b3nTToKOAXkJ3Mp8sgfQsSusISENkV5heSlm6wJXwh+UiuI
WLVRlOoke7KSB0Kpb0yZLfQqD/LVIRItIxRHXzS7JKnmIH9nc9IcJE7SXTz39FxH6ihgjc/Caocy
hGA0WHcWlFZ098ZlT+McvN/f0By8VvGdTDux5BqFUFaqSJMYfgzF61klWfkNLIoac9H/Mt06EHOn
pjDLVfg+YqpIpet0l29JJ/SRZ/jf5bXv4YdjL8L3FWxGBF2vFYnpjm+gBDVCAZtGHacyXKHVvpfP
e2K36V0G7PA/Wv5TwddBhsiLDLw=
`protect end_protected
