`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NB7s4mu4ZZaJUS2kL8r+M9sBaKUGSog3eBDqcoWXR8Q9+yt+xeJb/0IYAEFVHXTfhe+XzQqff5HD
wKSPdhhK+Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ofJbbZihSHWRuD1+wi+gYSohv5w6GiCBOvPofpssjn4UmIEa0YBLzbFkJM+/oRSHpxpXnYprOlqj
ZvhaYc9rOyWFCxifLvQ4UlaLFG2aZ9bCvwPPQT+4HLUtI0q+toAdTcK+bPepPJiR9lYBmxu4W7sP
F0JIuox7AhAn2u4/KLY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NgkwGaCzBVr+r/+RiPAQlOv+avrdDphr65QUDhtIZbB7Xob/uzFrSVizwB2bobpknkyyctc6Gryk
q+XJFr0OJyEzEagFpw8gISZVuOEP7uojkIEljbzPLJwEtTyM19g4pO2hoBTOI93/vS6n3eV4DMtS
dsC4IR+mBXPM0+tsSRiz6F7gNZx3fbRGqjTCN75hMXxixW9uAJkZs4qmzP50wOEO01yEgDFxMzTN
vdpJdYIriL26x/1rf/od7M/dKlc9upij4gHsRI8B1REHZ4NoSOhiJx70oF2X77+saX5gOQf9xfoE
VNZ1QIr85hLNxnnmSmja9moAfWZ1vJ128039Pw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uLHZi+C0n3JrfQYXLU+zTanGh34K3MFGL+eknVSHegPUzQ8dl2apKIQRz6TCX5+zvd0E3aDoaoFt
GOlFD0HEy/S5LMiLGuTjgw3YmZaWqvZiNB5o20XeNSyMnwf8exW2ZSWfEBqcngxWfAbJ40gnoUci
N6baEzWjpE6hJo85bI4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ea426SD4BylpswxT/O+cRRTqtbY+OnmPNRwkxOy5vwI1IOlPjnmqe5v0gWjC317hHnroCK4aE0wt
2nliyHzp6ht33x+eWFPbQI6o0cxRmgyPHre8J2pgZyIaUwhpZBxfDZgi8rKaJEsbtWZiV9pOxON1
oSzNqej5IBNwBF88qdUeW5kd1tA2C7+XlhAriifA8+cadXMeSPfzfJq6VhTyJbaaM4oZ8gotPlce
0phtIEMimDYUU2nmWusA/gHN7WKgjnGBSDGSxbxOUOQwiGW7zVH1Y8TcBBrZuPNvNnDDJZwmjoLA
f/2ISDKSB7xzqwXsBq2gevrt44eQHnOmn15bNw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5248)
`protect data_block
zOo8zd1j5qKg0fAie59dUnX7gNrvc0jDNqcjCJZ5upD3oCW48ZOM51ITLhnbGodOw/tX2H4M4lBo
guYpN/zm8USD5k0fGzl8HO4EwI2KmJgC6yKUwI+QoCbdZfk75tHtHWLUM9VNq8AVn6u4M7h1f404
ZIWRcmLY26RUvOgTkxjlieZaOMtUaxk2Q3k82IaDGhV3PgLDhKPhiLoQMqoCdXfGYqZUv7FTggSE
rumjHnkkXJ9CFgaDzz4V7qO3m2ypI+DMEv+GY0cfHj1kmxMMsKsnQ3w0Jg+MwNXLi9QEK1UoukxM
b3kZrfIss8co25XY6oryDuIeV9UV72sAu/UKv92c6KkuqihQwbrY2IkDcRhDwqmd5LuMIoYgouHh
1Zo6ziFEgA38Vg+jYO1sEeoRs93CX+bME/cdQRBYXiPUjs2fRgoXHM+rH0s+jG/+w0KKWRd6Zure
ibmBz2HszHYdBfnwS3m/WY2AnSCmO9MctD532Xuz8SM/fLxy2tsaKQk17dlpEs3rHt64Yso4SXe4
cKRPxyDfy/r+EYyrmOCvyQdjjkon8KLx81J6IAbHZZve9avX/fis3/8hZ6vOk22yloPNjHj2sGtC
yIxq16qsygLfq5zQDymEE1JSxK5XAVnGkvT7aLZqq/JSowgozWQgwdBY+3wklWVoLUuRZaxhWAcP
o3GjPFUDluP0JnxuxZlpsBBZgQ+1Of/JKe6pkDbidTlfrDAMHR1zEWAKvpRKyIXV0pSjeIYiLDsr
B22U4ezMi5ezA0z5+8eS9unKHV16wniUhxmBdPaEGLAMYdz3RGLlipRtK75+5mk3cybStlI0VZhj
1zaC/oW9+lSYTXIrHVCLzIyul0CxB+LpPULYyFYwmaB4WGukEoRm6q1Gcopy3hU4ceUIEHb694De
c+5PxgwnmSgFwez7BR9Ioenx75B471moswt70t8Sil84eB24lsvpy/+bXQ+Tp38L1RXjfsmuW9gB
2abZ7HoyqmNEA5Sym5kzSZIgnPAmuKZ8rTMgHomN+Gq63fF7YdkDgjhLbeT5EQYSwM1M5UCMKkPY
AozDI0E86AqCwe988HH8E6S3XlXnkRen58MmsmAi0L8xcBRqzeRySrDphJ3FYc7xPeSWdBK4beGM
dCNd+NHKIEVePZakxU3z6vhAhvgoYXJS/Kr3R6KliYceRfeijPeLykiEFlu+PCUbiyHQnpusBTLM
lUHr/RgvktIGWfrWSElb0Z1+LYHXzSjlj6i9DFys6nUpN0kT39KvA3Y+Bri/uZDG9WnSVU2iUKwQ
/qyDvgzdaXa32NryJoSrwAv+xuwcaASRluLG4b3+td1BIamxVdMApanr21XwxyYm24L//fpH65FJ
Zf0sDtIBuvb0u7fN2wR8TwpcTV1Km05qXLZpO0fXv6ccyFG+4xmyrcumsyBceIuRr1rKG93m6m2q
JeNes2KDFl5pzyOIdWiTnbvDZh0kEc3ZwS3cBnALiHpUyX98CRKfuDq/yfNuD7xFv07gIagmsICe
rrQQ0TsrLX1ucD4RL2Af0PX3SDVrncPOImnnFtV7oBaOOys79yNQjIKZDNbTNocienv2FlkBqdpK
hp5wZv/DQMVcS3rv05HdxNunFevtRictsQt7xcgcW9T55vjoq3NvPpE6ICePbPOzx92z0lxbf6am
MpHgYCjuHe2QYqmMjQ8IUsknesPudyqJbsmmKuErBBXvBmIyCueA7QzBPOZPzcsHrmfDlT1rre+4
JBgd/Dal3XVjziTy2EPYj7T4qPYNMZ+PPDma1B6okgNSr0j7wqek6KeCUEz1pLWgtQQywsCf6Spv
HytzXnHCs4mmANqOlb9l+Al1jxUDDLDSKERitK+2oMCVbAkZYCdWapmYWzSINbM8rxQADY4W+Tmh
9ivBbxAYQJ/XcBhxVGJKW+4VV4EI0k6OEjq1tzBiQtf5M8zcZvRWOvOTjmiooKtVzKTLXLInzyQ7
qEtu9lYmnqKxrJBi+zv7PELPd/XaYa40CuyyJ5EIX6p4fIYkAU/FOR4DtGOxpFFUXCBTeGx7Vf3P
iHtzbndlG5jhHWuZCAiJyf7GR/AggeImrh1c7/AY1XRbDBcR2yfD7pCricKbPyiSlAzZX7K0Ab3c
Bi8/zGEDc7NOoerUyZQeoK5hmm5iyZiXenjQxK1EjZHblmzm51QTKt0xVCY0YR/CFRbgg+Nj81Te
JGagBHTtPKIzfvpMbMkbY1JW0cWtjoz7q9LWTSzPO++0R/Zilyp8Ed2fj4/oV/TnqNJMAP+UadKj
C8u+N3a4VoFCM7/oV+FmA+O3nMZDyhSDcYsGow9/O1AgfrlFzed653ZsRktTAmrgyuN8YI2bMFVx
lGLdp+qT9Q76yNomdPeGQAOPrSbv6v5HpwuS3Z1eZg/moxvXXd5Sgmej4Hf12BAjouryRHvMm4w7
xLRJX92m64uDmi/MR2Y76CDWT0L3x3SKSPpKeFlYp011BiTFPJC2UE8uKN/UBXizRsbftQHzvDpX
UL3j+LnOpcxrDxZo/3Q0920DmdLEuoVfeZFuh1UPeUlL8L3Wic9A1d4IW4u4lbIK/Vb8EBr4gAT+
qS29Go4RYImRTK/+T74tvfEq5DNcUSCHWzbDVBaClmgXkw0T5hlTLddn2+LT9pwHALnnt+jHDdtL
xgTKlV2nPJgMZ69VmPMOEvnCcMGTqs1SeK3tWQNCRyNKCh6hJTP74KFxDxgE36/SkPM3iPzKubgR
SxNkvIzJdj2A94uoIr3NmePez5ymHr7J64fQ5cQmxvtii8u7anNItxZ0e1dYd3fuiJlYReHec7gm
Riq9xpDz7NzGqMRnUrLIlOWBe0WfXRJAI5NRkny1WhB13VgL5OcPX/1N457PdQshSzcPO95rW/lR
Fad9Ye8fcDCSG4d8O5hV2y9t2kO/Oit8GNHBiDo6Lp9jJ7y46CvGwm+cmU+jqZx35bOCaV1vtFKI
vr51mz2OqKBLA8FKQZWP0wNr9YR6FWF++939FKw+w4vB52A3Rx5VIIEgDXEmN9K8fDvSTH824tZ9
vfeGcSLOT7KclwLHJPRPrKXGYwNEU0I2QLXPvshEMoHK/SQcWhP4uGUYVZ+s6wqDLrnGSZS4W86m
+n51IQg7MCE97YscHXjfG+NMmAd7KuW9wGnLLU0D/kZqCIZNyPIafsQrA9VyR2NNW1Jz4ru8dt99
5cCfgaZo6Ac4+UeYSFcZc9LtylzbjCPv0J0VpkJDDprv7NgOJnfSkCRpORnKZQf+8r7G/JjFu4RO
85f2sWLc53bJy7ez1+Vuku/5orFuOeEoDrjwHmEJ7gOsd7Ogh0tQhMxUAlmCXrb8XTAEXAiiMqDd
N+oLy2RJjLmfJQMV4afU31G24Y5XpDuiDXjBwrhhMdjoKEX4R+sK8Rj8Rx0AHPbCjvonzLt9xzms
hXhpoKmkX7F9nQs/8Xk2jJe+4su3BPxHlqrqf+vFrDnluYfFj80k/bzlbHAPg4SIGWz1p+2JakzR
a4eIjtGz30cuKLEKPaHe+MydXSTj11/K5B5Tb9R+JjmCiPktCyqwKA5q9CuY3mlsDeB7ua3KXGHf
vWZzqkrRJcmCuaoS3ltYF8yu9BY1GcNQI7pMpUIJeWUkzWEYv3V2BXEuBS4RQyMBkjmop24awkjP
SqT3uA1vhlQyNW9hqas06rCqrZwI8iHyXSJoLTE6H+78xS//ecGuUXNv5t7wqBM7NCkZ6uvdrrA+
J+V8amVPMLqRw7pqKQGWis5jWy1Z+KwNr1uKfODo0kCW6X623zFj/5+3r2wsj0lkw3O9u/s8hbND
kDlWLd0tlObtIqZdxiXo+HvwrRsOXnr/76S5MVdAqCdD/LC0K+8dvdSWqBWRBZ5dNFVQUaD03edG
eGRCZ3qweyO2HQVIZh1pY9gIj+hKYHd/THwGTjh1jHv8EgBJVir7UmhxozfS9Y8i/Lci6md9L1n+
9Ns1MeGqFTqzcc3jkwb+VUR9Bcc5t09tg7NVhYWfzVvYk8vjBuRhd2Syh6ynIIc2iGx+ueWUz7Dx
+xNYerVfK5AI108E15EJML26DxXdVco3Nj5e1O5u0YGXez2g46Y62Tbo3eXOc+9Jh33E+hl564OL
Yem61KbQd7+4X1oDnhrsrDfNN9cru0AeHdVxV8+TtXThBw9KQh3bGjPtpt4j6u0cxRfNHZRsgbS1
LWQyt3QSI6Ivmln3f504+DxhdxbGXHM+ZlBXIQv2w2hUwI08KQAdS7+SayggxR6PidWNE0hLoxUp
39OUz1nePvH+PVYNNmF3szq7v1Py4O5YFh+/kHFb3Rpca/CSscVItlJtoCKce7U0MVR6NfSZ3b7B
vlaNcJAmZJFLmIkFW8jP9EX9j/ICOwu3LeAOYDM4jZDvReajc0QLXeTe7yzgunvdCCTtNlAwpiEi
rr0CochxPC5i5iHHT2GsWn7ePUoWBevCvOE3HWH9mHuwJHg67enkPxkn2aGlQe+2H96GpPg9ns5k
OtNwsaZMprBEcVPydBChcr3uWxZisVlHHKRM9OEVlrtCYbf0ih4GuTZ39Ui6JDKc/eLcyUGW5r2G
WMnEtrTxy41FBEBzYPphUnD7hYDjBKdBPjAvwiJH4wLQz7kAVukhFGpmh39VPiWHxLtP5hk/KX5M
hdnj6SLP6EsNG+cYmb10I8WsYMHOwwNCz7zyq1U5XcSlaWamDJ93hCqd98EPj63xFcGCn1JLkm7V
EkjX+sPpeYCq1KDocF1DyxY5olYkgVfJ3HIDpXvuaRRXIKzrNWdA+9sTFTfALqRFPwDST2Do59YQ
z2MeGuKdtuhpRimb5yQV3kqmt3G5Z2IFthyZ7u3mxCdufUX5VHGG2Ir3xn5y66gtBCK+H489u3pV
lnbcY+o7bCcGWOFETh2sTj08b5NFU7viQbAURWK/WjbQq3aqPYwtmNo7CAJs+ODDHt14HqAvoIob
S0IWI/5ERqE/J8yz6uMosndGu9nNtcqizufJ3x5BtUpkBNDyXTStn+mjTUi9Z0PwF2sEHI84ChvR
gc+s2E4fq4AFe4n6MQuJsWbnUBufy3ufhlx7g5KhFDPd//7DRksFJwkwJtKAB7b/LeThKgn1gfA9
RoRlFcmqTdUadX2B2RG3tSsCicV1g+v1C/iYUbs9fCtqqErvIOl3WNRc1Pej34yjjxej5ZKC5bGL
95MbeE8/SJezYu2ObroKJWshOU4FR00WbKens2V4iA4bI3aBxch2IpYV2W+OKIDscjfAHer/imrB
MatqMzZqZa3pIQmKox/eanIpyPKJiiwUFfrG0rnYNdxyqto4iJ/dUpf8vlGTY8pUOooMZB5FiJeJ
5u8pVPbZLi+aWzNei/EtLCZorK/EhIIjB7hZlWcfIwCRe/NTvO5yr1yfHluTNw76BimVXaYCpiDF
EKFX3jNTTgIHaRrqJSjaxys7RTLToqrHCmxg8U8Tb/ZWMh9XpNyEPWPTKs81WKqrmuRqlnhe2PD8
43FYnPKAWOkeWaUGD2/L7410x6P1Q1MNwgUy84S1wQiBXm0dE8kcrKHKw9Vu9mGKlMmCB2a5PDvU
hTrAQcaNVgY1gV2DlTYPkswHdjeRNVyryNRQBzrifGRCjJrZd4YrM1H+t/56Bwu4Bjk25Y+/HBEJ
EwFHF11xfbRh5TaojyeM8gLvaSCy7mvTU2mcbZIdQzxQDwJoqmhKVKuQc/lOWkNSfFrsHVLdQXMD
AB5kcfWpcbSBu/c3L+eqr85jqydiJJoOILOx4iSEPWXaUTKm8fhn3j16ykCC/+Dtrrjj1BVIJo0Z
65rrVkpqPELXB1AL7o8JzpaUQxdwC24kWknIiusw9N3bQPs8j88m3t1Q0F4/dSjhSBlnSxg3WErN
QDQecwQyNvY2nde7UIYQ0S4VjmzA5NJIn0fhOfsHvoF6mtXzQMNh94G04j4ZszQD0Mdy2B/lzyMG
h3X37oBWAGVT9GVqdjH4skexefYgaFYDc3Z30KqEMG6oh0dCFlo1Kle7Xa1FglV5UkIlubIwuG15
ZhxpMcwrWvBWE54gD4LO5oqqK61zeaEdtrjFD1PU+wI3q6cQLUVtEJ0BErQlrpynihqnJjyeAmTC
6+pJF05F907tkg37Amro1fSgVQWDBBGnIA6pH5TmGVm9csG78vKOf6pZ29H2Ts2yTAdn6ItdLYkO
00tjb26ZB06wj5wsPY0IV4v9jBrK0KTcgfo4SuZSwiaC5zH3JEM8vMRk5LjWWmLM9PqBk0RZRce0
Bphg+tcVV3mEVBmRDRLzVMTnemokYBuuq3oaccutcog/qi0Dx0I/1OfE9hRQ2HESy9YFH87uZD11
A3HCoUBa0ItGzWEaDV76AlbtEehigMeSUERcuVNpIO6o9kqNrtZ+huz3Ta1kmJyys6YmCQb06i11
ur9TGGhXdzyT3yRIkGwirqbNo6eTYkzQN2onYil8eAgfYohE7oUIjrR7XmYAKKfTvIaEWI32DGGG
uhUT0PhPDdT54nByFSOfp67H9Plthfku5NL8xBaPnSWiALVLto8GWzoWCKt4ynPsj41Ev+Mh1vjM
arWCprDDfIsmGRcLFKM+WD3CyH7vhKw28ipCFgSaAQaxs5ffuxiNleA13hiF8TUfksD8XaddrHD9
Uo0sLNCPtcji0zhKeSnouQHKWuuNF4VWRkCoEHm4h2ejPKqVuFryc97+7uJTkhu9oAEVpcyEogWk
sjhkF7g1QsA4/gLvKhMajlUzMOgoAUYpWRfapy58vmf2qkW5ZO0sSvYD3RieRfrdUvMrznZoftH3
Gb8Ou7/iermD8reYrzJ5R6eWvjwtJOzIE5+Lanz/53BZuOAmoY0fRXzslwIpajmwzLidrU9Qfj/f
gkioTiq1YyQBqU2a7/+MP+9hHTF8bUk+m+VHDqf9iumJijY/h1+aRoYjIcanxpwNXHhLZ3eRq73l
WopF706MwXEDWdZ172kCrQfAoKVRYqLtpV6fSlhKY14lg5zlu+HYwCs+tDCN1dQvOJQup9je780F
7sXjjQ==
`protect end_protected
