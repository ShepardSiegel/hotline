`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eDp7xAf5CcRdbCMmkqTpCor7vLgBVXiX6Alhbz7E68q+mG/bqYoZ8WsrF6fTwthwWNXe9afRZH1/
Wy3PalnRQg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bRPCCSfO0NN/nw1hDu2pyA/yNR7jMJz31cVDqFPol5yTBln4vVK/aFuhneJznuOzHedRxbeBb6/u
W1KZPUEcWwXM8mmBc0LhxJtREveKYg9KWb/USpsiHjJA0pmqkSdvG/e1GsRtBHNj5VEc2Z8fEB8f
ZQLxXUya1WT7T1fGPJg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kdYAi4rH0u1dF//zY9ExhucEKcq0/FrIRgZhf0mF9W57E7VJ0vaDrzDpMbiE4qtV5+H0flf03lB1
7l6s3KUSblPM2CTfuiNdv21to2utbpxeDW0eW6G9AauQTUQaQs4Rw/mgffy9Ho5qtj/7jGqvBJqG
5dNWVrtcWrpFDhHyfQVxPnDtYbIIMhPjY2qeIPmPMnLApJHZw7NdUXbflkc6AJpznCxugchYEVBS
thjUuNkuvFUi14zmw8VV+rAZwIEohg3emspfAC6rpNyB/nmssxQkA1AKt9DYD+IV/SdfeuSFb/p/
IWede4aO4Py2EiJef+aoBpw+4b/vxug9DnywVw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HgfTLetDVqx47niMu7/AvyyrFYRgysDN6RVHDqJmJV2N9innCJC/voTZMfhXk8Ia+8m2ZIG2INbf
CABPf+eS+H9ItM/eV2ZNq8d8Tiem2B3ro/2w/Prt1d+41ul3eme6/ex14TDV07y+hNTfo5PU+UbJ
aTHhT6t+OIOnwGjHdZ4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
blZHSVWXH3zjRbpLVY5Ak3JT/gRKLINPhGlY8LBfhuEkxr1o09aJRZwV5soDyBowEBDxebjjsVbO
F5Gt2V9l0c/1oqgTFXCRl/KPlLmbPj9E2O88WqfIRUsjop/elN/b4KTinugNYPDWyVZoyjBT5wIV
e4m4f41NRnJus0+Isqylg0vwFw8MS5qi7dYddo4dHBnJPS3MN32ZhIW0urwqqPQWFr3xVCQdXF61
TUSu8AP2/dp8la0j8CXgJCIJZ1MchQPR61R9axTgU4pb1rKrj+0I7e6oi3/ioNNOicAd4Lm1NnFb
VngUGcyxAPtsXWlkRc95ubjMq0n6V2uEVUW5Kg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 36928)
`protect data_block
PWE5G18EUknEoutO17TedpQe6FVGWskXkPvbxpl5xg3iAuOW2MdMcV5YkyOFKgvFxVAdd34ykc4g
RwjYD5D13e9+c/TNRtd4JO4iRIjwXLRbA8Z6teUx7bcQezIimAlVYKkUqheAdcvAWTYlA+uznsK4
MkKCbMwPKMFhIJIDwZGJvITRlLjJoAoM0GFxdtjCxvrxd8gfYop1AA2rwLaiA7PZ4w/0DNmeU3+h
FgvOGOcsZ80vqyIk0Eaa8NdgmNuNbMUREsjQZhMZF4zDCF7d0ha4tabcVG6cXl9ON2abYevS1wc/
1G8FlTNKECabgVtfDDFLTMyDIAbloM+Ayis6vcsrvYg0KtBCqLbALSBiCoS9PgDxZS2CwUK5RV1B
aAX8qKocUECWkOXt5hJMDcUARftDOwnrvngEKPlLtxpMmI+jb/WJ/JEpg+NO0ir/QmvnCH5deqq7
COn3m45Q9a6dMUFPAdn4kSJdjx5D3ZeBTKCTXOez5DiA8GZIsxyy7VAjs0M7c7xX/nnrgB2j8KV4
+pmVRSqiaIKMH1t0EXMzmVwrGYiaqgYuh3k3wcVbggG94Nvx8omw/ZLUHmlM1iT/ajkUy/77Fnwh
dqo5jwE9yg4V7fEtWoRTvF0Uek5cOKZLl4IqLa6ND1EJbV+/24bd/2+SkeWH8NQhtu1k7e4c8qms
OpxGxxEqf45l58JxfqQUqM+arvAm3bDI+nY5Ttn/gErSr+REAZupUzWmk0yNJsw+LY2wSW8oTszz
+kU1Jwfq/lWwhIMxB9F88WTDW31nmYPKh8XB0gAA000BN3BvKvD3Zbeh8milQ9G1WZNPrjaQOzhP
OXc/0xlo0a5nE+9sqZRFB3cCJ6t7Kxz2kDRcKy0tbOONFxEgnRGuY1rXhdt25BVCnpsFCiAJ2mwv
n5BJAuWiiII3veJCQFBR41g3TrX5A4+NFhn8onPrcwQGOKPk5/AI0nStnT80lNJz4LlHmrxBzqqe
trlEByKwbye7S0Bo7vF5vLjAbrV2Me/UAh0Gb8xvS69ccIPDdqvxS4wSZSA32JeD5cUI832aLeIt
DBuwCdJUC+MHesTgRVuYUr4qYWOHC7xuRIXY08QkxPJYYTja5rg0Q8b8ATavHEbQOGBpL+kGkFHq
Hg5xkidyJu4yIkKyi+wKWT2w2tWyLo8rLnUgZOrOxu6OJ/ZKIWVNJ4AZYPJSfYVlbfJ+QsMJ/Imw
3G30Lt5zCbf621Y3pX4rNSxnDyFREE/3yRrm2v8XmPPKouTEm9t1zZmOHHYrTAcENkv4P6/xxAo0
9XpvEpSbZrLTSvTlJppcklFNllg1jQ8LTYeGZpO8pR3sy5/VDCQ1gpHJhWU5gSuaOlMsPfp44ZzA
CvGw8yudvC3KK8NpSVToQ0KW6EL8JBKI86c08Q4qEAYQzmt7kfwh/T/AQB7h7mCLO571i7ne0BfS
0r4q/KVLoytz7g0saODLeYuVJObgfH2u+oouzEXkqPejRrBOTi8F2xClZh4QKFrGAEKy6/LzNoIJ
MaxKGd2I6lQqvHybAveeDvYKC1gk0iflue+gxqLKxYH4B4FxcwUFfbnB5z1yuwlmm76oOj0/AomC
HJLdZFG0LRWd4av89Zz0UPQZ/RYGKVlAOoE4Q0+7xqDFTGqCiOf4PeFqKJvAN+tQfCPmLpzoimPd
RAd6/tMYx9oBYnSq+ER0TjCFVhlQGfhrsD6jRsm96jOblYCSE8Jbbnt9i9keod4uNtOx96DDS5iK
uMiIpOYaTBa/UWuul9uiJhQVUjtVPPjLLMAwrI4XhMiLCvcm07FXKg9ofCRTTC9Qj0oFjlWzROI3
59rwp/RDQP9D/r1J+9dBJxIiuRIvCqcUYa9GoBzZV3aXnraAUUKz+bN7DGpWqp7NBRg5AkrPduZ6
v0LGysFqyqE18ah1p5cPACGD3mYwASsESSF2U0XCc5G+BbAs/x4FBUcErlAs6KB0LTqymB1zIuPv
XZnjkKjaBOR5WpDW2+6mx4BaBKAps4SRuBFU5nFEoouFozvi/cxRrt8pY+F9x1Zzf0NxcMTmKmTj
tju00/jM4vun213/2vejxFRRmtzc0fjPEBuxoH5nNf3JKVFzoegvgzU5+hTLDJ3IlFRbzLovVegA
yZ9e32cZ371ZZGsa2CwLpN4BVcu46BreDU2h2lmKzhq6K4OvOxqCuh+ikZfyFxCMZoLTizKm4efB
pQ0WWj5A9rpaTs7zPA2x+NI4qMtieXp+uKPJMKnrRtVBSIQs/XlGso2nesZQg+PomAIUI1VHk03T
2+Q0iNbHyeupXoTkPersROly53e2V6ZtPd7sg3ojR4sh3KFwrAc7y9BFgLH0drCXGLr83OhVjo3y
t8LBtvrwI89YudLMDFht0cc1bIcPjs8UN59gF1JbMcMHAAS7pPkCDNTRp6WYXrzv8aXdScHXlxJd
Lt1iXB5DdC5TwR6FV5XG8NCWjOdqfeIppSrEZD7Q+wGhY8erbxkINZ7XPCI/TXZh9dLtcb76gDcG
J0H0qZGzF6a11AmtwrqiqYguurO5ewlRmhjiOxg/WxtozRNnXZpMMMM8HO8gnZYGPPIlwOf1qYTm
D/xQrFifMLPUU3AEK+TEgGEbZz7lFMhif4YTVoOYmKZZGpPxofeFtv+Nsj3293sPU88G6MmfndP0
mUKYQULpaGUxUPmTt/vlPLu3WEgM3am2i3xDQzl5Z8tUYzZdfgNxf6XeKTkc3qQb/4GvdlPIPXKF
eaM/4Yu2NPR0y/ORn/zToHUtcTvZPozsfdZmFLYoTkXV3nNrwT/vBc8Xr5vBLyC9fM4GnQGBtsmv
BcKpyZcA9lW3urngIy6o4AGZWTWRlNvYR/QVptwKTy92+wKTJQBAFvi/J32esbxahUF61w+LQF51
jbwaXstXIbWmbe4Jdkn/9Xfn+QrwTW9BGIbYJhMt4NcKZWDrT+TDvVcBPQi5v9y0x6AINGycojeN
EV7jOtVp4gdBN9V0+Q056ETfZPIPtuqePojv9Y8VSNBYuj8XhW/eHwLeAtqDJXCQS/+nTnjj4M6V
cVk+5x9TATOcCzan+AYThhWfPVXiHiXVeCGm336WvXDqq+5RlRgBpkTQ0dkXuujnLPAv1yEQYcFE
uMwZ2a+I1RP1FME0YO3r2/rczZ6pEYe/iqxFLr8/fEq7lHY72LaBUzamln9eGHfqQ9lCRPdAbl9o
CRYyppocgr6XrVZRXdcyATnyA8cI13jRqJbEf3RRxssEBVll1euz/1WQg8ZsOdqZ6/gW5u4RLtAD
C2RzsTyHwoZO0CFNvGdlhG53PpK5vPXq27ygduuTlHBy1I2p+wtoXpU5FkCeakbP+UMYNHaEFKPb
K+WTdSOGli2So4ZQzaCH9Ojivq4nBut4GorjXZGwYo46kTHgWfDaYCPUjF/ODedlKIAl7odKeObm
XgFEKzU9zLp6GAwcxebm5sggW8ehp48dYmkMznO9sfen4Y9vZXSGXlQf0VyjLYNiSUNNSyRRrBfJ
JKjkRK+GCtXbHlx8p5eDTcCLUNJdsdVJ/OU7bV4pUAA3Y9DYrNUqfgoN0YZbRumesN309uoxixpv
7BREKrmeXYxcCm3wBgTdA3Kg0H6UmG9igVuG+xi772IJ6Wv3/1Zlg/mziuGet3QHb+OT/HzG1sSX
ve3g1Mr9moENVsfvDbpUlhzAEi06lodJuk7yIa1eRpTc4TtF99MPPMoosO317tPPEqTaEItQM9ER
bdbhXzbQ3igBOeES0fpCXaoUovUnKwl5F/79pNfhpd03Q5SQ4AL4ws87hOrrgsM5sghHzAesbIvP
DDKjMruH1YPl1cZHFwrHY2DsxloVOB48ihSnq6mUsbTX4SDTWNBAWgbtC0Ks6fwydTbKLFl75uvc
NZ3kRUTdFPwCrzUmz+Pgj9vajP1aLqVWh2tF7y25YUKLHy1LJoB2CQiMLYBvvYLzr/zizp4qYb+q
Z3Kz3bWPZ9YWHi+oCxozr5Lmx8vZt01uB/YKYcuWGzaWHsfbiGMEoWxVhAt4auPat8lSn7lfuqKO
qtxe3aV+/+oGSSeb3Jro4qNe8/sq92RMkGnBTKJ2ImFn+548sosd1L+t6hmHYPHOA3gNee4S5HQh
2/MaKRBhNDXNzGJJd/dRrNlwOVzAsMo9BFqFDWi6oontoR5TcGm0gkmArZjscpvBxV4H5Jtw+IFu
Ui6irWr7nLKeli/W+ECeSzU+SEf/cWVTJC6TUAo+cJHDIDDKSo18e0nyFxPbRSAX/dIKdSQxY3RT
0m1ZWV1YPS3xETaGt/Kjf1Ho1/RW7U6IaX6ukS+P8nv9SPWbGUxjTWd4Cbq7G7R6ifiza/c724Y1
ZTYIl+v7x8wakYrNZW+5EUmVI10UGd9tAVmAz/vtsxqcdQZnG+oAYAzupJ3ogxepbWQRWlO/y0Tb
2rTXWJe21CG7NYUg33JDhWsfrp8mKZcm3OWDlqQpnYhO9A9QDiofcPOc11iHmXQP/vymBKbt0y8z
OzyG6XH491vlP0+CHPEkHunppaxWHd9eVjxN6YQsdWwKn6TiICPpmk+CFAt2ebsvWBi18RBK6ySp
h/oCQLvV0Iknvkk9kYPOogD16T6MrN3Y5oJAp7XfIsXgngJF3w2ERCNVLJsikxS5quXBtvhNL3tL
lQaqvxyZ0SU+gmQ5m51FjWTu1yj22rLFyodR7wLzFANObxQZlVbhld9CuIOFye8dRoEdYFqH58SD
CIG/r6BGZOLR0fiUR+UTfvXFnirBoC835BgEcfZRmHSJqwmXOrjtLscfI/ZaTIvCVFnZFW7GkYyS
baJVm0i6u/JOydeaYGaAfe46/cR2CcfTbqwM7DeU3bNRucDNC5CuoS3a4C+txGsVJG7e/Huh72q8
4VOHA9NkVRf0Y83aF0P7kKZEYmNpi+0+AeqvRDTHcOf6zHOqdKap0kI7mlEbId0Qpav7rRKGM93j
aPrLcdh7O/TgLTTlcOcsH38yrXi7O65yBgPQD1Koaje9TkroSZxP69UbyXO8o79pz5rgRybz034/
L5BowxYPlETJBeSmbe+Gvryb0ksdtlXJWuj8zRuLmGVtjhu8aEIj/3TiUdMQB0wKMSlw+FXeOkoy
a9UVWMMxeQoQId8E5iIre1fOE/XaJ/qSnsY96AjZjlHwVdulWux+rgP3mgatiXPcZW2bI+I3Pdqc
Yno4eriEBgImZZEI5BX8WCCoRPAzi24irPkJOjRoIhWoMxmHHis8lr5zBATzG7Mf8jA41fQHut5n
FlSsO9+QkCNTN4N6BgVet6lYi2MVBt30PPYPuC74rpZLnXlOeS42TRQ8HhMbQnZv40lIJjcPm3D8
eNx14P+osFOZflWm1UXms+Nvp3zJ8WviPfzBa25w5bxomTiYUj8L5DYpQxiX/OAn3Fumo7Eh/dxt
u9vZE7Xxs4c9UiJbnCcbsy8/rckrfwDvbOqrdwdynkIJNCeAmZJ3VhH0T/aowAS/t5c/PQW5Hsfp
uHzWsr1UInHTl7L2rUXqVD3Hgw1TcUYI8wQeU55xUNUS4VXFYY9ox4hr4SIkNeRMaEjpcSDhDdYS
BIx4lJ0YlsrEG28wZPl9amra6m4JG9+Cpb0XB5qkUae46Uc+8dlnsCAy2dWTTU1JBK9AxHukCX1y
fb8P9atVaykixCbBis2R+e7tCttXxwYE9iQsjsg6yXwxwk2VpyioaPiJMsTYioX8OyXsIyytEtKF
DxexmZfr6qfEOPPwaoSvskBMCQPMaE1yqbgkgS/bJ967lygVKVeKGzktplFlyT3okycsQZTzqNAl
YEmR3C3MPhcs2dtUTpi79uXjbS7q8hsNtGauIydBks+vnQ3EzggtwB3D+l7iVRn2yYGWQBFEjAnD
AHWvG7HbYotmMcIvmr1IdDoOi+4zXt842IIXZkUsRSfhiyBHPYn+NhryUwkF2Im6lxIEmYC1gSF8
dGO0odeWbbeqzzrJANnkJ1f8ilCymjCVqHuJtuTMNUB6uu26ehbPonnKSmH/TzpBLpU4nvqXhBs6
27vSRShxSBPoKTmRLF9y3uMxfTMU3luh1GNy1+9IXFJYPLrhg9U48lcWp60Vc+bRuHYyev87dren
ap9VvZzPGbl49NvJ7EEGRDEA4Eeokx2Gvj/wyueeAGx+JekAaiFIuvi2sa6rcOiVozURLX5ewfHz
IhWSteFokmv0eo8DsPg+gbcThkjZ8TxPnhPo0Oa0nIOVYWPnOOvj0yaOZmGq23lBcrWRB8jLAb2k
aNOoTULWWip0sLQeRPNSlGqQP1f5n6uMxbqPA6QBw3itJE8/91y7RsSGUd4CaAeW4rH5t6N8jzFt
EbaCQnBeO35T2WOHHxoSCrsYpZNzq5JeNtY4aR4qUcRKMxgAJLUW3Jvokl3BzuPGiuyxkMUimod4
GeMX0s+zpt5MyLrzopvkTSHaysbp+5zVx7ZJvkYlpKzL/C0MjWyvHl1xHLJ7S210H+pgEJ0zSyLS
WCiA0/ivEwmmPzkppteDSwLk1WIVA5iBBzTgT6VFzxJDdOVxeZe7OcPW+yhJAeKFhJKwaOEUee8v
F5QjtigpbFu7kPpIa9TS4N4ZDVAPcGv6W8ZmF0n/Ve2bItipgmLhDfXcEpEj1wOouDDqWjr7sRdf
Elyk4JLyKhwV1SngOLSCDUnAHb7nl5St2HdOg2bg2WDZa1GcNi3IppFNGdLu/l3o0EGk6GEzc8AN
LsEbcMHQa6UlJGtOJjatfeSCpHWyR0jvNNNmxn55PoeEHvjzi4PS1Ng/wLz80yFvDOtHKhmdcIFc
wJYT3CUgY2aWiJmzsuqkeKzym/eplwGCy6824mVKfHTpi8lM5jbUReeQ3nfBFfDBcX1lYwJMzklA
21BsSJB0akPXhK2A3X3AntfdUUZD5YalvuUMJTJD+RrgTEBeeCzrRR7kIkki8JrZq2edJ7JrzORK
J8yktuLH3jZXpB02aqfTn4cWnBps/Ipp6PP0FUuS0PyURyUU+0CV7Yh/6aV3dkQ9plMaSJi/kRj0
NFdBTIBKsbI/ZbTi3vLn+pw9h0GIGj/Yj8CDdxKL9qFvibnwAJ2PoOLIcuqrEUM49j8JXItLPa0V
KgD0hPGCCU7uUiEjh1Q43Vko1r2fxX+3S56qLV9fc3akFnGY++9vw1OlVJVY+6j1kX+ziL64DEzP
aRLzpRX4wP6lF2GSHRnYngjXQfovV3V6p87K2mNySGfKeoX+b+DzVyWzXkJ3HKaJqq8BIuzKht2V
HpxJSRV4lNNmpqAH8my/vQRB+wEj/2B8B8gPKz4PA4GXogAUoGWZFAamNhdNTi3gBNi3agJfna1l
hPikuiG36HDNRmWamasFEJSuZsyzWYKqWui7o1GrFFB52vWWXSCqokrcvCVRI0xAmf9b90LCqtua
tiDmHXm9xZ0NcZkqX8dPjodN7CCqC48c8fbi2ny8ufpeK63N5fyZZV5rwl7xEsA/xgZWk1abrz2E
NIWrsyQFXTlAZaw4w47VZSeFaTlnlueFhKA9hQJXMMiupGcu4liHT45AUNzX/2ti+Ki1lbj/VuQy
ulseoNZj/uyEX3euT1euzQmbTcfAgHoXglFp2wYh/sD5PbawJtYvBP5S2M6p1dd0rI6C5lh2aETa
O9GHtvnVVHym9ieJL8D7r73+QyYD7gTMavzHC4iUhhDkyDzY9KJ2Yy1+z4FlGJ1lu5xSsV1tPoNG
W0Uom4/+2wACsksv26zB9lzgkI/qlXqO3X50cxuUJNO7Fd/UcoeInKG6xcv1OpmXbjteo6OSAupb
7msQnr8XjGQMPCOeSecrsxjqFDkCA6KqiLsBoPUMp/cv4o/kZcvoaQ75yRxmvPri2JbqR4o4WpyZ
51ImOFVkz+IRYNwkO8h/jm5PqYQGC7D72Sufq+CL0FJjguIWkN+Qh7veirHvRqCLh3J9v4xS1Qg8
Hf7R27fp+DpM0EkxWgtYBXgTyppYXdHlchU5OnJj1e3647mi7gAdzFkI+2NpPo8LoUQ9bnUVn8Ob
gRp7WUN8V2vMELCostG+RRCFNoFwlIxaIfgQUnkfIksgnVDQPzlzOYIYkwVutVE36qSbzPCnqay+
uR/dNvy9fCnnRhn4LE/WywxqCfkDOu/D7iXNCg+yJG1zV9XCwX3rJZCauNX7AdCbWxBe86hSxCaa
Lg0I+sj7Wwyac3BLgXzVQxiHIDkNbdKEJXyj6HSVgQl2X4AAH+90aJxsIMGkQCpMZRmwIUseVSkq
5cIImCACl6Gotygxf+jYv/eGlwYJduqOeGJGqbvvPYfqLVH+gafjFTGKBHL1eVfE+FaHUCssrwMM
fasgRK1i+O9l6h4bum+8+1B0GbtosEXSy5w7Ma2EHUelsvx2MkYefdC5+Fvf79I+fQdwGNXnNxeZ
+S0b3YJz94PqmFxerUVS3dRMPoasmqmFZ+3l/5PkU2HtjI8pTmJ1MG5ufktGhKzzDsb9NeJ3T9Vp
R34M6JgU2OMwxZlQFplilDN9nK9adPMlUF1P9ukcjt2QZZYeq4HTJ+GK/VvhMIB3eNlkOM9uBwQn
8h0r7vEb9+cCqF9zxSPQObLvKE5eDQP3MzHSZou+Lq5N2D2iGraeHcz3xXf3vPCFM+iuGXnIN7FF
/Iw977dOAtjrBsA+9u8WflEVzrUQ8xNyccR4qo35Jrf4iy09kS01KfxvP+3HS9A6v6o8LWIxRBPv
J3DyAN/otlxBJumoFSkE4Wh7S6WSKvXewpqfubRt+ZEMHa+xxM8fSb6ld2EcVgBg+pjFslzsjVto
cdocIKMzgiXl/ipiBmE5edhSq24Mg+WGBooURrbKbFunzs/fh5QkienWq6qi7V7TwMhpod74Pvl/
UmXA9WvpNAAmrOhZRLyMy9CSpNejBDyiEHmbzEv8T80cP7YMwbwScH0hb8DjcNwtILaZTdp0pWFx
T5UxRIg6Yyj06oYVOjlwu6Fp8/GfVIBuECH+tOSzrutTLUG2hoHrf1itEX7Z2kZ9FPAc/lgiOQMf
TqGzP+Rs97tT276J0R+xomorlDzqgj+4LYI8i0MQvLurbBIB49xLQoMU/Qewr2X/plWutVQZGA1A
MFdIIwQkngQJto+RQVUmY/YrkSZx15MremZ1XBus8xLuRHE9o2lFwK7hWgLqvF4eGFzDdZij6X/Y
UauqYsV+bVSev2/oWOIaZnw1Jh4gx3Nq4xo0DPptKOtKOGCnsGcsCyDVmmyF3xQ1Rpbpgk4re40d
gyUrFSHBVW7IjcJj9MUMCt9+iZs/SU3564sUnZAjx5rGDoeIDxK5B7HgkReuFD2hZa9Q+9s7gDUe
QkDm58pgqECfwbRMVfa5F7kGO8gdlEC6h3rtttoaHdV/6uW98R/Q8uPu4VxE/J3u/pX6n2l3gddV
6SDdPgInN1VZla8uoM2qv03oUOMayeA0zfLxEa4zJIMVJv3qZBzJ9mk6J9Euqf0+zEEVKxK5wl7q
4j2sAWRWaTSuvM2guv+Q1pVkeb5/PSD6aU+JKtx5ZOZjHhiIchAnnTZkXzLQiMxMsITr+j9cUfW4
4ZHPNxrQNHZ+XqKo5pXWr+Jpl0FUMF9eZwXpgjIqLjz1tNYpmmW3AUejk0xIf04NhNIBWomqRNZA
6gQNPY8zzqTjYhbYi93MCDawW0fRkvqKo/XofxIrAxg5K/60KrtwPps60iXup/sA09wPJi3pKjTp
n7reVExn4Ukrky494bl/jE5UgtVETdRzILeUUIlUYw2nQ9GijZcqmdD50H5gsDqZ7G7XenBIdEqj
4muxOv8Vj0ImKEzmdDcepF8+APCWjUD+twK6DpMZRtDVtSoaVyOSrwBEdRVVFQBsAakHKA9rl3Fw
+xaGsgiCxaCPfs20gBO0XQbsYj5qZlTS+3XXw26QoyTlRs4A6ZrEQBcD0fo74QPra3CvYymgy6ey
D9x6KahE+OVap9TIatULd78/cEtB65n+sMlJu00nNiiQlUUhE2V0DuUnWbfXtVlfVoiVOLak3ThX
i0aECgXM1SA1CvRt6cjwDuavLlE3JEl90xL5aCy74WEo/OezvtG8QTzJjpWDV8uQ8evNPiixLxWb
seUYtUgLz26Arvyif2FoGajbHPYTHBD3IRy43l5KkMOIpfleZtqVJcr3bpxPdARx7LssWG17HQ5p
tgRZHHD5+2XVZBCdX2It77QJxWK/JlvY2ZBS+A0cyAkqnqvWKXi0wgAz54hjpLqDx7pxut6wlnmZ
k5PwH97RmnA4z/98j08NIKuwJog+zVtVs5SXUYdgr993eSKbFDRYpg9fT9hCrcT4EByqJ36BXw6L
1WAiV3U1kvFsbO9i5kZskRT5Akbc8sDsmrL5eKS39S0ZnDY1FE+4z5UKrtYYOKB8Odoyvuumd3/m
ssEWy3G7iiKM1KPX8sHgcYPnbNMfDcIF5iV6Ngn+yq/phFxESkG2oI+2XOYAi8m/Nx+CQzrjOcJ9
dpmvtokgnDd1x/sH1Azr+WuV11xlHRNHfAGcPuCMmZs8uKSdtte1NKUOIV1oXi7H8II+NqBh5KTT
/Twr3vX7K1kqdAesMu8qC6lCfvSwCCS1vj0jJL04NFWzdSB5/OvPU8xnqPIQJTWkIM/9xkvvVGRW
BZ5AT2k6Utevta7G25NpHsBLwDL+mO3UrzJkUgp2/Eu+Ruh6Hh5xuX3R+O4+KANip03nfNeyDJXE
eolvzjkN5lLvUhEuKBtKuFgWHvBrMJo1O/FqeNLSNvpqmZsPaW7iTkBFiFZgnkn+/ZzufIl0e+WC
Eiy2JIodyE+LOveQ23CUFle/zeAvkBLO48ZLzMdQ0x7B2yI9myKZ29NQi4vTFwXMAlWe3VSV3oDB
oM8KwJdEtrw8vnv9n0avOqlmpD4gp1UBmwhSU0Qs0xQSC6tctvV34yrvl/p9BWNe5hydDfKEe9Et
fm11IFfEJyAMqElepPwCnAWhANds44AMgFgppUeKKbJPCH2XjfiSpdKyJvdu69Z62FubgBh1u+tt
Fbh8B+m3xawUFqs6teiVXjFaXcnoSF6WYbfcKIX7jh3O5K+QwtVPJf5uRuwigjN2YQXVpeIiehD9
vTAGPrAhUuLzkmPL9yxtVA92g6JgDAMqD/9PMX0RmkJBDKjiZhl6CaLsSi4nv8h+p1BuOZCyWHPZ
4l6JPUKCYYZeUysiMlFuqSPpenqOtCH8nTYwn/CcT3y9sD9ckvP8rul31NXecrZY/7dsYKaHfpPO
r5cBSEtm9I6I00AWs9v+h/1CeNoheEmfxW1rAXhP3X3OwxMj/BIzTKooVMXse0yZIlHXSwXWpaoX
2tsQ4qL5G7i+3ySF3lfwWmd7Dop6jmlaZLpN3Tl5pWHvIPMYFvoYClybAmictY4gAkrHX/zmimKS
xY4u3vgGL6KcvkO4gOVEwg2urRCFrfx74WvrErPEa7Owf3/sJFPh53+rD36dRI5NgRaQhVypbsvQ
YmXqAxb5HIt7+1yiqARLiFCbxqp+9Qdgg0AzZqoUAugtnp7JUgrrDa+bt9cweMOCzVTaBfvL5+Bd
bf9lqjBLsmS+3pjTFAJrW2iJq1C9pxJwQxKx0MrR8gogX6rX5PvGU+o4jqEpwJK/XQiSdpqnxD4F
Zlt2MtFXg9sFUU2StQlrpcDpvrrqG0OygkNi9MB/9MyO/dyxmw7Ev3WnpC0XcI47gQa3mm7UnFgJ
LieBx+SU9Av955qT8zUi0umj5LO2NRRFUwwYmdOKbHNyHl6dx0oneIeQzndNm4EZFmm8oW18DPt5
JANONXz3Q2Zb8DD4KIAc/PW6e2MKmXM2xIWnA2M5xmXUDRZ2nF979qYNcTV0PPrKYd2QUOcDe9IP
NzHjomAEUjiY5asdHFfm0qYCXlwp0lUG194bdu8hDOHyw3hK+JFKLHlnUJ4Aiikix7phjDrbgjAI
hIsoueX1eKYzw3nnNkyMlMfP080iFyI1wJHYo3Clss24uIP4kEiBEoxU+ztX68GTpXAuEr5jix3l
Fh1b2U0veiu+e2w87oN6dCSXl/oXwdEYhbPvS3dcftNjKiU25ypZCuTamUaCxCejrMLp8Aw0g2xK
4YnWJtxJKWSB/lPod91u1QpMzFhmpAgrDOPPAr+PXJw4xV8SE+aeRAeOONAaaB/v3WkAaPitvcdr
h3mj65aTwugS+WrwgTqU55aZwlHnZit4/djl7A2MP+6MT4XGIwGfbdT+FQGeZvhMWJQiPFFjqkdJ
gT6rJ8hiCcysY8I7/tcjrtUNcHbTyDbBdcj2UfHnDa8aHIqGFnq+JP+Raw+Oyr70/mYPgJhj38uW
G8gERnWjVsCxpTlPc/PDqACnMAae+uyihhoTh/Gb0QcUoQQzQU7E838a4Piv0GgiMG3PbkFin+2V
vVZ139ghOUB8NLyLPzWEEBp90elz+a6N03ETmnLLu3M6n4YGwGJs8TWbTgc8YjlvZt74fpDE0Na3
RHtIxIVIe2/63AcPO+D1SuW8ePQjXDXoCPGvMcVJxYSB6ZJOZTklYG7BTXsTGjZ6PVP1s+gFtv88
lIRnUPM594y/Hzg6b4VVUTpZc0OMiUBbJp2rV48Q3Ht6VkW2CmQ1ONgt5N5o7u+OiAIdZAQv2aD2
PlgNH19AEtBAYIU9+R/HZeAz1lDnP3EY3IMqfju7l2GkrSVgWhOx25OOl/TYsCXUk49XeFgOu6oa
cFLN+0o41cAv5MPbaYyzTE/8OxEshOxG/N9j1VJw9HKUhy8sfPqv5TXsEt89bfvZcYbUlBnQlTgQ
KXAWOvIf1ub/yKkH4KWZIMHFewMrMRZbhHWIB9T3G/o7HgCuMiQBcXsi9s5N51KOfMY/KKl73NU8
YOd0D3l5DwEsBtGx2p1DSOy0b6OYnAArv7BkuG/IkSzDapHqkBUK8O4HasKGn0N+7xaYSePkgRK4
FJ/+GU/CHwzYgVGCqaFqUZYB7P/Kkyci/OV1jrDAEGgkyAYRSddp+2lPQwcynniheOrqw0ECTKU0
Qs76d13+/kj9Cd5tGfK5XROumQIGSfca+iZeYx6MLFN+Y+V9mMoB2f0XDA0Hu9ztLiZJhVPgVRjq
SRvMeiAMf0FUHq0Xr4cT8QFmTFarMJrMTi7gleEiogcSSLQQJfKirnjkJP/cqcunFR/e1aIc7GGY
OWTTHkzS//fAlDBRq4Ho50zdiAFds2wzZu8A3phkPAwPWGFD82iO/cjrpqeRlkRZbBrhsN4pvvq8
ZqYujvQod23SmEoqnF+xV7ci2xYk383karpTxwUUPyTSAAKiMQ9r8IFzEr0/+oQPmnWNK1Q8j74U
25YJCdQfd+1j+YmcN5SOcFf8gVdcdwwJ6egzf9bwp0rcsOA4KzO6uGsd6MUWSdeZs5dOR0vjxNlV
JFHfzVp2iaEfOjN988BaonM5WhCrbNe630suGONqhYJgGmpAKiyloJ8xHDz0pRgc75wl26WIrM6K
wzbUazu0EuvTG/Cv2jjOpFfEmSOFPvltWKvNYMoHreYKPuzf4YucQUC6hGyZls9FdDLqEkRWn+En
ysxximQBJCbVMdKrQ7koq8pzaHE5hGmCTPzVVlQsA7/O3YAPOcB2JDDT9Bcdl7XWrwM/BgiNxUsv
NEc2yaX+vKKYjabSyX/ZVq2nPUS9Vk9o8BPqzAlYF29znCkq5+H/PRjBQloBH918aBi0dHH96Dif
3rDuClRJLVKSNwh+ZVEJCZObEk3BQpFJks2NW2b8ftT7wmsjzhn6gL34PByVe2DHVGCLr/sLqXc6
jLlQjKOHPppRr6Yw94n5TQwg2hI7YkbAiVDz3GDI6isnCFSMXzpVaRHXVpNodTvz+3PKo2btcR6F
7bcHC+V+omrEG/wcQ/vA7Nlxu1qgHPnNWaA6qtLJ0vfdSTYSP2cw754txpuwXZTv3lsE7yhlDOar
k3vbK7VzOG4i0RsNlZzz+Ta5gRPtE210NHtjyTW3DpKThScLnDFcIrdbh1sakwcTKtmBhietbXNo
lzIxboGdqvc+zxZN4mW2914QlXstCQfrNrVQy7el+T9M4zsgl9RtQb/A6K4n9zUBu1iYLSczOwfm
izXPo1bS6AhXNA035GnJrl6NIEhXO92LTrQvz80E0PLGIRf5Tt/UA9E9MWwDox98RqV7+n9EP+ZB
FBZwJa3pnth7OJL5iuoOHddm25xxqeR2tCPrAoIWd66UPEjVZZSYTzyyr2wAk5nr5OHuD2iABr9f
wHqyne2od1Kg6ESelweJg66tJb+TqPRrF28K4megQTuxa63cRDPt1RYLCZ2aipA5ecpoSMi9yovH
Xn2dzK/aGJfwy6Q6UFfc3FbA7s0FrR2UWi0d/X3zhzENAMPdyzvoPRCQ1dqdNmMj8kgOmC9bBw1J
VFfJz5kgfr5Vw6JKlX2pzRSKmC7sSsCv0n6rhtxbdXtIgvWtFD+YwUbh4noQfNcsWYSYtdPbuVjG
rWOUHG50Kai7/m/r6c7z3pR5cxxB6hNv4jmQjpXYCOYHY6oxz3w3Ut/B0hWogKf7ZdoOUiJ9FTIA
2NebGDWimm3srSwknq3ZoC/GwXB1DNC9Rp+5rvclgobifCqKTPBQn1I4U99LC7dW66yzd/ZGt/4l
eOAneKIrg/f+WlvgU7GdK1iH6K74c8Ghn98Ppt7uMhtzt5cOauxKaCe9loC9vSHyzMRblLmBtiMA
dJx9ksqoEPBa3lrG0OUoxSzKz2lXCDCeD86KWiqgNbgdEfdBByqe3zpwYvrRYjp1bx6VyhkRYaZx
vIYLH6nLxvCPF+oss7RBlbk+G9z00WBq3UQgTM6G6O60d+XJ+mV80q8EhLgYIh/ijhfezsojP0Wh
eJutwdQ2BdTaLcptJ0V1YArOeghD5bbEwCh656vOJdzTkzOiV2Kq9uCgybHAXAKSdZLQbfJdhe/X
bxRzu3a3l5qaDNpOioiOR8RNCWXwFICiVJrBtG+wdwIaOQ/N2douZyUESlgG/2BGOKsir5W1pCJC
RMOMsflj+39DZo69sWADyHCgGqIuCPWB0A8WvEL4nFxEot+kPNPHgLGZkOBzaS9IhAAPOKA2AWQ0
uNtIiCgEHdS4MmeUIHBXU1JJbq0FSOAOWj87upxawDHY0mU/5+raiIPuJDmKBu0KlLH2c9qGSUH0
u8YuSlNMzhsMgrPEETuz1+krFJvvUT6YKy928kj73htBXHl9oSU2OxQqy1hF6gLfBllxRUwigsca
uwBH3Ai3nuI5/iGzcgDizL7fi2NKcnfoDq3+t4O5ssO/cukwGpBGZof1e2qn1lFYZ/hzOpB/Tn9B
gnNuR/ygjtkyGRK3zRLM3pnPoXV1137vGY+v9ginWMpGDnqDUAVqh/HnM2xbj1XXJeiAKV8rTVkH
Ef//gMc03mzbnN+Pru9FhV0YUC60Nzw3CH/QFfF8IgBQ5mDMOZ0FDcGJGlSzmwU3tpehjLcqOCtS
wcHtvSdXbUzr08jjkC1cXdbc5CT2sJ6w1Hp+0kA+IQI3EEM4irOymbo17zaU02yulHh60VR63DlW
FkVwEwd6R4N0wAFok2HQlZqHP8+C4SXyP14/MV9c58H5vWYqShqqfVJ/TBhPdfdAodMH1gqdZcXc
QTl/j9BV9zM/SMex2oJ1gImzGq9W8o5Q8xfUCZbTMl2dqaeFZoowm6zt7wnE9VYXWJdKf16Vh3GM
3hEr3lA8+SVKpCPQi81oJ0IPUyNnp4H34jo85uAvCOPbeRIe84S8cKHuL2kixDzc7AjY6sz0H9VJ
KIFGPDeJPBq8xXY14pIzeR2JPaxAW4xbPiYhhk/LtJ5ltCQva2uAA4CbcewS2TPw7fUnBaifAlQ8
1G3FevErmhhBL5S0UswXFZeJ7mKl2ckfZLyUVmhKZcuekLYvsjUlmlyHe3mv+VAuoGq4goABbTkS
0kBoYzAqK33e3IFQU4fdzDnKDWYugaqJLbmZPQ1Do48xlvopojKLRfV7hXCKonQFml3g0KLlOEIa
cdp1oWUQfCgubDwdvtkkCofqQB+UlQImj3x2uRQGmbhCMJGJ2ui/qWCh6nhQzc+vGKzx02i1ihSD
WBUR4L7Lwk7IJc6LdR198CCpp0NHW9XsjgHNWBTcaCvUe+buvQIpV0gFIleYYwM0JrA9ZbcOIa0H
9+dZYEuz8hY53x7GvIZii0aqxqkuxb4jiKNTwnvbtaXPlpf2jdt3stJ3N3B7P2RRQYQVadgV1lhW
LW56o6eEIpagu5RjVHrUZ1BbJwiNeP3R7TN4c7Mg0SYlxpl3xPR8k9gYEmNBqtI3jo5AzdzpWA+Q
Um4/peBxeb4MMaAKR/O+Cbyk8FxB77oUEufAIqzarcho/u4ThBoGi84L1K3tLnaYi5hDcaaOE9Ko
S6+IH5kFT5kV2hseITa2PC0B6Fp0qbZqkTT/sYyXmYLRsWUbahHKM/+S4YKhse7boHTJIpMw7NOo
4RH+n5qGPz664NUiTxwpGIyhieca9s9hYvS0zHOaLLF8Z7431O5BzxLCRLnjqQYLVBD/0cRmE4hf
u7ne7BPEdSYYuRERPGVZqcwZ4R09br6bYqeF4ztz/8gmoEPMKb2EdwY1ZKS8jU12WaO9AsbtcK+g
tFImk9cYgFuckY8C2SZzz2+0Ld8V9z+yTy5jFCTlBmUFmEdLQdRoUWwru6CHQRvmAtsLqU51vof+
rDVbxEF6fkqKPnoMF4Z14H+CcJ8f7IvbFqDWW8aXcIbdAS3OPFjM4gNel44YJEbBSlgnrbFp9sw3
ZFKkCJNF3WTETPaPMLs5z7RCp12wtCTCqPDQkVzXQKgdbl5dvogkvvKtpzjsWdq8ulZj8eKaZaHG
liJ0n/Wh2m1/J79QMvHCE+0S61XGKGtWTXjXeM4vkch6imbU+TxBc0KJ0MPn3hHmf8IWI0LoR8Of
9oRUC4MeLdcj/USWMXm6QE9Pbz5E/LRZIeUxV/dkNbKj1iTZA5iKJG+Gyyxtdg8sn32NXAVtc1GK
3XeXC2G9XggycTb8/AWbUB8Qz1sY2IeJKtMRnCYmN9/ra0enar1H+0LL04PMmrgNdGf2aakUJiSb
/Odali2Rlw5x6NRGFtgamConaqh2jj3OYxBQ2JuA1SJsR1Q0CvZlXR6YBdd+3lDoM30tdjYp4UUG
iKTH6413VS/98EzOjv4Go/5pxTAPu2NUo+5PnQ0+YTNQXLQLgX+En+74DZeWU/rW68cxBeo4Uwf4
+hySHbExiYyVrTl63VbTj4nMReXQeBtehev2IVyU0MYaFPjHQHQQoM3XKIgw9u30JUHPZsXKUcgp
kvnvThTxEjDsIWSjbKUb4bgXURSX5AYlqh7E6IJBaSoEUbHjfgqQz/uDJmcI6xxbVli2OKbh9mwl
uG+XVBk1Kc9GNNjdkudnQwYKB4KGmk6xrTfujdMeIfSIhEB5BaY/G1OzWEzdB3tBj0ftnHQm5P7+
oIfcti4fLR5oaDPkpJpYLrwjanyrhZm7ttsM/fGUIYoAwrbdMoKgiX/t4B2fBUAcao/zb7ZPyvu7
l122DIiEkphNIXsFnEW8b2fikxIgNilQH3Vef7iH+MuH68i07ZTLCta2rl191hU9L0lwC02zZ1L1
R1EPxnwdlFifeBk7XIhqHDTl99tETApwSrvK3VxtST7+GqpsPpfTmFHKhqn4z1uqP/HRH2IZG0Tw
Gl7ceJNyxUWGRHg5recTE2YtHPh7PvaTVfCVfrenwSUbpme9Xlrqq9d2W3/POxSQFYvq1hrCjqHj
Ng/YL8ApWA+LU7ZnNJ2j5LO4f4ZlSIbsBrwpxa7QHMjv8THpVoKGIMQHI4+apNnfsE/5XUe8X42a
ZiCjSSIGDsBQvi56+vHyU4FfE8kfrR8ah9aQrlju9ttIl+W+N/ZPWsClZ2WlSYYsJvHaIFhUlx/l
UJes2f8BXUndOtinLQMtl8Tj8mOJlddIyL6plX5wZtVWQmlt7jYNEg5CRl5EqnwYv7WwJf9NEvUo
1cyI5UCpxhPdyQnfyMvSzEgJ/mjgZql38x6M2KvbK+Y9Jjd9OGzoVc/SEvCsSLnBI3QjR0wGhypT
RIWFZdtdQLetzcWoN1F4Fq715ohfNt4zj5HCGhHHNZCPacfXgC6U5T+VhpccmMEh9URtzZbEEmZt
IKlF1YOQcL6ykl2Lc3dTUVJ+tl/mXH705Q4zip3PE2GpOUCpSqOz62Ja5lYZjn1so9LFOz5gdCkD
b681pz2H+siNU11VORw36lWnBD1ofoaJuQ0qzVw5dDJjw+mXGf8pVMr0LvnYOlkBm+B28mRUtfpl
iKpnzmqxg+JYPYMzGurcAvX5qPxxU9XlqcqfQXwg3+XYen+AwtmhO6cw4cFzcWhFPvPQJuqZz9/L
4e7cjDAnvPd/j1bRQLZm0kCs9LZstFRGY+WRDNjezRBnwnKaQp4FFwHhX/TKY+kYa7PxK1Av97dk
1QeoTlmo+xihMK0KdKmSjUiWyBp2prVYg14VX2siVIJ/WVbs4r+k00uxmQ3iMIJE6stFS49309oH
/L5Hss6jUNJPdOZcsBw9OJJ5ZuTxuMnMEuuD5SpoIROxxlL9ZmTjJlzIZMp9S4lUjAttpzNpTA7y
U5mm6qk7wo9jH76PyBYI3Yh5bKb9G14Y9OZycx6oDuVWRw72765aYHx0uFGnq0O8pnBzswpxkHdL
4HN3ZphKEM76tCc2HaK6+uz47P8jsyjg2LdAfCxOCTzrlmfiSLvaLzbzWN9TMIlsBhv1juPH3uQ6
/FqIidn6XFHuQRB7Bm3heUHcSojO6/Qe7NqMaP2m/1LQgi+JqrllNuWy0dLqfyvmie1MrvJC5dMy
JHyibO9DYI+P4DToQDyF9nLX4LNkX+bJ/Ci98aSorwXfvneIYt6evoI9xGEzBitqw928vSxgUIi3
RwYsmUoXmKVqKUb4oWwMc0dX8xmR4oZHu1MgDanwOrcgPIe/4q5Gr3jHhSDSqSTyoJ9LN/wzDiDH
dF0jeKU/+w2ot+m3QD/6M4y4KupCAiiIdw7+33/wc2RTTxLYZ68Qa1iQVHfrSHW5BcSKAck9P9ou
GMngd8jNQ1Gbo7So7hGvs7hTVvWUTSbpObRwnGGFNj8NNBL6hNq6fJKHhXAGW4Qg/h6k7aFYSHEx
WLnpey2Yop/1a9obRDLLBuC/HLx1r8peH2m4l+3ZHxEi1Jvb3NmvWP1Fbuhy2NDmgQhLjco+DB0/
mWug933yeO/UXkCOup2lGJhlezVrmW6AV4tSDOe+upoDb2+f/I7ptkElOHwT1WkhEAFxgKlIoEfN
5NguaYf5QVzx/Ig6Efjc9A1QgNckEfQfZItBC1d+WYfIQX+4c90Vk4GFmYJbFh0q+4268V21dhWh
SxnSf1dE8ub0i2rbso2Wc47ukRXCCXPmA0M1nVoGqbuwwfc4yogBihSS1TmoQsyZGd9uYnyvSQ9s
VLGvtJZUGdko1J89+d1DBQsuPd/+3lF8Kbyvi5Jfsbq8LTR/hIf6rYZxAVXCetbuZ2KAZgTatD4i
Z2uUtXCqFi3fO2brqtT8VVICEHWAOK+RilS7IRzE2lQcZLR2EKA39kPMPhgWx/pqlrKEQr2BXylI
t++KEbE+CkTzMyCPE+XY4wHcGmHgtL/NGbZ6Vin9ocWMUNr33xCDIr8Ur1coQsVSjqaasY3aTzHO
0LOukdAB1SERr4rSFsjJUlmO7Nu2lydAkD7xcIacm/dvWr9Hb4Ra/BRMA9FW+l9d+0K1xHvaEg+6
2WUikl7BHLS1VA2+RheTUU7kALpNhjXesuM4irxNDa0o2rxS5sZxuw8VS1LfYC1Isb78uuHw1hwn
TJDoyJXGmcYvYVXmP3H5T9YEcc++Us2PC4W10Do31C1r3BKXGs8Df7SvZ2u9/AaRI9jtPYdgDFuZ
1oOoooQ7gAEErAUXMi+KB7QKhAtPLt6YNxlV2jzBLG2v1Bpswx3Jeyj5PDZBzrgo3r0dt1gCuWPx
4we4wL5idBSJ4GYjqKq1p0IR9CqX3i6KfVAu2nMyt7H2tqrmOxrR/b783UEzr9XqVfyCeNFNcAmc
/eIag6QBDZHT/lXgqjJYeqcXaUfnJhbfAFkLlbyDiX/6STBRkpok3RlW/HD6yg/K/tlsAMI3qZ4F
5W2KwtJWbfk2LnqQ5fU7cND1ZGqlz+KrOOiI4w6wCZuKVPzS0dwup6TfRSyag4uZPFMIdcR1PUHI
KXgbJTx9teUdHgs4kPaNUfxaZAKQyUDDR8MR+PyfBJB5xpWZhvZhkS86faGrirtkuvxAU17TzTVL
U0vfFzYQVKTk0y0caNU0Uc/QUS9X26Wml32vZTxeeGwR7H1g/LXffs1/cS8xgWttT5lS2fUVt6FR
z5NQynJRPJEq891im96qwRzWfDEqf4emdgOCmyBhC91pmxhU5LVxG9r/sRR8hjcMI0KJZAfSSHn7
v17E8RcocIUPs5+/PoRhFj5nb/qh9FU+iQhugi0kUoteYut2AIRBbXiamBbTESLO3dtHDHzVIz2F
/qMpzXey1DBUlDzJgYhtR5x48/2vy1aZ1MFx4ID0UCMVQNCI7BWsSADbA+U+5nvvb+4vGv4PNSi6
CFRvhygzZ595nQ0nF/LeGx3JKc37yQizfoCsoknewr9vOK/U3f53393c6994FVXeE1X1UBAeBIh8
aSi454nX0Kl7PqyZ2VzKim8gf+tNYQ0uyr8Gu39MnVUhea5TqBJwMCN3Ot/B5axmljA5pO19Nx82
mXBI/aBytFsMr36eLQzcWNakBHOau5qKrZYPHW6VLwNHDk8uR/1QdQ924ZtC9rCTtaTxA3mrr+ET
XZZ6rsEgyH6ZXfjRWr/zbbR6JLLmPYQrFCcsk3x8037w8sqBKaIbk61ksZ4SlQHwA1WKBcK/C6KU
u2SD843CztGArLRPEMB7jHJyMYTcKfNT/HKqzNRTJ223O8mA4mC9QlZ9/FvaqIMPWLYBALshEGiR
nfKZBfEjCPWuy6LNRHTU603Grswl+JTmLqdFA98IE4Aq7PzVTLejP3HrMN+zfoOc5zJsT3PDKhgc
pzW2pD6811oUZLcurKimnMc5tF9gM9HSVBn18nZ53uIn7U3pLH3eSkUQkPxtKIJf8qqqGqrzZB64
Fnfp+87vtIAz6Ttpu9AxJLmavuFye/W5dQdJU7eWw4Mwtcpw1Cw+Qcdvks/EYtzNWgtcBJWyO2oZ
SI8APJZ6n46O2llXG+ZMRsn1jQ7ic/9WezaupnUH0+3JHEDEw2fvYbiLiSlI6OEsuajPBscu7r6Z
Jkmickhxzks6uE80fGfccvikSPHcpnEQrLTB86hSOf8zg0ME34eYl/3kXcyzfxMqg1U1CV1c00vq
HzGrYHOpKNpe59ofYhjNkb1SGbyufiGrQDXzNtOBsnm2lOQ4R2Hdc4BlWOm39xG4tQXv9vjvWT8E
nJpJy/QvvyvJuDTAOAYWKexEX1LK1Xgq94hP5xzghv/kpFxnv+4o2l6S6NACzxOgFTy5LDJJ/Med
7dIQwZ2q5T7TztkgctSO44RNy5DoXUBPskhyzEuv4VwNH0ZtNz8OMYgCmgk0R3KVoF24RkFhSAQ+
8GVEFcDr88357nAgffrYLDxvQWWZLv76KMRUnucenJabQaOq+CIWDEJf/2N9JLLomYb9sM25rGjv
nZU12RUuLod3kZSlydVq3qKQqvHCT2xp7CuA4Koqp+7UeHDW/nP7hY5iO+EUauj72SOsvKobUzo3
7mAdfhxGeUYxDwfle/DaPGqXFH+gLc574lDTIM/m3gyKIvIewXp4kaLsRj+Nv3B26vLM8IxgfexE
34FB86ncllr3mOdJvSCRa5bcVZIzD6AsRiwmss/LnkQfZwalCFCNK8qHetP93USfiYrFdyzo1Q8C
M1iOj4ktFeOyO3XfZfrkpDh8XdiksZR2A/df5eEU6p/sBSYfzwes1dhfcUOEpLm+V2xxaNKexh+U
A0ls4pwn82jkkmcCxbW0A9aXrXeBlyosr4hZxKKVqunt9kxkKiKoxn1lnjwRSzuyv3Z0Exn4i7ep
XyIuYacgl7ySR17apE7C03+XaPkP/qavFV2WJBDWfL1ptL/1Hh5mCLU+9HkXg4VmO+/CH90N+MM/
QtmR0cPO/JwlpP/xFgcZLs02XoQoWl+1tfxOKknRB8BqZBuCeHhaup+PDLWPhGKk2HAgS9WD+Csw
eEZgF7qY9Pjjg4xcQ95lxSdglHqEjOb4bq/5O2u8ucDOdYD+zNr1J9nJ7ke0996TlB5jCZQlBjob
213Xtjd4t9Yce39VaUvaQIg/gS28UFm2hJ3hoXccXdx+dKYAwPfCWG7Zd6ZaZxRwQuIDGsZz3d/I
8MYFsVWXCkDTOZZRsN0XymQvXxT/OhsRsiu0z+UTnEwmUE51ppO1CWxKEIaqSviTU402O1rQdLMl
2ATM0nOrhNBvsv1D0MACQxwP+km33HqC9ckZPzUQ4H7l0PqSUszZuxpXDbH2UOvoTCFN7UWCKzbq
QXaNxmHaSBQmQ3gCZQH7dCN65u3w/ECHfqnczMi2Pa6HSuXO59xSAYrFR00pvxdd4oau1bNCd1RY
4nFyJd8IPujCRFianjimYDeN7R0E/JIfUjdJg81Q5p4y9w874R+WdYfWVtEI4kcAeq8Ftqy3syI2
O1ifb3scZF7ZajU+0oTWk/7Bz4U3hAZ3IJC0lmsqCoreGxl+4puMFtdrb2AvAUCOwGVnWKjLw7Gb
wa7whJsMLWgrunYNJfi+jWCai0m2KtmL4SDCmuh0ZiVhhI/ffJAWGI6I0S+u8bsjuAqHS6qihsw8
TgK2K7nujmd/FFRiFOkVboCrtC/UKOm+FrQQQbL5AKfQ39lAeeDnpHOBM3rN3ThlVNb2I4weuHrR
DEQJYvIY/E8okmqALabx4qMVT46cwJ8fLm6WSbZSHelFK9KCWfWbqhpzZ571n0VGIEAnT7r289pR
9nqFN/YPnkh/yHfxE6PlMArybWnN88RW2mHi6OP3os5/hF8APoTdYFHr7hx3W/OXWuOQy0PK77mY
052WzxdOaYJc0B6fivXk/32DPGN235TSDNDmUz9c6tHMhEuhW5WAQUya+XjIs+SRyvHqLFF260a6
4elsVxqfc0SRC9rjT9RXbTvu8tWd7JUlvMU0SOuX621+r1Y/ZH8R9+vYij3QnGdgI0+FI1MJHgfC
MjdHGsd+wm4b0xuvZRuVu3oEWKSKL8VsqNev7sO9Ccbv3qbW81Qgpt0ZNLX3JiGlm4duyO6t/ESK
+Q8ZyFyC2IQ/2Vi7bFyLmKN9kV4x4Ar1UfLZgftVO1s9lBV8scnBnE6VM79sVmoiwIQxIDC+gp1M
hGkeJqrRnwlcnvZthxfNu3BjCADsxkYDoIXXBadbrXv8PmLhf4dXXDJFQll4CdLifWKB+N89LrlS
8JfmLmb3r/va/fYa28V/L8x/k63M/p3ivnZtb0NIptaUzj3gxz9D69kz2TeEgng9eFW0MapNPiv2
/WoqpzXj6aCI5n3870KvpcAdrRbMJL4ljXDDFEa4AS7uHEfdRWXFOxewsGaPjZwPj8Ba/od1Hkn1
b0YPOUAYJErw2jknwnZ/LpWFHsu12tlzVx7LYlVwxvNrifhU9DTs8pVA31YTLTc1eCqKfOErnFjv
yeMcmEI1fMjWSWY/CLq5C3O3xOIxGwPds8rgekYFfgCT3edJzgWscbCkn1o7F7OghGEaDtpl17Fp
pOrLy1F01EVHNqepp8P8xR6WSdjm7bem8BEW7t5SfFbRFeCF4ZvGtFCCx8OmfzbP0tnk+K4KzCp2
KIFL7TAWTUv5JHS8T6w2UtM/Fe+76TbVaa6qtW/EgXl02sII/FjtC3fGswbXHE0JjBw787tQCEAs
6jchP/lRWTJu4xZ+BOJJDN6AZQ8YUeTjvWVHlLw/Q2tpTZ7+G5CexnW6YI1xy4fiRchU9Vfe8Bzo
O7LIIjlx06Xo8h3402Fej2e5GMZAFYsr/UfwUlrb4OfFMETA0MfJZREExlRcYGP/ciBqUf2oCokJ
esuydHIg0hIgm71TS/s/dkVR97gsz1i3RH6DiQQZsEpoeC/81sSmX2d31ypTzFljij4NMGOUuM9Z
ppLskmMNLNTomRQzIt7q113ePjjPUFRvaLO+u571IG/KxUeHE6KgXcA6Lj1G+ejYZ1qe7NhjIJD2
kzgMg25aa5kHvdta7N35BwOa4xpWq3vBoTkJcU3PQYaz/Utyl4TAT1me7CQNRrrGZ3EVwrTP//rn
ZgPr7x9zU57BVw+p0CUoT/uYXGWH4uYZoJtK49hPRnnjvXsznLuY+PofHD3dEp+UTalXsh68do9e
fVvEMf+QkUJQ/lCmcXx+exsw3gjYSz75lfXNL1P1r0xw0pC8BxU87uWUVpZ2Se4cMwzR1a62WIbR
cWtfzYIQg25tGvKvTee8XjN1/tTHVH4mAOclfB/cT2BP9bOtKgp2K43Eels9fYPVJ1qVs9Q48AmK
4Iktzrl9puSyTT3oB2wiHkwlVnknsUNrWjLEMMFOCsjM1+r/4DJhk7s9p+Rvqw/gf3R4hRSMq/us
arD1X1tEfFwMMSWMSXYGnRkk9PAsWiuq7Ynv/UXz/Fp79YH/Xxyn676Op6v7PQs8Mlntfb3Lwva5
A1seQbcL5VU4pB6ZOnG/63Za+8BYp+rCbAmUPlV1sUPTiHdCLPERCI/KGgoKS8yWsFfnrp0RqcZ+
a8puKj43htCyhU/dduQqYembcjS4nStL4rUlZZgV8tmndY0RsBHpbEvo5iQdl2qaD1pebezThr2R
tLExSdWeCYadkc7falPh50m8mdIovWd+UxH9fLPVMu6cV2GICjNC1hpCZXzu4E969fcb8INBZxEy
ngfcwV3Ty9hbza0jJbd99y7fynvxShQYLOua+mYv+PRWTY4Lu4YcaNFYz9lpoI3+Z5ag9PIKtESp
ofvUGTsn2qmThYf5bUbc5ReDF0Jox8QJtqPIIHek3/HUjNbRumwi09Q6rjjfIfOYw1Aydm+uV4nz
V3bBhqWNNTu65EvBo/r+ba9NOONutuUomv7an9JWDdBcBY/ACffJcnT2pdmlcFFfXH0+XOOnzXW1
leOrAS1gf7g2fsNGSVtR89k/SlthG9UTvZ6IkvztSNyCXc5DPSc0J/Q4Ba17NdMmSzRznCRa/bXg
QbkLj5v9mM2VoE13AmrhdpJFWJHSY+3ANeyVdBxJiDkJjGMu0Hb4wvj4E3/OHqE031rTnPljusaW
LU7SGbrwjrk8wYhtEb9mD85+O8xWZen+Eoh6htSobK+ooTvbgmHQ9oQQcN5YZQ//gBTOnhzcDGJ/
tRipv3nWzD1qseo/QIqRbbi8SqB6foIVC8ELHGhZ1KCGtDqzBwG9UI6kvp8xEkt91q/WK2ytNv4/
9HUxij4ypSme+BGifh/col4PAmW9tm9ZpFox6uFpWIbgYxEk3LOk9qOhmGYzvAkzAqw8zRMlfS9p
HHYaenjKqz9KHPeFIZVHNe9a3y4iG8nUEqP64EvPHIU0jS8F0durynKF/5IcaE+2Zcbq8Qeqebth
aQWJGcl4AP5j42M/NIjqFTcNXqVhVFeEsncvDquVHx9o3c18B2u+Qvt9pjJ4pqWMOkhHjZ/4hXbH
fX6FfM7vDAM3ycknXk8izgF1/rpqBja/JaTifBQvtf201Yvt9mE4ynWsMBiICQbaN4h0cY0U9/Vm
IlczLn7/MrZOplhBbKG3LOZjeiBsh0W42065N2yi2onGa5wiHikwpmHmgt+10eFGLSQABIHCEogd
yufEY9RudX18nD5+5wCf8I2VWAvA8gjGprXoPelJKuPU+mPFqvFK6WB+O8BjnUNn/NTezP7HBUoq
zumtxNU3SByOoumSLQQNyc6Hx1WEZUdx3vadpB5ih7ODUXMfq7q/njFcBZJxiKI9XBcVCI8+oKHj
Q3KQ9tVbuoqetFXcbsyNRwE6PsOLoAXqAW3mKBnbIfv/gjng9FlRKqHA/XvutooObF9/hYGBgtWX
9UZXE3albQRvFTO5J5PZgBNpnlxpcTtFAPIuSJw7yldIFxUIqWuxh/zi22ha5jptBCKba4q6tw10
z3s01JF9mDC2Dj5MxZ2199HpTjfYY8RFyARK7aeUOZZoAoP/Exhj0Rn0T4HYfUTdbM7bHIiShgdI
q6MWnSz9swSFqm9+fY9lqRmQ0Wt6/O3l2jB1eWpXd1nRLWwX9g4oTlAgo6bvm69XvepoPze7YKoq
lW3twvORxt0SzKR05Tu6hzDzjjd3DagHbStAKZBv5NBB85G3GDaeQrZzAvYiIk8RFWi+ULIIrlnr
KOdqCM4aRvAZ1A/NVLk1lu72NRFpYuaaPecA24BAadC4oMdiTvbxxS9B0wcP2YjlZnSSazODPPYn
1toAxfz2NMUd/Aio94oYf8qSxUpaioQb3MkJS5cKHaT3kDVBCY1FOflUf8rP58ibhc7m98dOIbH3
MKvekV9KHva+IhIaezFeUhGFXvgNq14UND9naScV5O5oGCOJoiaZ3b3rGIbR7IBd7NEBj7hiCaSS
iV1C6YbumZ8Xf7EV+Dea/YMEz787RTjCJp3DF9zDilPPtBijKGvBfm2DRU7uQnyp76jWjNMg41I7
8dE4JdsWji3bxp0IXdfMG7pexmZd6EQJF+k4RF/f9WrYOHSETT2/vC10JLuTUWULynBgD1KPB6y7
QKfNIDhjjR1+c09WxEF5IXdJzQKg+44oLC2JhyBb8RXYn/LG6Cn6udAzJ4Ns/Eo/XUmzzxHo3MOH
NphowY3HUL+gUQHAyLT6vpOq541Du/DQFv5Nwww8oF9Q4QSP5MqDVOtS+QxIoUXxCf/EGAhv7s7l
xisjaTwgDdZVRgjveEfh6xwD9W9JYYHUBFanFQIlhJPwjls8aO0braL5NcIYdKlgM8UbeiBMLRCw
oiCfNlfTH2mZ6U8vr6/BZL+JApb1/a7FSxORnfZrt9bU3FHC1iWVNPrizdExukwEr6Z2p62Em8VO
99Ah3Xti+dKRVTSsq75w2+NQ5wy8XWe+hy/SP8NlNbYNZjeMODnb565h6lOaDdjF8IXasxkO8Upn
sY++CR7LMZ7jGyIK+jiF3HKtr8sj5rXTsFMxxhrnKsLkWVTu2noaux6zAPIEDhtl9ZiJvR+e1vvh
AoB8dMtPgQyl8qkMINjsdo/LQqG5wrFzIFMOoW1IxLpZELnpKqdLk05EUWBjDJtKgAqW02SbN7qv
AWDulnA/jPkcJFLlVOcZBv68cjn4Scs3vYcEvtAiD9t9Pt0mP33wMB6FD15ikGiaPuD8PQSOLcfO
kXzq+8nhGtiMm5ovcasJjbSEbpC6QPoMhEVmpG9NkYPC9Aqr45ZbYLrqHMPfHq5ZuekIeoz2u9OA
uNHrRBSx+vCyQilaE9IwAhmwJU36mp/zWOFk5ROg9CxW7BXqK0AVGjs9G1FRYWa4aJqsee/VGzb0
gaKRD3sNAfXWmqoLkkl28sWS6/7SdtuyIfu//0WUuEQ5lzLe412kNpJsPyLf4yiuG8+6Ydk7I0Hl
6C68J390AY5741FU3ncivnBwLGU+3r1D+luXF5BcVR0vis+tMQS523Bd9XsgwsRc0JaGKJohamzQ
LA25EoNXenLlcdzYolmWjtaZrl53c+hurceDXD0G/3Ao9f3Uuo9Jg6ybJhryG4mfed5Dfi+dK/ET
+aTqiTjhYT4xz6FoeWAqkxZTawls8EFy68982tHzvgnTsmYBev9SSy8uv/q+IxzAMRlGM0i9KNhQ
rIv+WGo5Xk91w7KSX54a5uVoiV0KHwlcrMnI9JjGVnrF1ak8XqjE/92ZRClX9UfJfTX/jKux9nvv
y/L8lrMfOFu4u4az286maWJdCM53jv8R+oiehPfb6vkQLhn5uWRKsBY+AYa5FiByvHjo+++PTbpa
UJGT8rQqmZWParpxdAPTqRKiVkNeG1IY1R/CGH8N5rZ5KOKB1hiKH8giTAgTsP83GZrWjKim71HE
0ErdB1MSxgUzpCWcJ+tP7nXyjRW9+nNKJlaOmOcdF4nDy1z8Onma8N9cfbd2qzlzw/7DiF3T2fG5
7lzuVYuniiNCEOfjylv92yM5zk29dI7p2nQt6o8YMYEwj7ZgjPAQHsfaCK/S9jyN046dCtjwKEB2
IGQpGSl1Fup259B+pa1k8AVEZvmMgHYZRks52d6l6uoBVXtl8dz01YKoP1JPMd2GtA+gzD0WISu+
+wyiWIUNzcPL4PsTia8wNueR05fGFEsnb5+2gPTUr/OiR7HH5EuE5QWqh9BsxKqazXpBXxumpTue
gJsaGuH/ndWxDGryiAj3ZURROSgoOpofcexK4I8ik9gI2/bH+gk4QMePdzEWDzkpjmAJAOSawqNv
tyDh9v50GeLYiMuynvCcfk0O6Llh0Qq2ZbALPPbvslZ3S3QfapWsRQ9rW2lBM/ev0mgK3vMnWoPO
6q0KRAUvd7/XpVrW4t2oYKp8KSLyiJQ6otMBmm36UhqYJoXM2jJ3JxYwnRBznhS75W48175XkCgE
M8Aw8Xn4rlTfpm8FXkDs4u65xoismBGjG1X7fTIT4e58OYQ4WnZtVAFewRic7X09kacyQzosLOp8
36HKz+ZAmEnYRkGr/vaHClScuk7Yal2o5boh/kDoPhJELXQhtM5gEgrFIXda5rU9a4rATnB0QZXb
kH0UI1u3c4317VNwl6ZS8X+ADZc9lyWlPZGZnpkujzOIShAiunXnDYLtPKKGo9SxudRjMAQFq9dr
oObWj/G/zlddH5THzOg88gSSI0pDZHo+PBMelTix4mR0LOX510JLGlJJh5XDSW9MWeGEnCxOp6Tq
ThsqYViwzMXKcAT3gIw3AuVTVIQ/tvuHhYuxraGv7qoKLNhpBFVJ1bMEW7xaguFsYHZVsAjb2Jmw
Ob+6iF4Qh1ZeTgbKJLh4oSUh7civcj9vA0mmmSZsbi556C1YME2GR1EDImGneCRyB8a4qzYd+XLS
EUvmmKw2rNMMyzYq1JHifVRdQIcPffs5c77l/bkm5RAjp5jIvMZK3q/hl5v/Bw2H9gMQpmy1pnho
62voLlf/yP9h8OgvurTKYXrgFTIH3sqRvXpihwoifqAKaIDnR/H5N1XjA1MskZZCSM4emOEnhg5s
/r7SFNra1Zi2jHioXSrvoCCXSOM8UOlzfn6MeyUhbHmC42fk5i9Uo0HtSQG9KdPeVVh2Rga1qL2k
OqzHayCajUGWHVeR9iXMAqP0T4SVmh0e9dsVIBu9/9uPFs4r/KSI+o/CO/d8p/9hO8I3KpzU75Iz
vi6A2khZLB3/LBDE8l6ZRMlrpmjURTedf0JmdL3IN/I4PQbTRhbF4GFkYNcpHhn9CcXmK/oxTQsc
6H6xpwVq4ufd2A8jksPZ43zPTg/9KPaDAdUVYAVm8Zd2tEPSCYn3hHpmJeI/59fX70Y/X8OlfGVw
GBKa6Rj94lBvQtPfwSUjqw3R9uZ5hYmcYLP/moK7bmYYFJ18xncyp1RDQx2SHws1v7ljZlND/WDR
8oNIG14t36fO3MDBPVZA3wWbxSPxGbCZUe6DTwt/v42TqVHxo/w6iOPkLiR80Dp1LASdGl5nvwB4
PKp5B5ui9+JqPEBm0xlAsT9O6PwCorT0Y+goNrDKpyVwZ8hEDnwoBGH06lo8f9lNE6kxNnTOtdep
wx/hZ2J7PiUHqdcJcmdfGGvRUjXkzoCPrLyGhAIKWOyXDx2ik/bduXgvcGexfKCSjn8/CM1PICln
i9c9VH87mS2lPelDDWacKpG6RmMZGR+yWC+Se8U0tR5eqjJVru1EjOj/tg0fapj8B6d3drE4ICyC
ItPr0smvVzEX7Q0BFZMeyLl/y/UJ/PiSDJWtCNIrLz8225tod80pjFsg0Ga7FUnv707QyVDwMOgS
ln6c/DxRy0Rk7rmf/AYiMJAYwN1onVVAA4rgTz72+7KHv8glrMJjt1ceZoIvpU5u5EOTUxKixlO1
b5q/i7TS/0lqZH7ZqwHds4191bvUaX1mbub/KgNavM+cqh1vAgRT4uhs2x5xm/0Xp6oBDxlnzyJ+
qXTS+LxZGF3onvCUCluGixNDfeG81ZnmQVgt5y1FkGIinOJzeUkHPzs1imnTWfX2deAvLPXOxOvx
RxwnsThZXehFW1GyWbuNSQnJKRclCR5PHggcdWGlwy7SAbxEOtiNafGBOARhpjayKayDXpQY2EYx
FRaDHY1tzRUOD/1Vm7VlUbAqvUMO+bpb87LU+r699sLoaMoLcTNwCI23R4cnjc2hCLw09oTGhzsW
M7Yy1QhpLZXyxpLfa+k2G0eV00oFKZsRkrwn7mw5abhzpCwcT4XU7MpJQElE8kIB1BDBQqoevoph
/W2aGMbasUqEXM7El9YKleifJT/+48s+XRvK6hZZ+OJ2Em9JJaih8GJ96oarLa39KMl1r//zgTsb
/AlfpPE8TFJZpNrTIdxON48+uNpjFDfiW/U/t3bxmGlW+YKYcK7K8sloxDSj2eFNoyhNWwXkcdtX
yg3B1tkojLv8Y9dHw+l7ZItBTbkrxek9bdlI0jlMFYdlJ+aghnZzpt55B2Z8B0p061E96prFkCmW
vebp6AOqOW57dpV2ULYmJjn7U7mviMWe43eULJ6olW3Yqn8j6P4jiNYWFtqW1Hi9wAP/uM0QxHmg
rfzAgJMdtBjEAe8rw62kdjqcaFMrFzZ4g30oAp/TWylRjk+TIRpDdlZ1fgEXuqyz2pvLUuqVHNJQ
Qhukw9nkXat1HCJPiAYR02JMv30yQU6f7BTNtRTQG0r+BKr/OeTb93pXpFrqAqghxbcN1sI7nNdT
mQ5qH/bDZFsXgUzdaB3UWuNGe+pvHtvd9G8umHnZskfQwQGt/E4jrpyvogxmLKKAlLbNXhRU++Ml
obwFDFlWIsGNM62WTKLIcMG16/d0QUqdJU7gMUenAekdomHDUw11kLhVP7mRc5c9zYEzYq4a5njd
i9Rhe6SikbC7nNYSI7k1JEOOUf19RzT0fqyiWATRvoI8Ra6dm9WzHZTyQ2/UsXSy1puEBnla8USI
bP5Y8YNdtBinVhCCwCxZjY74YQtrETRqcIch92+CmUkXCcR/CdJo60xnXtiQyhji099zpLHZ9zIZ
g9s+CFIr/vQjONa4GTiL4o2rPaUeAS12tBBNl85BWWu0wuuiH4suN5YmOrVLM3fY5NC49ZIQSyG3
XTSfW6Tpnj7NDYzkkZ2sjkCj/lpGJmigvlYVutNGyuWAsjs6zBHhFqyzTMOd3g6qA0kq6sVtpCTZ
zGhRalYwiaWElg0lPoRwzMZgiJiwDSP+Z6qxjjZT5biBtae1n3GjLEhbvtG0MPJGSaaiqe3MBNUR
A+a2oVknB8Xa/LaIOM3u+iaQDycv8PF/lO7Jh2IUpEOrUFc38tBfsKDRr8FuVA0zv19fJI46fZU3
2NFNC8/xw8AJ3ztCff6BGuy2CwsMI6CXlTuHsJKDgssFjh+ZEwY/9S3fK4f4GnEoGYOS0lEaWwEM
TLkInK1i3dSBUA2s/L7apcyG8cdi5L+4keYLKQaWGvrgAPHRKakvVuhMLv38B4UrIozbv4BP59ep
n8dNlcFOM/M2aoBLy3jypmPGAvf5Ad4ybsnGKhu82iLLj1VF3ahiOx7EFgFe8J8XjrvI2TsQQTX9
keajjNjsvSy3LJYcGvUU5akTLROoTb73b0nFa+D1v5CZFdTaDjmXpEyQlC4H2C/FYstrc2p1Dy2S
zZolQ1k2hahel54ljrB8LZ40VlrcegunxfvOzUuh+hX6AnMj0EL7CJoYUBhmeMRUsdir0fOHxT7c
6jMVploaIWP3RZPt4e8xZr3v+xMbo7/N8R0YPi9xVZYAxeEc9nLTb1Zb3wUatUHtoTtBYCumzHzP
zxSZdES1yNgAynwMQDJa4nm3uPHYcv8yA52SKYl4aTCAT+0gYE+Bz9yTBJDPUylhI9IAchEkQrN8
ag6gJZlTh5TtzHWMDXCDoQRcotl+0zX3asd7NviF0vJFSaAmoo2LSqdAD4PaWSR6sk9gEL7nTo6J
lw+LVriXgLung6oRNVp6I+NXlO3sBfIzohQaAyd+Sk2Znrne0Lc8g+rf0drJj1PJi2D541s2tACt
2r+iG9MmOmv71lkrtu9ez0RnjHmoYFsngDtYedvBOa9ewe6LoGeLT9EHQu4AVtL1oC0fgn8nmCEr
Fb3nJR6RR4dd9HqeNE3yERnglNBdLd4TtgZEeuVZXj7yFyQtAELRoqFjpi3k0od+41CBqZGZLX+G
/4aldwjGhwWhykfJretBnZA2mKcsIcD4K+w7E6FUPJVhYJe74AongglwDx65TJv7OlyRXb903V4P
LcQM7CJC/mYvGf462gC2/TSumiv+QFPAxOHARMoFUzIzToEY1t+Qtnx1e+6zyVGe3BEDvWIcBtT6
jhm7UfPvqa9K7IwX9TzP/kH06PsMvmbvJ0JglcHYL5AISYBOWJMjWsXbAi+QfTJkIIM6AKIZ4rWW
uPVbBy24A9nG4fughkOGuPCuWPEJOUGUNptYVc7vKn5WlTKQNFkxnj6A7PeMN0s2aLl4vyUkKwNO
rr3BNHG/yN8ez0vh0IAtcja0dJe9ZQmSmqEmLtJJzDVGvd7cb+fQTmKYdOuDYxMBUrbPWpy1n8cK
xNf03dmrHJ/zG7S+NGgQ9faq4yOWXHebFm4nYq6zXjZjMEmGPoED6JD7FLnFEnnYjy57Eg8qxQtR
wx0fs4Ad8s7qOfVuy3hPA4J9fwviR+dPqxD5xmWuGz1zDk3xvy3BvEVPHw1BWJyjvyXeY7kueURI
r8mx6Rx52veI5oRZlvSWz8s/aKoIDcFqJ6+nUzowQ0/ALYKfKhWYXOye0YWG5ImzJQgoI16TQDzS
BgrovXKLlwEZl+fliLvyiPEErvCvzApIl+mBaHuxcG3bu/T/5a2xKezIcqhxGJJzRTP7dzjbPqVo
BuaM21hmw0QB0vQeaUT0RKoUBsrtV7/JDcx9avXSg6kzsFNBn3V0kMsjFRkOiAB8Nfws6Ckx2/hY
CpI2BC4jyUfwLG4C+tgmJIs9T1y60eHC78YuYq8Ko6vrkkF3oZSHa1l2osdjQSz0TpCHfQOvQ+A+
GHG1LvAS5Wuavh668lY9vA6Al90oTtgU+Afj5lAm94YtrFsPO+QqPVQ00sxxp7GsE2touSJLIKam
HCYNKJI+aK9DrfuFUM0b1hdAYzwcQQ946rmrl0xce5mAA5cMpP+cfTF2vbCmNbUAAWiWg+WKldg9
lyIJfJvavD/uGKgQSi5uF9LTTGj+k+Ac99C34LI1hk0yvxBMc9eHyYX1FRDPIsYUhx3vOmGVYRZ9
Cx7j53vKOVk6/yyZUzBjteXsmtBwa0vG7ncl5Gc0jMr0ApgJj+ALnOQ/+v+H36jknm6/BjYvwJnt
KveGucDFFDM2VTZ7nP5KndbdFezh6TXNPTMDH4VUJrB5ktjJrc7EYtHSBnkxV7aywpDwFiV0QJ6s
BY7p5fh1GnPWSJRtBRI1HKx/8NpzE7RGRcommIQQG1xqTXfvZmvi8znp10DlK6Xdzy9TSspsGl5S
u3JwYiOoOTNX/yoQZhLzrOOW/PzzA2i6329d/eKuUGGpYtFDAwAQDgLeiaUHtwgcYKL/Uzd8ZUBq
yGWLMVDaTuc/LkrMLTcnlSzrWufEfic0xpIHEfbqUHcKptkTkbU2dkZ3ZgzsleZKFdvWmfHKE/lv
Vak4/NltoCX6s5yFIjbPscLj/S1kAtaC6yJmjVwNca5E1L6Ov9+LdOOOHFQfoE2hCIzJn0BYGaDL
DmT2jSnfYsKXjJR3yrcHQQrxOV7c7JMbfWFC9srfrAPfaXNLVGMemxaSzzEMwsOowSn1J6zXmrYa
08qogH3tlcZgAhJz9nBqUbXbBv51rr3J0wS+Qv48y8RClCJ5MPk1vWYT+h3qzVVICvsuwhby0vH0
/mBVEzzbZ4t9v2p+uw4ML6SLSEsS3W/cQCpOGDCAHmv6wmhCDcrhi/VZrlLlrKK3+OYOyhVnRwT5
aiNVo1MhFmMS54jDl5tLTQWTdZgLB03jQfJXcPYGsrbqY33bG2zFoE+6IwwgR/dR0UFnU/ESKV2U
0Q73GaKwrkX2Q2P8m9fbMvUPAU6KdMdkN+PAImHsl2n3zPA/Ipnvdl0s55Ly4BsnQkWakhURta8O
U+g8hjHeGq6cTKPzxtIlmPwL8bSSEGA15d1aPNWskt4LniRdovEi7EsJpAwFg4aYmlQ4lXZUG3ES
fzrcwTuJeE576oDUHs5MjthQ9PYs8cnnh4YLAgnQxtaIjIf1IKkA+5EelVWsVZuALDfh2MUee6Wz
xBHlfbpHQMQzleH4qf9l9Hbt6g76Ev8vFgmQNKdBVWbmTlqo++d8WMDoFaQ+2HHV7IUTtGcpofFE
9Lu0y/+uYNt6Bm4/WkQbFRGaDHYkvdnLEQLdKPPBDpJzk7gzD7oJYQLRDL0WRi/mSbMdNOyVw0wS
++3HtWJVLqpOkXmm3gyiTvV2SxybggLf4mabmcKKaMhtNerqeQVblGX0y7UM3aPo3Gz6/CWdd0pK
8Mq0E0SQUbawjvD6YD0VvuOcrjz3W5RQV8uA+iGXPx9aiG2RlDhJtGYZNq9SzeQvMAR8Gx0+SVCX
Dgwv6mc0FlhnFqVdMDSY82m3V6L9fv0mA1hW4Fni95FTeJ4561k9JNulkyh0i4YuhxGNGcn9ub84
XWUi3SuSe0C+E9/LDxrBybC8yT81p+O1YDoS7xpMAXMljM+WzFbMaWeQJcRqxivbWsBmiR0VTm9k
zKXkpg/rCM2csijWBReKDgUwUMqAiZdp1aa+tS0cM31xbGLk2+GbXM15g52/+RqjSs6ehE/UYVjA
/gu6IP5N5BZvynLLpWoMHopCn248aF5kbsiAyUNCn0fTJAdTlb83DQr2Tjj6bDZhnAgcpbf4WZ4b
gXxpjLJKBhw9Mzya7f9NpU/hFuHVSprcLRIzH/njg+rT4PvDKxLiv2dp/LBzkb9E49G+hwiwhfEK
AjrlVT+QqjwHZWmNrypbMgfA318bv/NzEjhFdcK74Et58W51sdQD3agAR2iOEHuUchN6DP37GyUw
xVVk0GTervJlwNOt92W5NFsSAJc4abPBEgyxl2blo4H9XX9Eielz+ur/CUojkErIom8yQZ5+bHHc
oYx33exJE9bPeZiPxrrZHlIKrazAJxKSGE7uEb4pHGhJlcgii8vWNlwxUJW1OWPw/Syvs0HsNvPz
gQFEyR5yvK4H7Rm4SAoyP2ydNexMWjLzHJDF1J7UGzmtdBPuxCFpz19iKyHlH0khg8mCQRRjnl+S
tyXizQACdf2fQYJu1nyiARz/xp8HJifllATwR84sWUP/plCpnQeKSmZ4CWNfu7/Dxr4GyLpVkW4+
SzLgb1iTs21++zM1qgTj8p4xfdzVSUizKEPGXGglGyebSKHMi787wJjKTy5XzMO42Gn/49Nzxxcd
uAA1VZtidNgjz1pVWuispWOglKstyHlxbaL+G72aapZbpqTIx0T96FQJX9KImApSGSwyCeOvAOkX
pHa/I2gNg19tuYpWz5oHhAPkNG+96qxsdxXvomCSG4IziyE1K/VfeS9dIeTcjik548AHZmozVqcM
bJQrLi6lpE5vvHP1DMSDDUMHznVcDg0d3RqyHfz1ywsYNKSO4UfO3LzEv9D0TTMmy1XxiymMb5j1
CncOBYeOr9p14TNFrxzTIOanE6sBM4W6/TXdlG6zMcON67L7tTp3N2Qkjn4GKb4wA1fZsU3cQ4aV
w7pfoBq/1OO1+ws8wVLCp/FFYvz+6glpvD9Ig1/tYHE0CHbKdRfqA7W6KNXUvUTh7aR7oruQ3ptm
bKP5kJoNbn9AOcOTz8T8Dg1rKvRG5smVQzVtpRhJsl/RmPVyEBV4tNY+Lxh3iyMsH/jI1VwL/3X5
9+ZwnW29b+DcXa55Qyc3WjBWsFp2AnDULUGTozyhBkpYgQZx79noCFmJrBBdhDP5dmtGhxxtrBe4
b84Nuz29xwinPTG3bUkDi0+8b8XXGdTfV8mEDVRY+yHzmNHpszteXa7ml5IfjQ/5+/5Wojv5bpsU
gl1Ksx8/4ByhLyncq3JbrZdWLM72rtOW3+ox+h32U1I8eMu/9en62Q4tL0WDN61yKJvnvvJTzyiF
zJ9VHNG2UuJ+gIomGYPIeOfvSH0o26FT8ncQhTgZXn9G4W9IwQ/tkmVyS0g4glNsmkWPZoYoUzuP
0QVa3d7p9eY6TjP30UAgKt7Kf/wmw48w56ekxsbDAPXMxpJWKka7W6DVRoKbQyocPw8RuOOL8l/L
nOCuq+ftFWfHfKuLVlUxegKJegAjKh3UZZMpiVVCDSAoIINKJXGUJWHaK0H7sv2u1mF+/p0Vpl9q
da1rb2FawN646gb2WTQPhFYMcxRDqIS7S13A1CpfzHxM3j30uaFUJcUZolqAy255kJRTIqfa10aj
Py5jBKG+P4TIQyEkG0JApHWPg1ofN2KJte5tgs3uaR06swgxr1MiV3rwCBZQO40ERtB/6D251rDU
ctVpzF4JvcZz++hTUT5Z8AVwSBX1j5aqv53NlwvFjSrTd83eI5ls613Kfvd+FjI7XwXgay0cuHTz
pjMTG4cERqbElF8rho02o/nU7fOTJ0gP86suiEFLC7JLgEtEtrHRUiSHB879dKTF4Dpqnrb/tqd0
LFLyETZgZh5z7Rfq/gcvEivV/przOfxXQJVX2TytUkSq740yj2spOdB4pQBzftwoaZqU2OTBwAZQ
7EPn7tWYeNwWugDwcSrspfOU3g08B0idSF+bXwO7y5o80Pw4/c98bP55s46etAwqbiK+W2Ma2yVT
iHLfukxxwNuWmZuuzLF8ZK8bvV5y5x7i5nusumDenZLLZR4ywlooJTRDf/IVZ2sIb8WuygBFay2F
u7qSBFYuw9MvcuWOZZah+DSuMvmzsBUognHnm8S1RT8w1qZWpFCz3ys4I60hJ6vQAErQ5Yx4Cp46
7GzI0p+cncC5GVfUcEGB5aJy3sLr/0Fr7x4X7600KGNugky61pTTNhkfAyGlz5mwr1aIdb2fuCRZ
T/6DJlMwAiagSsCgpPwlZbftfxUocFivZ/2tyePBAqg0SgoGtxlxegNU4s/6aauPo948Q9devmvo
ur8Up+ChFalImWyrUABsQUAiViZ8FF93zjHSuIl6uxTRAGBjeYc9rzpT/GV3H8+BrGhwCok0LKo2
9oEng8LaC4asimc6GQRg0PGtK7EjdjaqFudQdiqIAkBrNHZ0Dv/RelPKZzKLCVjkemPArZBk9EWL
K9HLJkrZPfSYy5y3nM1kAgNR4gK2tkRklfcB6fi05PtA5ex8XiB+Lg0IaUexuDXhQgoHaISJFcN/
hcHmtok5+k09rwZcQkiTSJGis4SAZzqMxIa91NEwehQTDNFTDDk8exRv2E25iKeCFC1oyR7YWUUU
yRL28cqzvIEloKVIqW8KPkmEG2xTs0LCy8yEId1hLUOdVEfJqn6bYaXYjNbgGleOgTkXyw1aNePf
LMdT1dkoVx3hzHt11M6K5YZvaWOVxIf7It2ZyFLtTWwDwUMHph373B7K0mwuxbfMQ/M4FlKWOOtp
+D8UzmBLUwN5J9Y+PetNWF37IUG9/N1vEaPhnKqiPKTzqDMREprlbWuu50bLFx5qKB9DOTuTflNm
4FFORCpT3KlbGe8KfQATOurt98k/jK6Bn43JgNq492nDTwIVNC7Q2JFLiZ4hY6InMergPb2c/fWU
0xg9BjZL7bgvC6t0u3eagb/gnihkG5dxTLP+qMoB448CykuuG9DV8LDDWiZ4GfIfWtFxywD0AdVH
peZXLqolw42knWz7mROzPVVWWegn73gwIdFePSrzcM8fZmusW/SaKDx1ZSREMe6NbgOJMoV5P/Gb
5Vm1nFIpvNPaBnGMyJodW64BAfmRxyJuii79DpezvihPkKjIwwwpZCcZOW1pENFVhUav8wXF14V1
BSJlJ4SEkvU/mr7z9I4TFkdql7B1YFUJ97vqA5Xuu7V+gHvS1BgW8/I9InzskM/vg6mu7bISFRLr
gI4i6Exn8FgiR3ZFb5qSbmEKjnYnb9+RCkAGg+9M0aKXkJ3vBeXEhjstoAQR9rCcAkIaA+LdYHHW
QvUbd1Km+wHxrPZfcWdBOfabjl7aE3olv75ZBXCwibneJUkN6W0TcJHl1glCdyG0ZdWpWpqjpgUP
3HwY8S2liCQH4WOtgHdTPyIVXVPjICs84VuImar0wu8V7cTNXoYlX50BRapYaYl8w/QmmlA5FMxE
jm2hGJDsX1/UyuoYPlEpnXqFoc5VTdu3K88lqRq+ZohlKZd/Gs/n9N9BZ69hDB1tqnvGEdDpyVlV
OeviW96qdL/838MAjpRAwO9n1XNIkm8pXnHWm2m/9CVthKVGqGBawZkkYUVcEoQepkOIoYLgOPzX
5jdCBpaF1RiCqPnT8UweXKcDqYrZCPVnFC2I5rG0TmysckGehn2wKjxd1nraFnKf9ImKYXbG+OO1
FB1d3o0It68BvERruWcKbd4AukN3b03keGkF8aJCv8kJ/n1aRrDjJU3nxuQbghLVW9fdPIV+3Cte
GlvF2ppZIJ2XSvyr7VznlY2o4F1Hg2Ysa9M7NPUWlitDkhQYx5HwuNkun4Ra6jIg+JcnJ61f8cKm
p+D5eT6hpswzX3Uf4Wal/9dpDUVfd/IC0F0GXRD0fRpjPH8rjwoIuguFQOft8QUCPv6CBeQKdwNl
mOIGaXpLLpBUoVolm4tuIYzD/rurQmLwe+5KMMw61OPb8fJ5YP35pqjBBfVclKDeclIlAsiUajld
iqynYe3ErWZMt/GerlG6AKh7hkl+3Hw759gLIRH2jZTALLDy81fLQzK46m6t86HHnC4+YLD4wLxU
VwTMyyv9LOW1gN6WO6taVdGmJE8xmg61DtYA2ssJ8BxHrsGy/YzvnDjnY52jkad44azjfmJrq45s
c8n6gTgUCLt2RO6mLZaeb8ckTrpg3/ZDnBb7oZf0TY8WTxptUNO4Vb0lpx/0wDVJCamvG9NGAlWc
VxL9a8nnqrMO1dkHcVHZeNelTEFmYU1OoVOMKsF3nLG2eD7sf4fyCO5aIQ22FdgdV5xr+dbOCoga
CQmzaaOdEf0NF4VQe1YC+Tz8SPmowb+pLPBHWaatAVZvLIJOlS823lGYXoPIuBSYZn7BYKd2q1Jw
cMUCCdoPg5W1wYam11LETK5Lwd2D9wsOoL5WUglG0F80BLPYjNiD/8v/VE0RrDV/G3kmh8uTELJ2
AbmW3RRZ8rbTC5sgvmiYjpGMOzd57IZStXR6qDoGQEV3Il9GqmhL2Si30ufpy+3wrFNDwy1plNb+
hWBaCVnkD0JhyIe0T0UHYdPFrGL0yGM16YHsdI2EXTfI+DZLW/IAVdvhNHgr5QdC0jUlZj1Kgses
1zJ07VWWzlJcghYmuMl/1db5mm6VjGa5XYEZ+G9TBaQ4fIJVZkl/R2gGNtoctFjeSdbBM3FaaJzE
tRgZHkf8SIvO7akJDum2al8CRAL3wnk4o+2pWZkLtrM/C44W/O417LLNpW7GoyOpEJZ5CX/8VHKo
vgcGwos8MAQ7zJ/YcU2dKesQgE7DWd6sALuvWcsO+RxuSNbJ4YZtUrt41jcuvKYFO65ixZwftk4c
oUgH/t1fitfHn2fGl9uFcgP2hHmU5kVN5/Fciz8VrUn905Lrji6Ij8YWzq7LOe5dRN0ICISu2bA0
PEb069Pkwdkd/p72ifqmaqJHvHYsIRTQcUVzyWja+NYl6ZJel7+cP/sCZYplfjppwpKyDY5RM8Bs
N8A8kGtDKQTuy9MjlHazmN4yL8rHZRgOf2LwN8X9i5B5tgcJnDd7JNLyJhcPbXATXjB5fraOK1wn
TJmRwRSI91ZcduLFmlooJ0WHMJFbnsIsp3V/PWUcO1/CPHwmq8urvUEQFiUFjUXz26N8emv5zdc+
8qiw32QkMunfdhCM+giP0pDr3DuDEeGtrCfumn6SqD+f6gpO4VFGSj6lW6Os5zyCGHv1cdH2ur1O
H8dTF0UGx4eFswkBq3Mx+gK/MSU8l1fz0UaFMJXuEQEaIP7A75BLBYZDTMi5VY1m/8PQZOmvX/Do
VuHssTfAhBiWaM/U6558ZvSbyhQjGXjhz/o27+oB6XkHsQnfETT4kD3TprRi3luKmZkPqZxZP53I
OOOx9OiezWVzxPtkYSEeRcP57iyp2JmTKfL1lxmSIo7mOp4yfAev3o6d7eNL2QK53YcCa2vM7/RO
01j+teeymv2zesOYDAMZoNKDZ8t5waeZqgDbLNErNvkpimJiBVkr74Pb1ZBwrOh3k9RXj8lfa52/
XC2zGre+3FE6MWKG2MVbpIy4TG0U1rBJ+Vbhbs+g1xyCP2w6Swq+AOniHtqsHlEmY5M2tSHvYzZA
gGmqSIihqh938J0l8pvFXUIW6CySqitjZdiRmAjWg2bixR2CXe09OHl50JDvveqtBg/XkNysfIdL
vXk7K+b0gA4/hbADHs4eGbEjBKwOib9jVQXBnUxzz+EC/Ke7Lpycu3NGz6mgOmJfCRmll0Cwjsd4
hDbULERBDxtLIseomSNj5D5noAAO2SmScLw0AwKgaC2Ji6/8ko39IJsb4/Ygrv8pCB/XsvDdldIu
L0CimrJD8pM9XEuBo7fPp6mrw334raNqBI5p6Hv+8VKwTbG5VF6a+wCHAZmoNKmxDIbV8HV+UiW8
y4GdSDho6Cn6h7BlOYKcfuXjVCQGcHZ6g9mw73dKIr7t2QiKlRr8mS5+JH9foPKXZr8SJ3mzgCvY
eenimUDM7H/Ne0OW0/7sAJo8WqCc94ucsdSn/4GWZ7nVdi0DAaTChNcCLxwi7q/LTR2BeHVXVMVN
cgzr4AQkRkybA6/45gvoSusOEaD+0zbcAVx6Vw5R4Jl3ym2ZuYKaYMt5H110Hd0/kTun7aPmZ9yd
r23Ki1Gyh97hvEChom6dsFkzAmqZddeeCqgRV9KTQ8GXztiFbNOy9N2+/QISW1Wh/8mvEa+UVHzx
4nv+tbzQ7YBg6FlbzDEzNqM6RKJhSa9hztnSnpJkBfZ/noDVurnLh4BhAnJspmxtXALSfMoDqjCK
ilDO6WXURiTS8aIiAl3hDQs8H0Q1wBgUkacfnS2DVLIbRUJWoZaiwfQEJAFFuZtlQIIMvHYiwPaY
mQuDAuBvKowkYpNjprd25u4FV63qMTpzGxXfsNGCkd3TIJZkmBLk7/4LFZaaDnI/0qumRfj1meXU
vUJi6V9ijAOnJk7VSJiarqwdohJk4bhdSmCXLKEJpzmM6UnVk531DPWIDlsVtOsXstBPeCWPFI2q
Q7uaDDBIpo1hNk5atjaOLOPc4Pjm19c4Fpdm9+qi93/FO30MU2e+KTyKhOMvGEnFp9Da+1v8hH7b
vSnAHn0gZ6ZElPhh4JbFho2l5VtT5mx7pke16A5kLBBIMctwjXvmIRMr6pLYS7/NMk0g0z8P2xL8
FoDC1XI8N2AVv1F//RxgFYt9ccdXt6vjGv975dZEldgcHtvU4/LK6QbHIzoGDpMsP3dLwdUbqLp/
gHZLtAYmwJXdjAMRBYIfOHTcdnFbXN3UaigBYe8hUVDRxQgdkA17VJrRTkOuTQBlkugxN1vV7Anu
SEOb1K1ufHWT90UeQSe77BwVZi+lAXtwQrUle+1gIVRAM2fJSlF+0dYC3o6a+bE+WJJH9mW6O184
Ubc+jsUroZDdKvpn8EhPf05NW44+e20Rk6E6Ks0Dk5ErUilr/ENql3IW4h/quKaN25uIattBCTv4
kA7KVnD7STumB+uRk0/OK9gpRwheJxEAu6JEGXenXJwKnvHO8EKzdg8LlZQdd14u95X/wZr0FPd4
YEZ3kYPS7YCsTv62u5d5OJdSOCVASMb3L+uYTC2vw+NJm3f98Xg8pccgxX+GJ7WJKEArsr/EYeWV
LnoUlketeDfrGhYUHLZUxRP7UL6rngAUFMrtXKdkeSNeVnBhZY2qLrgDTPMWsE4Wx1VaSkxHfxnF
SsdB82iuSEoo6A1dgnM3sC8DspHuHm5sykOp9r09ZoSIuQchATgvhR3h3EOGaZHZ0GdYuZ5WefTW
LsloYF7h0I5fpYQZ+vhQDJc7czDlurNl4m5ZU2oJrhj+LDZsupf9BDrfw8asm63rVFPf7FUimgKL
ddTfoDFnvkVF4Tm2KTnZ05687og/kYowhQqQ7o0iriCgY2zmsYy3OqPttB1rhqI6+qB5Y9ci0+Vg
NCDcTl7pmcgOuLzpfCHT9cRAxXokGAKIoVLnVFeevwGOxKRQa95Kv9MMhtmIIgSzdMkNXzsWl/J+
2bffASsPVS1ziKLB5S+xMQDM1/DisqCWOXIT2ivS+fHPQhgTlXc6NnPawHfAzSumkLeLZfuoMmK1
uPl+05e3I3MHQeFPz4fxyoCKOR13HQxF7dP5DjPxaMowA+bpRa7wuili3QMqUjKXN+34i8mP7pek
faWwvh8XMh5oKT8op1kBD18en/SOclzxJ32dLlh+qzWiAWGfR+Jp5uJGAiXw8xdt82+/z9ty0KvY
H775kjIGv78IcqNdDQtLDA8Hl1fpmfQbEr/F3JkTdcivSn9n0HWt9F2p1TCu8ktOYdyTbMucczi/
EBUMxNKpRmH/hzvcBoXZDKcQqLyRJHJcc0U/8wVoBC22Cj7Z97q7N+a9gwoKor6U88OF9qHJqJ18
i6PH4d3QNbq/yoFF7fa34htYne8qVf/39NoT4mYX3uWQ/0STVQHyBOzhZ5GGe0GodtS0+lXslQzg
PaeNBMniOLJ+DuYriZIaiF0unVVbN6r3NUVFpu288usCD9qCYHMb20hfZ757iogYIMSX6LmzOar3
12P3byoH1P1HJLsbFKRv78z5f+x8UagOWTtQ94tL6X7vPQZzx2L5+IRR7d195ujTNRnjWpR1aGET
AFJ66oGSmPItfBFRwOJF3XnCSC5SY17vOUlu0Lpfq0Qlg1NuAwlFV0iU2a4/74//lM/vkFWCSBGQ
rd3q17B9UZOEUzIcabD9d7SR/XIjNg/UjhiUgtmCQDfQanRcwqd64aq6eQk2ciFn/NdrQ92KlI6k
/0juWJCXPwn2Rr36J7uQKLlw3lDeZLFfAhwl0mhW1+Tf/O+tfSEhrgGUgDt7623Xv6GnBBS4m2ab
7KjbdDYAUhyoFrU5Qm2sfv6+FBbDgc9PNEvIwOtSxyWhIJxaTNW2PTXxO49oW9XjTYK8zMUSaqoO
nYDn6zXz3IUD3EGyT0iajbpPeJwFO4/wyWg4EafKoSuo4gK+VxUgflAA77d1G7ZxqF/V3st4hiTO
Z2TyyI2afd7nurlsTAegoAItNZUQWsIR8f9uVA1iyd2daJaybCi7mascicZlHVsF7l0bMgd9jClt
3bT2OY2MiJKzOAPActO++RLPCAu3hCNb3Fj+us8l517LGWd5JOGXDf8rhdoVwovJwYg5WYjmXjut
P6pTnDwgYyssKvqmcIrUGnPpU8C4yUyG1/PJdM77Et1+UvGTW0L16TUwb/Dk+jBl5mWsLxZJJxUV
wR6jfdOv+QoE2J3nCzGJWRMXJES28JfdxIxuZK385nUjCkby5O3Sek6TcMZnMbVNSSd+jwvSn4t/
ywjlXy4j05dmaFIymUpaO53bCFO8eI32Y6OrvlaBEEBgCZ+9Aaa7TPos3A7pWfvhPALKGxtDjsea
4JHdabtPatyrkFQvJBodvERGSddLjl08woe6/X5QbLJ1v/qkysyLdV4bkx8HVYZe0ALdyrjfcRBA
B1d+x47puax3wsGLq61v2lWdRlvx+BE3V9W5sloEQoZjfpBlQ/0l2HJH+bEgfLduuNkDr1Vyh0nJ
C059rvyYWebO18M0/R6CEuyxao1zNfvycOU82TJQujdP8XCn8iz41mT+ls2FWGwaCoYQqN/xLrqf
qy8Oyq1KBADmN+j4cRQp9ldZyDqqW9FJU3RuHphKTEItbS5oAubksaOd40L+wzIHX9GvQp40RZuW
24lJwczcjW54qWeNAG0DU13Fq7+MrpEr1BHQsqCDIuWzx127wYj+FLcehUlRuXGIvxYnc1hpQ7pN
Sw4DlMlHDhaBMw09d4GQEtc3dGApiYVkH3c100vAs4sPziuVAP7JoEHYI8zIwEgq03Ul+mQeR1Wi
sZpdtkxMafecgqo/8Ff7gBbq/dTF4OB8SWslXwnzf9YznvMKU8KH5Owzfp6/umwspeWIGJt8aA14
+3HdIemixaD0scyrdNHSi6S8xPyKkDZEUVgzhBYFKax0Hjvs3gaQNkHD0yGQcXmAlGICPVsVnXzF
Hym4I62SV/3bKrP/N0wU1PNXE013U09/1x/xGrgrmEZJEzVsfmSvpId8j8DwTEVaNbjafY7sWQj3
8G0j/vee9JEy3mqLsNER1jvjk1Kae2ypFDRYMyKzgyKZBDWpNiCQrjArDlrGiFv54CmyG/jNJbp2
P9R3xBSFAs/FN7+UaBQ/OeYIDbcEh656E37gXHf0Ma72wC/HZgY6FtQCYdOZBIAWsC4gQs4iM1Yn
Oldg4mxtXz01BsRmqETHrIrLe+MteMQE302FckZa9qzJv2jxoKqKiGS4A8a3MeEUcXsrLD1vZngW
InG5FTILcsAQJNfElrSoWPkNTi1EivEsMoNc/gBU36zXkTe8o0GpJXn/25fjDvW2UHbo/W647FZ+
kF1EdsDn1ljgey980Uov4TLSdlrxRViG4p8zPGnP7fOdcyVWwcqgvPvpk6JnHh9cT0CcmkM/MrSO
LPKQaPJaRTuMavFhxSVIZrgO45c+Av6N1anXJDgtzc3DTVrH+qiaXGA3Nanx69vPX7O2AUS7yxeX
kvzXU0eDIu4wXeFRQwUZFJus4EdyeX5K1+7/cSmY5sqJb66dxUJgUD3lwMuGXd+QxHM5rHRXb+QG
cyWMXUOvP+ewX8mEh4wDfiVAhlUp9lI7IZ8X+8HEk7auXZsWXsnfzE4wwdINvTWnYl7+I+q8d/LS
EIzd7lsRoaOx5CFHc5t4YK3RBxLX3aOwxBwNTytjOC+P2DrKkWfZ+/d1h7wxSToftiEG8nMVRmiI
T+twOOxJLAVzdHjOszl2m2ETSrrsBrPJUZ99R1MxYqbDt7FB/f9Bs4DYz9fOh4f3JBgaSsBY4N6M
qg/TG42Qr2jZ/9nN6BClwpwz5eycUXZJxrHQ4btc70FbIk7pQ9zWsVn0UxAZ0K4VJ8IhWCk7w6mc
a705EPTWZhOs7EkHY29xCsZ8moGh9KIs3EnWq6kTSiW/SD+WERGCU0XhK1QxanaQTF7UypFPnirS
1R9sUbe0dyzu8miQsqDuExxEVkkkvzS4ItP/AQYLh3OkQRh25Nnwzy7m6T3sJgMe2Fbc8MnPFuh5
7vEWsLhmuXU+2R+bAExs1K3w3iu/Ob+5K2074U5uQzzLLny0WEXHj7l8p5yZWy7XnlxlYorHr8SG
I0PvYU3gtIa8+gS14/ol81Bldaz+Zjcdqr2CvmWtEV80WrE/Lj7ak1ikVK5SZ95rKiUeLgDcriKQ
fpXu9F+a+C+1R6oTyiHitoy3vjWK81P5kXsIyq7L/UkQlPjW5VsyQRxholJJXE/y+S86xOyFMZBv
fQi8q2E5W6cbRQpTyBNofxpRIL3wc+sNoEastVeCnvYB08Ox2dj0AdJkXF3qj/sbAoY8/rg0zT6S
IjwfpkqO7+kFNqCCzYQKt8pqAFYyBznXQvoolz66w8OmVbySzNGfuWk76Yi1U9ZYRkSb8FXpMSQa
Y2j4dPzBRdJ/OAr4smZ3DHbbURxYx65H6GM19DfOw5/2NvrG2lFF7439UuTyEIxoSiw7Xzv8z5UG
qzwFjnYEZTQbFZHfqt7drxrKVcBpKvNhggFi6ih2LwjD4xIsDWVgeB8laFxaSdUbZDecPCosMDKu
hoqj/257vPJLrUTJzJvlWL54/BprJoKHS45zQa70fWxXP8J+iSwVuW3olzLGgawOlmimCrhQZ4Ot
rag6XxcVXF284bNzetz+Ie0HtFtAKPv/du6zySQ2gyTUgqSuhUrdkR9LRWzJuMUY/PnSBtc/ocP2
W5LrQOdhlXr9r41sc/ajIySa7m8nzqIdOVlJfpgH8KnhROTU/uWAEPynPUz7Tt/cOv4hY9UYPTKS
/+C8R6uNW3pxImbW0IOxdLVmRchs/3kNZYENvVGf1VLEHxGkrIn31vjTfti2PyaO8Ah1aWw6rGD5
LiZtFRyGnVThMubEKqrfM/sX74mXTpAJS+j1bT8+wrp/nNeCcGaUoMtElEsTyR/jgcUjWgnhG+ST
nRkHIcufwrvx0SWC5QTk8e3L/+y8vrFv0lhZCiSe6DFfiigaw9P5GeNPUTsOCc1U24YkxAJd+IQs
c3fFd0hqG0wD2dDFLJQUKWWlXW45du2LZFcIYcHawbDMIokTJ3wCgc7Pe8sIuhSgCljLOyJ62Exc
Ps4TDTdhZnAfH5ZrldLsjb4nuO1hMn2ilpiYnYi+a00aDQ0BvmVOA9jidxWagYXk8MB2zR3Rcrm9
luA1ZhQDh+cuB5LUxZwSoma0+1e57L8gnIXWWbpFUY+bxwSrBGus3iOBJsKDKBNkiUBwMTvu+VcM
AZYpne942DKIz/saMn4noS7YD6ULNA9FSHhNSWsJW+jXuSLhCZ86nZ4MIG747FL0A4ouKARiXelV
p0pa8j5jJxiK/M1BA5fdF4XyjxTmq6yl8ei+cTI/ockNnOXsEm6HhZU8pL4ZgOkyprO5kJHlcr3J
bDdh9nSz1WJSlZu0YQv1PB/9DK/NXO6xR2YpnIG7accTpktO6DzZQ2s7wG9kucprmYg1roIID8Y3
7VoV2dnUepB4+I/6+FLJmYDUDjNHGHA1brQQdelLK20ZhUSzszHhRmbCB3oG5AK5+rLKET8WCKwr
MpH+rDJAGCs9PuE1fFACau+uvRgUScZ6JcoJqjz46LV5MkmFCDRrBZIu4DK9va9o7qf20WxUKJQz
VxJDRP6wwz2yUpU8cZyYbJfnELcWCzWn7YSsjgddC/ttPhFT65cC11XzMa5LDxvX63DXIcrqYlFm
QBiYSnHiM51BbIlJfAIQ1C2dZUowAN4m7+f3URl3LFxongv1Nam4MtEsPHzqLO449DJH61bnMA4d
J0fDI+NMrqRNSa8ucDk76CBuPoRT69abYnT6fD5/lOlXY/FdMMVFPD9K05jVKoWZ12GM6SJb0nBk
ZNsKRYyPhx3P7f6ZyQl7squCiu9YjYv8k8k6tg1PSczQvbMPLMKfsegF2jie8yncPwadjDc7VioR
eP7++4wu+pBHP08LedYx4qXxYtfGNV3ysE3Rhj5qLNpEN1lFpuP3xVyHuh3hfSE0ioK/xdTtBbLM
sXfuh1rodxxmxZ1r63bwzmw1KjDh4GyOMqPKgCPMYmZqO9fD7U/9t+ZxyY6KQKICRyasm0x8voIp
8H2yxyF1fV2bHMsTGQOZQLSRX6ycXjLzQD1OirndayALL0yUeRhcxiGv4Zea0e3WBKVqJ0ar3ewd
pmKXzVbvNL7WUWvCXWCc8YkivlihXA8wLryTEWea9RECcSUngapBV7hGp2JsdIoDUByFWPOPb/V1
I6kJP0/7lcC5wmp8iKHWGomAFiDoGLFVfK/1wnwuNAAaESk2QoE+qrizDCAV45ER91QzKhyF9evX
0hZWhlFGZ9b39qs89YotCibqMf+6iY43DN4ToHNCs450mrsqnUrHuie/OkY0ttM3R5lnIOHmbi5+
JdVezJpCrx3P27fAo1xfLK/lKDvePEUvGy9ktQ9T/w3WFTZ11ohg/N3YfRmM9WwZj7D/cuRX30zq
B129Sz/nbbQUHBiT6Non5mhi8GzZYeYmYUZ9w13GHnZHjoPTthHPTh7unahGICUYxnY1sv3riVRU
zz4ENzJ0X20ND5p2DepT1W7OqlblaXlmdTqZbZNVRMPVK5cKMBivIAOoLHR9Oda58WPAaSPrWzNp
CCL1w4W4WurGY2mDK7qtPZ/vBdw2CSj0ATiOhXXxAFqYxari8yQF0c87Re0gHXmacIntEm0sz7zz
aWutOthu10qJhOcqq3IlqQU+a0lDivmJOrGIMDm9UWpICjjnvvHyw9s36Vzt6yU07ddltqfErXlU
yaxOiZ2XaD35MlgJPVOPqjyI6AZRTz455Ax7T9dWqk9iiyaZRsGM/NVGyWuy1ovqOzeu8DmFwtuF
RwxhEhdMHcrHrQL8fUs6xCcrsuDiWzugqK4+vlw8wPszf6OWWdvg/A/WsRpLGfMpR2/9WZFhrYvg
+tF5keMuhcGUXV1BeYJnVdShT1+fCFAy0aVRBkqXs0Arf3srZxnAAqnjZFVTEwkgCNSo8DeP/Mom
Zer5K4L/WZltvzWvhc+r5Kza9UYRfmH4qS7nHf+eZG2/PoTPjtRZ7b1zmz/ejT/GcBcj3zzlGgsr
7/PwnASsm9wV022CR/aXCz82Cto7KeTNNbPAeyxbbKSEZbfUzQ1EjTBTKOO3YLgriJAWxwItk3wW
GviSkhgLI9xjusz7j3RTbuj2Y+Ft1VY2Z9Ax2JLRkNIFwMVRs1aaLOeVvOmmPFEE1uUlVIHWGa/G
QWL9MT6jNa849Qe3KeLu4NPvifBH4W7NaYRzF6+BUTPis9L/Vh/vW+Lu2ICgLH+X51HxkbKA0jt6
JIFDFJocI5wNsFTyUR1a77wIoTSIEivEDMovDwl40LlP3gyWoPSETDtWM8TVlTxepFPUptze4D88
1UBYb06MQY7nR853dofU9NZUNsgnJ7Wy0BSScNA2TkXDQEzpoq25quofG7DOEyelcGOZ+QSV8QtG
7jcxItNtmV1LRvgrdc12Ug0QOvTo1ifNekhLkfyfmRj8vFx8EaE+DnMk/SpgISitBDqH3+iHqEw2
lReabqFZlQLqHVMNYC1ESHLt1uaOhNGzACAd2PVPXX06Tgcf3xdUiK9aXPBhwSIUBFALHRhgVj05
SxJ+ioZfKqyMceXVJbAB/UezVN5qq/1fMPs1SmcbFrQ1gg2k/yDjwQXkjd/MzBlzHfauy8rxr5ji
1DxUFLveeVRQqI2DWo4jDWL5XZSvXiMjiu/SKRLarnrH8MmEGfx6eV6OJuuQWTArQWhAopsddgXX
BrBOdeyPkXZSD5HGXPhphOFlF8+OR65a7oGKTwGmVcDuEFw8Mgh4Oe6D8ldqqBT3vCLWNwr7pYaa
YRv24xtbhkUsYuyA3SV0VSHKyPLdWYVBSIa1w531qoh8Nohvhe6ShVhLRSoqB2seY1AWzMBtl+1h
Wn7qP6du31HcETvy9t59grmAB1VepQBFyE+CxeZvsObhZmBxan5XAvdkzOfltT5yt+zfy3y7D35F
LmMTOnXgCIUZS2pBru50tJCFRobZnqEvjHXKqmkRLjj2TIUfU69txhvgcrA5E8BAJXYWDZeRq66C
Rl4X5O9rpdldKq5eDAtYyOzYgsTOmpJUXw4I4Y0cqfj4cpiQDa1M3J29PRS6a1G7jQ==
`protect end_protected
