`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
H4jlUGYNLDZxooRMBbWt7iq7jqPasIOOHSg2G5nKxFK5dFgYd/2IIkmGt67JqC3eZuAMuaRlnM/L
eOm7KjUFZg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Q9oK2CFn9OMnEQ6154G5zvUIQA4eFuSooV+UuFre3yW7170bMRKFeJobtYbHzDGvzDOfTl80dfrU
tqoKj2rzXHOHsv+wzu0t1FtL9nPqKXjhYzCEwittyV36S5kfczI9OR94g7cGqSBphlSIbBhYBrKJ
Ry59wLe6rNGJJuIqGQQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AYkjFKJ8U9Cqld2JHskZ9Ai/vfoQ2+IwJ96CZC0Vuh8SGilaaT/LaDcWaYxqHdUdjzCbEtpa0qyH
BVrIbTTxT4hdndaB+G7bL+yYvEUl9+UvwL9VzrcZ3aEmuf/E7yOiMa91nyTJa2xXGqxQEXSsByOD
D7ZjD0fvd5aP+zHid0hSHQ1lOTyTmeWZRtbXw9U5Sp7cAtYoY+dQ1HZg7mEHt66q3638w8bjQZsY
Jz+y+06lWFr83e97x+QVxXXYmmIqn0TywlFsmn6/kEh7Y9KVTa02bOBZJ9iEyktR6KedbGkixDM/
JtJukpVv7PFEr4uX999HondwY1eGwiANX/4k5w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lsI0mGR4YfmcEYhnEBrcadesVRtCG4LHmwqHiv5pNtkj7yPh9Qv8zV0au+5ZERPhebEa0Oyq/vhd
xG7FZ/uD1zFUT26XUo9FMBL/9lDCzEg4O1l67xEGv0w5k7cN95I55ap7s/TsMO4SIHDCYdSma70S
fPPpfjtHBNvMl0+zCHM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BbYLP5gyrqBAnRSoVD8CFPflfHbGpLp47ljuEC+Qq9cJUSRis1J5NpyMQ9mKH60zMB89D4FkEx/W
EsqjQZPOft17HzVFo0k7OwJxrlL/9OCx+IEkxz9DZaMlWM5Lnp2QA/y7mfAmQ3GzXGNTwtzPaBRr
8JeLrh/D1c7qGq5/3HMEAPsziu+SkUObYgwKCzNmhxg1absFY4ADgH0pY+iEBvWW5wjSPhT4LhcX
J51oIZi3EIANzErqayFaZGHY2HR5YlM3ASW0Pvr+Rn5hiQLYKk/+zX1bO6ptL0obGv18UBWtBx3Y
4bh2KhDiC3jTOFfTqu2eknboT8b562N06nZR9g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9952)
`protect data_block
51vt9MLzJ+2qki3xOmBxL7JecnZAHBZS8IZM+YIjM0zmOioo/2ofwFNpPJJDrqKjabCqjW3MH3hU
oziQpmJwGEXxezafHElCAIOrP2YF+S1t2f95QDk8ftm1BzCL5H4nVNtk1VfnhbJf6v0Z3abSFbQL
wsmG1bQB4DQC/DbY6tC8gJjbN/2EE+ksBv1tuZeMgrMJrmNxJHDjkiefrGpk+7zlhV+SeCMi6ysS
9T3X+5xLcVHnqDSSYnY5mizkJp3XtRMRVBDOPiA89+Ho1QnsmVKugYK6VbrSzTZycbde4CNGdOdE
E/q7N4D7O5QZizGISIuGFNFBbLfFooapBzOhr/QQAiJIlYOWZw3Y4j0AJowtEUxae8G4aVMb4RW+
3ql+cFH4uxD06XQnL24dHZ1tyt2KwIXcNdV8oWprqijLBL9D9gVPtfECE+JMnJAo8XVLieRABDfy
5K3BzAJSYzWblCwT5RbckK+sG978cMCeSDjqWDvtg965a1bLG1ewV04xWiuIDs7c/HVxOdbg/pb9
ofz5UjPNVKflFgm2q3YySABZygX1NBFjJ0eQC6ppFiQCpsuzLqiqw9X+w+ULHvEsryif0xlf7213
kWk5346eCVyd3SayiwQ10Vmz0Rpf8wYorx+NCSRojerp1aLzqu3embO+9BZSYnF80xL9hZNqXv0v
sgoHxJzr9yBCzWzR5dFtPQik74QSvOLkeyq26wV7/cj0ezGGwqzSrnS4t8hg1wVa9/P4uFNnu2zT
WLaqZ7Wo3XqqnIeIGRbkO3txwt3nubJlCo9eweIKjDGDYmgKTCmG5mD8TPrUTm2OL/mfabRQqwzp
EvG25GvWEbZ1lbWHcmyTYx4CASYRUnmvQD6UKQvAKEutbyrXEW4HqTXREHD1EMPJqLXf/fBlQyNg
PstZBaJVqixjQ/nkBj/r3ZlgV8NniHWTJa5BnyVYtm4pVWZTsd0sSBeiSrnhhOyMzyvdekTzl3iU
CNzLhlzmg/Ujqv/LIIAW4xK59E0NFEDQ73H+eYavYNaVVmTbtpQ/2R4hPhUgaehHKVSpadJHbgm0
bGyhBktUmgPM5m8VTScOumLYF6Okdrmfhbr2IuURdTMS7nxaK6lUrspsCbA3WUl3CFRmftrEI9a9
vtLPr/FUL5ayAgKw0TJOf2okuBzeAduO0jl7wSZf3cas2gC+nKkYkrOP0/6cKTHFUMbMUXk9yshL
C1s5Ch9lGYUg51HzyNSdxoMi1jHDUeWUGv/sUKgbAFaNfm/EvLGiTCaF/KlBz1bRBCvfygZ4PpZc
29qm3QsThhqIS57h9M5Q30Nwih3exZAI3v3ZFhTgdkm+P/2cD4ac4CHLVNcDxupzUIcrRrr76xpU
vYqHJTLgNULqT49Ng67lTjKt/622NrOtpGdX4/6pQXyD27XkSGSUds8jyswXL1LBUgq2sdOCL4I8
0eCf5vy6CxTP4i8qm/E+Ocau3dTOpTAHRLzxQgFmjy2ifQnUsm0ebNPZfvcFQxQZuuVv9gPbQMhM
qRiEARYh3kqYwAiQp5A3bwGKAAq0ICyoOGEZAXbWBrcTC26cvOGONfIuFq7qoBijXcy5CFlEtjI9
ue7iNri4/8YEFT1stL1aQdWjVTJJqXcAWEvf2hq4nMrEYHsGpXzS6sR84BMrkzmMhnqgTHYZY2ja
yX6+bJgARAqVm9Wz9IsIItM0YZPU118fkvOfyLE/Onlzas3uVGyqqB+DGNQga2WkdpqSFrvilh3n
+gScEY5dLk1x3kn9jigqnpXdpzBvAL0KzAvb4dftlL3+eG2z5tBpMm9HycNP18fDEJkl2BMyex4X
DKj/RvqsrSYwVw5obXdY9KksJw9gYvrsJfLLjaAcTL70WxR84KLYhU2Z4c1M1WiZLYExv2I2CSet
/E62qEDkYSXsrygahitjjW/Z/mdYa2LnlXXq3RILMhoYhw4cebRGMOohrNJXlgb0nZ8gPbBTManB
NKdyuo5OgZr2ksqMgoRRbAlk/FJAERTamz0v21A3SyiYNXRnwNSi5Wdjg5j9T8TK5FmFHR2aI4UN
zB6hL1e1S0mYWqsNfeEBGY/plKtdkbzN+lPq9m/w6PaiqlGBE3PktBovSXxv//a85KRCZ08FVg0E
hmXOD81G5Vii6dWe2tp5Z756cc16rasuEDV4SRT+UrS65qT9NxemZ/z6dOOj9rea+K02njoOU0VH
5oryP7Gt0BJF3L2VOBZzkERJZz8d1v00i/ElA2yvs9nT/67fQKL2Ozi5rJb/JaYx0vi/OUCf12Uo
vdMKbmTSKbERQu/FxVqwmMtetDVgzkvJx9TnzrntfxAsc3MAThb29OSsL+vVgwOeVNQ5+A+H97We
6eplhP7ZzQS1HbN9r7Rb+UkmN1P7bUtSwAz1tF+zlyWWBEdEt4T4wRv1yga2DN8hd0VP6qujcemq
xNq+NjsNsjmtLUOHmO6axx4FMWBl0y3OlTGei9SMDVbAzVcl4JoWBzS7jKAPU99tvCQbtVlSUyOd
RHs85gOxaxpyz0c26LwN0mmK3425ZSrd2Eaz9HvV0l7hJcgo3J3tHSkn/kBcDPqXyi33Ww4kg+Mp
KPKQ9FrdlxzdHD/niptftBgkWHaBCTedinRetuh5rQCZEvt72HBh5DxxSfOh5mwVmuvdkLDvlb+O
Nul3mh2UG6fVSrPTbuAGH3cF4A2p6ttJ+/BDg9VnajeTrpoScTlE2QR5DVZvp0f438WHN+5ybEst
eDsjlSAqH/m1zTQjPb4N2ce1y+QXGCAHHXZb+wu222aXJnCjE9eno2wgjEk7vxUu3dpmJfA7jy9B
FcZ+atQEAuiI8ODTllvlh34Tzjcs/iw1EisiXBFqX5JJ49PiV2dbvfvzSg3kzcSzA7OhCAUo2mgI
pvmbTmCA6F7DB0fU2snek1l4paXhr+6TE5AxR/zP0w2somJBmypXgeZeG2Y6k2kBPT7b+uMMxEEh
7ZiobNG0qKbqzEr1cUWZLbsKimKDMww6C0cZq9KZa1N8zXHEHp84Qxrot2F9hOTSiSrI5CUkCpNC
f0pSRE50b+nGsgGPC/t+Gv0c2emntZ1+tKa/juGUw8pa+0Xd54EtigQ7Jmt5+XTnXlzvbQr3MlfS
QqePZmnyWAvYlbTJe8XIXtBPvv1zRhWqVAkcGnvo0TOMKzYddXifC0tvMV4pB2OZ6rZSra447YVv
nMCA0nOe46YUhNp3tNFL83dzAVZHZJGx63C+FyRuextYg1wC/BJzW084tbA9n4egXTui0HfoMg7h
6+wrZ0eQFyKkbcBHzB7OPiajDdIEDyrivnhgtmnUqb9IYxWdLdM/r/DlHM1/KeVVopfj49z9EpON
Z2xi2IN82Z0MlHQ4yaYLMNQpHkRZb8vRzRz4ei8FttPyFIV9MocHoWxv97VcuPJxfN6pIpgScTN6
NiedFb7Hkk5WKp4iWIRylbnbtYw8bi3QDLQgNaAagJRW+ANszX1mpNe0XPfNZ4mpFpHuQ0lchb/C
WdMu4g0ZVA0xLBtpi6wTsJUr2PuWt1B9rOm1ibvlAjBF8ECpotwVdMDLs3I+aQa3E4kCngOpLhyN
sAZK8lc4RLFbZQqIquQ5jgzbyklaJw50t6oWE62OcKAP2/2TIFAf/zGWBubsR8sK8diSS6+uRJHS
KNpWuI4aru2mw7HJrxpXrYFMY3bQuPwroEju8Poi5Q4vKNbTxmcsqPfaLgko60xfLAk41gmoMSDC
Bu2qEPX/Qshu2yqCmoDOI5sY28Kyfg5A1EvOB5r9dOsKQ+JUo/srB6QPR8u3/eGac2+tOr01LlZr
gEAlhb60hDoGLJv9dQpo8qOe0tyNkUBWX2R7FBZmcbiKw19y0Au9pXJh/qYA4HvudH8ViNNzZsve
/HiCiSsnEJffQIxhbzVfwsABeq/93om8qmvMfZldvluwuXpYx78oKbaS2oRI8xf/aWtUYBv+E+tT
/ZBla6bO8am/Sj4treWufuTXe0T8pnTDkuaUkiDk9gEWowfFc3WeSt1toK3PHhqTnYdxaRG82Rkq
5KPeUDOZOXKLsGVY546rr2GXXxLYqGMOmC7W/jUxUamGVf1tXKmkwvf4jDXHtmB9UfNHNTXvqj0c
Yv4c+VmBEWfoDYfl1M4FAzL8q7LKPlUyYTkSFlV24bPY9GhbfPtaIM0w3TwH+5jbRjNnGs3I7Pdr
p/ttyF8fnI7IGL5HiZ0SvfBnfah/w9gWJVk2mibr9V6T+8MVV0z8TLpncj3RMyVyJ0VV8ce+JSs/
SJAj77+ElMNL1z0d+3sthuuigytdPG7Ruowq4AGVNOgqh093ekXa/RlIZUsG8SUxTninMabeknzU
w0fsKT1kyPOQ28H4TfrSyxFvE2Zz8aWkaaLy40Iwn1TOVd0LXLmvenOd5imo2sIfxt64nVgFzfPT
Rx4ndzRIlI2UB8tTdYRtDlbHJSbMypokj5ojnuxp/buUwawY9VyywVEENu+bz5Gf1ywhjHn9+HfE
9RUKgRJjcRaMsO7DwWZBTaqEfhJYe+oSj2w7WXbIKsN/GnEWmVOkoyMHWGC3KFKXxN7/qjDJWMj2
/ORjIkSXX/IG3vP1+kjpafKtFaJ2tKk9Gk5rjp/JxwD/CZSIBJO6O2Z6p2hKARi+zo3y+bXXgUZA
zuRZr7xhtbJ7PinVpknE18AsDFOkUYuPq2Ak2B2mqv4mrEmEkFM2SIhnmB18gCLQ3c7qkJeV/GCL
TbMidOTH4atBrjndSbDRFmd9JjlE9UUa/WTv/UPet0HTaPq3q1nU+XvTNK/vJUR++Z+XFAbX4jVA
afq/hgemNQiSxalch9vBjQ0n54EkixAwn/djFFnZeDe1J9pWdVXa0xa4GqkMeqUFiLl3gjQ0UwAN
HzxpP5LXkXjAHs6qxvVv+S66uHc1+z7c/9HKyy9KLkRUdK0kJcr/lpbA7qQ8OYCSRbgl+Q2is0yn
v2MId5FGbbImWqG7RBhW/3P3ddWL4fX+E8VrHdwEE9c29AwOyv6xyGjaARrSXqXao/sYjzddzKYA
68o6dFywTobtV3WL7qYAAQjQRIJgUMsrJRfIvm+OPeSX+9ZmTYxsg0v4ORz6mFvMeNNgJQOeeIrm
HxRkXUd11ERftih8FI8KBei5cPsSFMT2Si96CrlOnbXvcK2CV7CVUNgnMuPLFHV5dshhW2RzBT2O
ej01DCCFQqXsIsXB+1dcwKbIoJp78SNoxNVO+NSwdkyHLMkJjMXZwceGymquh3I7j6JRC3upOa9B
rjB6aid17rh530JrcmMUJWsyuSLBRkaXviEz1KgaeLe4ApF1Xkonw0R8VlNX5m5mSxJlk9QcW9cD
loXqRZPaQXqzxWxcHPFSJ6TeZ9vAyMclNHHQflaXC4KT8L7fZj26x+rMunHxwVKTsR5IkWKrWwMm
9vpdJNRJft9cXEckZlBHaJt1wMLZpMMuwXpLfyChNGW3/fS4xSxGmUD0bJ6xLs+FJBh2yvnY7wZY
CAVFADvNdp/5mKZInpFetDyp3/es4Ech7LCWOeNKXbSMcgTMEmWoONJxM3AUmacZDJpjp2BLTcyu
06r8cpcI2wBZjk45VU8FQEaAZlLhhqWXwpEL8Xv2OhLElL42NlTb3IA/LZ06aIZ8u5S5MuQ5LGNQ
Uto/3nw9EByKPZ0ilxsR2CVXmHfjQ+FxxMK937bjJKYY9Rk15aIWHKNymUyI6EcQXyUtp8+xNcRj
boq443yTp0V3zWZhzAoqIg2v/KdQUV4h53bngVSH4APWu8ebfUAuNZh+Ou4VpVEuhoSnrLkUW051
49iT1HPtpB56DDOfu41+q++FALDDzcCoSjzJ6FSB6L5TKHs1u2vIc3fYu03af1dzJ9PiWULwLIL/
x59k5SnGFszDtXx2+vjsLYXpFCrW6txxPcS/cR07KhoBTOGZUDGqKTSdXpOqkNJFS6tcqOOShTiV
TXpTh2jjFo2XN/QvqEzOHwCVSeC6p/w7cmS3LuNIZNUgiiGBZGj4gaJPsvDGngFY8JUxLzHfiRKp
pDt+nTss8WGssCykYtpQfvYzRv5ebVZtApgKk0reQq/+IcvezjwcWjBx6Hjkk7Nogb7q8RfWTxoz
vPgenRfZwxhguCk6SuLnyoqDYhMaHoXx//T8WqbjlOe18cgI7CD61dkYDIpdKSUA1edFHWH/RVF9
l5p0kLgHB43hG3T0Wg0gFjznQ4atNjKWJNd79b88jEgGR+ol5UCiC4FHDkY4rKuVOTRAAuShGNcT
OzRjgOVrkarYE4wnMF1qCBug7+6RIejdA7w6jqChk+75t+6WFkM/1OT4LmlaM9RPYOfwrlZYtYho
e+UiOBcx/QM1/Q8aKNa39ONoFGpAXM/zmWOPSoL6Bhbr86P+KQjhBRS1MRq0OrikKPNMB7RIyKpc
5J+w4djcUB0V+6HEuv16F0wXQGEznxi8+PcvTeDKFE+5LNOo8sfHhj8KfG9LoZ26MB1ieDsijP2b
utg+ysxVLeUkNFAYcHVlboPHOR3iaA6A0FCI5rMqXet8VWVZQuvy0uUWU2/M8Gr19Em3ltM21N7I
cSRkgeQKZMyQZSjgN+A4NNNE0+Fkv5TsOtQ5GuiaIMlLfrAQsb8Um6rB1ag4JMplP5Y8J2DMqqvU
igWTqERGohnOS2jPqtM+llgzvYy8sG460WZAFygJwjO40L4oGQdfteWQ+A8cclcZ49n+V6dsAUuF
kyZwYzFsrpDNfOjB6DUFdRYbMYFfhPVxVu6HPoGuj6dplB/VG0AQAUFmCvSVTqeZeuUgND8n1ZxF
ha1f5Y6EFp/pP0T/WJQLOihSW0/tBte95uIpXnRNH5UA+w5dN66NRdIytQdY/OHq/Y/7xHLU9BhH
OELphs6U4QNYaJ30fLrj/3IwBT2hrHB5xwHpA0YiffUeQJs4HbQWFnAL3uSezjt5zmhXghYqhrBQ
YyWh433Ms2AM5PUc+q/k9RKt1nrusjZfCoV79boEf1kPPdVstksRzVQFNo8QQLr9bp8H9ADzh/If
clzBAGTEfSK8bu3XoYugTjDS9e0Df9w4Gtz8y9cqJlJro6YSzj54/nl6AJkUWT7C+VtwmfhLOaql
7JBZR0teN89YJFgbOY+LW/Q/hG0nmhsQVe6PKu0sNN5uWUTTtVgAfNJux6mGRqHp5seu0MsaRsAx
qRGZZziehWfz2XoXcnRtbAFkXNnf3xL4FZOMboYscp5DvTi9ZD5m6FdZzZXinDyRZC8mukfIsFZk
fcDQABAAGqfCC14SYpxKKK+NeFvScEEWg7VO4ghCzK2DmveiCSFHiLQATAroaO5j7LY6gHYXgUA2
s5wbU0AuVRBuHyKz6xcX9WmToseRA5Pn1FR8kbBP71iBUE11HtXkAKLygxcCD4X45RLcxJVGVYCN
CmSlq9NbUFRqURHh7DCm1a4qu9RjwQhkoRONxAme4OjRksPUBeJelklGASNWlZwT6SVgkKrAkd68
EDpM0dQBpfok0FCOauxXeJUkKVK75inf03y2gitswIZXN/d7mX4YPZHt2nHYiOkw+6hObiyxFytS
vx+xfPPXNXA0R9rHUG+ztTkIit9HXrdOCToah9GlQUkya+1oDanmm5rBPIhnWpZhvjn/NACbx/C3
X7OIoV3w/rkEQNtTkKSulpS6/Uj0xuI+pnMA24SPqlIKyPKFLlegIB9415bOGOuldFpWETMgXNg+
L4IiOIIIUoaE/9pxgTD768MlCBJ0M+bBP7FKOfBYsbY54AfkJkS6s4LVF6XSWk4bUqN2nddwgX9V
CCMxjmlTNvfc2d1diRubPeWCxk6CwJqBiPJl7MVL8APitnxusjUQOgsW2A8kSmYUFKuD8342tuuO
DMXjx8i1R+9oHLpHRe6cRolLBngf5ee/L96GXmvwheGgGHkuoWBqMoA3/ssT7/dR2oQwNcIi1vpc
hN3akYm5Xn1ry1dKh8SCa/tI0BYeI5WPfRGiF83lhUGVHzgaqqYJeff2xrqhHnmsSDwzFgsV8l4Y
jzdHvQ6f7dlrHXn47lR4tRYy66hGjA0J/9yWLhtVx2wQ3NIKPYZ7u8e4nZQfEeljA7NeZv4Qb4wB
ZM5cYa0d1mrr4kBAW54/FRo0I32joJtw0fV4QTZUeRwZsWsbOXLp6UcJWWWB1jlRXxT2l2qFcq1e
OD4CvnjTmCaLAKg7uyH8yaALfX98agq7fTdwEpfRMpFLCEVsXKVPm0/xybYcy7RXai0XgdvgijqM
g5RuovxScWLXuKXJJRFG/7/hqeJ2EdfSMRLlfhBcakcnv9pj/8o3yBUYMQyCTloZMa9bRiVNdLc4
wmZFt/ijiWAFjYR1OHTPeXJUVJ+tWgBSp10EWLr/4Gi+hslrfAnveAzC4J0fGm9U+9T4tJY9HYDf
jG97DU1QxsxUFcoRAIeD8XpVMyAdD6WHmTDWjID4A8i297NYM+dWKKAkcYSRVKtkqDF/4YYcrMF7
zJxTLRyUjcWKyoUObovtdGnBNYwRRMkI/iZYTdrTKh9dnoZ0SZJB3j7kHMa1usppeK5rQRKW6H5C
J69kijcVh55aU/aZehAEbVII5JcJRtNlXC4w58G9ondcNCOf1ij+yBN8332HHsGwlbEdkRvl0nEW
SRiIpaH7vW3mTGobPZnrhOw+C9Puq43iYWxkXiUc3/Ug/FJlEqK0eSghIEg5lw1kYm0PCCystL8U
AZjLyiOv4f7D7FiUeYX6w+R88e6lRQ9rr1HT4lvZGfdVUb7XKSo5FaNa0KovXXTocJPxLi/g2sFo
AsiskT2c6PnnN7RI3VmgZcsl6EuSXWbaal9bf98C1uKju3xAHYV8zsO5IpkhuRuKChFkwN+shbYA
hhn/CM/WCyIRQO+thTCAv9tKy7UbifqLht8WVzL9u2z3OjJeGLi+VIg5BHgASLGGB7GWvEkN57No
NXVzKqgXPH1fHBjMITg4iaLqWScnjI4b9eby8K7k2RAzwBsTWl04Y+Yql0lqfrGp8Ol6D7/7Vbab
m5rSre7RSd8VwYwaKugvzeUg+mIKAyAI7ATwLm0U6ogab5FujIBfcwufQmOfsKCuJSrZlza5d9q1
ByGPFLt8l+nTrF5WPZmHCWAYH9/Ot9J7O3IUQE1dT96MrkbtDGJYmYlOjjlZqepAzHUzBbQUAq7E
Hc7ZRoHglSNtkcPAxQTjNL4saMutGKcEefSHgyMMR8wlzk9Zza5l4jiObOQZemGGndjkuI9YJ0IX
OL8TH3yFmOFmp6KHSpr8Na+tgkBZM8S4yXZfDhCJW3lgFsj9vfklFDu6Um6+AVhg0sBAGy5G7thM
3ORlp49za9GrhtbPePamqQeJn5VrNtigB2gS9UGR9ettB5hRIZLWafCfgdlK/XlaCMYFTFo0kvXR
SfzLoRVYTq4Yx/zYGjqz1K38+R/OeGTCYMDtSjNGd1Tw3lt3Wp3qLjgJ/zacfcQJ2U3h8im0Khtu
wsJHoDJwCn7rU6/iZvbMPGZUfRwjJ9GjXxoq4gK9OGtmgL5Jt5679b7EnNSgNRaVOKwLDXQLshWF
H1ZJuGqpteG4tUXri39/dFWi69QdKL8+5t7TJsAr5MyG8/7oEagxKugeHz+KsrBW8QndLEbO9B9B
g002vKKo5uxeUJffogrx1A+VdhCKOWHY6M1Gpm8kr5MBsEcTHvtnv56DTK0YDiiSyVQXuvnbRjbP
YCnP/AxFU0htGHqUZTcTDof7Ft1ZcZQK0HmAqdXadnN57gIF6JnVhHo66S+GqADYRZEO1Xt0UxdR
KK6xIxP8ND5IDQb2J+rGWLkaWfDYMKCUAr6oU9szaQ8r22sWyWYO8s7aY3jvPC82EG2RHWPRdqq+
eFmyY9rxUcKA+XZ+4UYODd/WuOiGKE6a/+LU+m5dQVP5uOaeZtAc2O/xRRVPKGmpT2yFiS/WoQ78
k4Og8VfiZ6UaWJtP7WRuSVym2HTGfA8RqKALkIjrNuzBWSRzQiyNjIrgoN6+hIiKMzueO15Ix4g8
fQm88Mrb4gwXDHJhVuplaDt18S4dThql4AU6tgBuSTqPRIL8t7lM5Q7uH/7MzXEOsTXQewi/i++D
XySVVkYtB03H5QXI6iBVJsdtITCN2TG8j4y6ERIipcxy7NQXmxn8rIZl43t8FmHiZwlT0HMS6kXo
/0LsKFfDqWsbZ6jbW3gnwP3lcl1Q7yolMEnliDi9WrzK0HMkTTaYl/isJ2I08KsvcBgAT9S9TcxI
l8383dtJHqpBUNucUMA8pi+IdcpjMM1JhjfqtjPiCNa94fLzSJWyQQFriftwSxnhKVrF5mRZcngm
7x6/SjFHCdt4DIVfMCirmFEs9n98UkaEexHwkOy3XIu0ubTMoyhXJmUJM/bIBGcqaK0b5hPvtezm
hPbPtLVuRnzIiT39RluxIP+Qm+ZMuxyv4HCsLeO7ofAUcYXF5RrYd4IR63Vz2JEekvpFLKcEXeMW
qRw49abCoVx5hjrT/huquvl/H0xKdHPlwGT70LY+CTzT1FTylIKN9zWhPWvUNjKwjKclnbQgnRkR
Ef1xnn/Hv7jpsEVdljHfFmqjEq9pNL/Jc87H4blkoAWPDyMrFqeDoOapekQFvd6XwEhzU3C1+807
olWEkLCXPSpFqRzlPvsdlZQUjGlLLhOJPkozn6uXqORRjK7mEv1+KT5srzou7n7ZUBRNsKiNXTkj
BEH5QTO6MIIx9I/am0CsCs/wF6qVWruGQF4ktkKpVPbUFpqT+mmIYVaK3Z3OBgb1bIf5uI0BtbgF
DRtgvyBFC8pqIq8KxJ2LdtBBRAtF9oGp87sythH9iKjHBV+uzPbSoTTJW7TMESRpjLy2FzlXhr5S
GIu/610YtUeEIjVwNMoudzvJ82IOe6ateOmx1ZP7FSvJHT1sTT3JnI1U3czoZPyUFgIdgjhEb0fU
01bgKbAkaS+0Xl9b885TXLvqeI6e2kOz8x4F/VbtPp4V/TgWAHS7crhtHp7lNq+oibz8YK9X485C
wYJp7c8dCbwvRGvw6tsMif8NrX7PAo4VsPY7mmSh7uf4tcAsZSUiWqZqM0tnfsbh+mNN96e46eCg
yyDC/rfO79N8CrCr7RSs4CTZFKtIvlKMl1yQmEEfhJ0w+n093yg3MuglKdnUGXU1XI4d+3yGdidq
ZWfV6qhEqTqtBjI/fXjAT2HXFMB0xp2eg+XDvSrE3TBWAeQ9KHn20xNzrsFaH+k7Ag5QKwo0k9aa
4kRD3Q2617WZrRmcc+IdEari/50WBS0OQAsfWLbBHSrf1tEProOrU4x9DSTrZE6J80oG2UzlCeqJ
1M2oTmMzuQA3u9PiIL+ct7AqHEFku1U92TswWxAsQtPWzYYw1FKXztczO620LiwkM8aSUXKW62fJ
7aWTT1FMldLrtOgGB9q401uE7FeYC0vcnmEvRlaIxHDSqY2kY01wcT800qecy+cVyEF2x+5CrbIu
erj3x1/yiMWVa8skUDxFe3Aob6g77xsV1dr2bVUSFxoJsJrnMlsOr/sfhlvAnHaZqQVXNFKs8pkk
CwedJZfN5VrVWzYmoh2xjupKUWVrhlBWzmDN0kPljg8lRa8b/TZBzKUiuqTP+EzT+W3ao9LlLq3a
JdcozJOF+h5mjYzyGrHec+42xZ3+SGcT5rsJLdkXANmHNvErnBXH26DU9qdgQXoRzA5fIlU5d+Vp
XC3LMpdUPt9pXhUD0k9VklxEx5EvoaV9AzNKte8ER1xK72c3qFiUGmGb1717A/Mnwd1UGriBgvFo
7KVOrAvzc088shg767iZE5taelD6WLZ10e1gbooy+pPi044B2SECm7SpIrFO4Iuj/Agv8vmSqhgH
JYsNFlYK+lO4tWFeFnQ9IWLXCEP3rzuEUtpNCGsq88fX9bXKBqg/RFLJRpnp1X2RH/GDGygre4hn
vOKVr2tHNCotdY6Mb0q3pHHyTpgz3J9dUvJcDgUkRFKMJyLMRyRFkpUsbGcfQCtWALvaqli7opHL
OcGDlpuNeQvp83gyhiVSsZeEDn51INim8aFzBmoRGZjO/B7IN3G6cVoMr465IB8DF5nxuApLBin0
Pqy+4PwRWUN/40cDGqWLEUuyaE0tL1C247QVzXhi+ApxMdjke+xWR/mfhcDBA+FIUpaBzf21s6Lz
w538/BHZLgU5sWskTwGfKsydnNkBvOioet8A3uLm+sm7+icfLcLL5EQ0E1BcCAzlzsjMZSFYaww5
gg4saTzYEcuR7SdnDwtbuWkNR5LPq6dDAZV/y93So94r77GEbxgpkYcW+sSHLAQP4Okl0Qe5tglY
PHiHJKmVBuedCOIihL+gmhDCbP1Lbek5uUFzcSRdwg3HvBYrSyG2WYr84Vw36Jcl4+TcJlmviTsy
06v/owqTN+Yf+5vV9H9sBvWcdNlaEBz78TfijWT5EyK7T9GwuKElIoJnR2ivA0tCMHjR+i7Zd50Z
ZyZ8MdeQaNhFWMy0VEnMrG+fCLm5Q3IHzJtbYfR+GPaxGtZJ6//uS8eqqQdmC1AFaPvq5D4mQS7Q
UHKi5dChveeZ+ZQjzadcgoi/hypXf0YXVwXJGgjIx83bF8ZykwqQQAuUAW8IbBDfMKsE2kNT7llS
PFSW+NYsmdmeZmzxwEBKIES2SzFuiMnTykzkCCrEt6xR1ngyUWd/pEvKnC8+qa1zSLdb+4rye0Vx
WTZf9vXQU2yuBdC3kLlptTqyDGiOOWCkraB0LW2I0Rz7luTWEquaETalctEN+zYgeNJqyWx+ETR8
/roZjq2vLiqRl8BUeDLoQrfYRbjlGhSfmtgJKf235QzFl99k39A7E2z29hkhByVP8N5XTiCO+X9z
Fg3v+991oMC+mI2DQMesuPBGo00wPCW1G7FhfvD79IkzN4aFFHcJsMVC+JEqBqGCy+hxPPcdKfea
9VKygoqWEYhdbWOYnPnmIE4ydSsUxxqYlNkeItdD23n8Zpwm/QcnPX6ffB18MWHl9KyKepRquP/T
ufgAVtE19t+ky9M5hFZogg3KymWVcBrdvM52OC8WnYx2xVndzCpRh0Vqj/Z7rSoRSAQDDOMVL1MM
TzoYtOK29Ez//mohx9Ud8UcWrt6KK7dh1ycOGEAZDDxDP+0lyXdDGHB7J4ViSBjksJLGlBpNyBUi
C2/k/pPNJx1gkbWmLXSy2M1fWU3huRdvtiwZwNSjPbapvFcUeSo+mphFbR7sdlXRaGigoYeY8wzc
OcANrLA3ay35rpBU+ZN/U8174cTWLeF6JOoJCDatgRB5zSdwdxRB/HYl3sdAgK9JzXt5M6F/ZiEb
IYJF9/Zok650tztFp8oSmnNeoIEohQp3KDu7V6h7vZLO+A==
`protect end_protected
