`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qBkDoL+zq9xDHko1dqTIrtCysxt5T0Lw/5e54UpF5yo58YEjYNrIq0nlen0CuQF2h3ec/uZmZk/x
v1NNPWO97Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
U9faUy0Ig7WxX2mwx3ipr8dxzWvz6/3DmBBJUCg/0V0O87GRXgh6H49H9tw6ksGFstr1ana3Nq7z
TqUDkk1FKBN0CrEb1joThh/MiVaRSIjra9tfuQ316L3nrIRA3D/xAECJ2ZxbpXJjUFEermU44pPQ
H0zKPNjpBHDaY07XSrI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UmL5euE4JtOuIZzU3d1qUMh63beEfLkjQXARF9oT/Khw2uFy/h+bImTk3m7BSVyGDaaBL6DmMVOr
LMI6s6zgYu4PBx43ATkcmwyu0PjcfXUkmAYm2WOQ7gtB8It6GI2Wcd4vYdBLZeSiax1aE2Eswpr/
askoaPdCCTiX+yHaJcaaHr3XR8M/fz8VXx6JkiuDLzqunJk/zv4yneFczoBGUP/umtr+Hiwt2RXh
+MswbubCL9wwB7wtb3c02El2M7QjZfVF5LqsURNtnTK5mFGaPQzuIh4FRG2s8PihGiaKOX0FGK+I
/KOvTP8i53vh5l78DJbcRyhhVQSGmR1zt9IHWw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WjRHmOXOt4o8ai/6NYQu2Ce9yHhmGKw1+/zjOzkEZ0q6L4OS5hnd66COrIFzpDixlu6bPnb9Zls5
NrykfHi+nk3IZHTYyNVA+vRJNl9xLci7ESJrZepS+JZer5SquIupGrPCE7Ln7fq2ksVaSeXhKT4z
2DKdyJfVnbbfNnsM/Ok=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VNKW19tiXS+n1eU4hh4+rSs6MEq2Wk9753XWQAr+bsnd/Citm69FjGtlpOBVO7zvMVQJYsj+XRu1
88u8zxsniE7DKTiOxx+fc/EbdACgngOyHQScyGalEj/z7hmg1CijCCVNe+CKQFXltERmhD3eQHRZ
L2aX5nb5yAenJEIK0tX+AxNeSTEiITSCcEl4E3FCohjSU1cbqAVlB2Ha8LJ1Y1ZfiVpnF9y8H5aO
8iMb/rveBvGS6OWeaqxHMKrC0x5rjbd8r2wbDF5pVlI3olzbWkRUGnzG+5d/mMUUKEubEAiBfyOX
nXooz93WH/DEKqE5yW7+IwB/lmfQQzo0HjAzoQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12560)
`protect data_block
I09cshl154RtbLM/VrCC2IVAqpuJkw3Wi4edwzsrGnPPkdoMC+joSiFzh8nIuwq4+qSZ4SqEjiSC
VGUXCxUyHPSfO1D31QVBHbQebrjG7iVZy9JBXBaqdIrChu9XWTOJDFtY1x1Oel78Bc1ANLAa3gpt
oxP8cYUtl+7AbMH74EnLnEtBEyFpstwlO9/qGbNcASXsFuC9Zv0WdkPRvW5Uo9QiBTI+UEMDKVdP
XI982HAmM7F97wM8MIAjCTRWxBu2jihuP9j3qDcZyPBBPnX6CONxxyFGTzKK81JesxsYD4gJ8AK3
Rp2cqOIhCC8Lo40txXcTanROdXxtiutQTHo64qotyqsXwBKMbZNt+rnuk5fSfgVQt8ilMJbxSqVG
5iygFTmAPrJ5IWLyklqATfWsedAIEL2D49HxZcKYwTBQy7SdFnmAbGkYSOWmknW5K9wqqda82efF
p83LSxGOucLjezhUFMb8MYfOSXCKCi7qKDRLgdGTMgNCHV5ItjamLpwRlkLf3jQBARxLLoJhgpGS
OxwTAzY8FaT+3ozksC+TugEGcXkZp5S8fvko8ndjCT7/PsqNe0JYIyk2WVPCh1tLli/8KiW5DRMP
beTJTSjiVAlq9W05I02ny08swPfhXu+l+XBBszolpnsQKVR+HKg9V7OILe8+0FqVTvQqc2DmsSKy
wRfeTGY/2jsgrMe1IGvC5BdgWSceeeDTyILIUr2T4scO12zsebztfAk4Gk7LBgcm96ID3ieKfplc
Xe8UiubOuBQMSEP9G+huXrWr8pkNmioQgiux25SvWFso2C3eFALUZSifT/UnYXMvtKkKVchc97pL
LLBaP0lanjXlyXzmMpwyiI6CTPHu1j2mfAt0W8ZBB/vbSw1VWz4EYvnwuDtk8yQB2U5XkX/pIpAJ
/Jb8rvMbwT6cucallt1O4ukd+nt4Q2ukfSB+nBdTrETfUCXKvAerD4oKNaFTrikk63ai+2dAGAeX
aL/7SwkNwQrDJP/CC57LWrE9TIUPfQng/Le+wSVlXd51nJ9CsWiEQjuMtxN9yFggI8sJdQn/m/eU
ZY18Bk2FH1j26WJ+D44JycoQH2z4krp77Btntfrr7ksTQXaQHCJ732uPXlhbXsgptRpyAOI8/8ov
f3dkK32ytAQvhn+1mkuiz9SPSzghOHO+Swwes/HfZSaXnwbBvsKEddSPFi+HrlKPFsD9tHlnQK/g
4ESukjDtkWCW5Zel2pLcA6f3QexK/Xbf9ppxVvD+njgTto8wXGCkGawpRsUuT7Av/R4K2JnAE43j
/Fp/AOrpwkw3zEbW3zQ5f3sWLWopP6yhLe67p1Xr4cvQY+aSvN0Cs33/fJ2PeolSER2IVoJ3lcQb
kf6bMy3ZUokSQlrMU7ZZ9mhiPFt3VFpY8pOJck1/zzChDIT3eYoEmspYsfPcwne/Q04qR6afQATP
9i/bwUAg9jfPo4loVRXpDu+AseCvjtm6vQCdggryyy3vLVQRqGom7EqV71U2LXkCjU5zoJHyT5ZA
c/tQJ/h6jcCPzbOqwnfpI9YUWA3bdmJcxMznT4JGerIPHuLvu+NH5kWokVDMP719Y+K36Tgk4Wyh
JrPGOTmHgs7kfNRlAO4Yr9ZUoa0lj0E0vkthKmlcqQUprbnPq9aeUcdMud8GNz2/KsQrRc2hvZ12
es3iTrOxy4FqcDZmElCuUgx2KIpxn2DrbPRtsGtBWMwZKvCM4jVlZONITIUhaKV+ax3Im391mO1p
F/AyAspMMsAmb9m7Bu5AI356NJeXIMOy1GW1fKtLtHJbOfJPtlmjN0LQlc5oSLm0bGMlVfHHicpH
X6cDNSCDyZhRk7JnrJtzLWYsJNXroGVu0uD9aFJPOgqdjpHhVYK0mgipUVlcVRZgZUXuntgr/wGd
hGqVWxBoLjF5XGunqtQeIf3DrU4vsBzddiSdunPU0SoMvjYZTYq4mlXxboMP2SgXLpHiGmFlqhbw
fEBSevSfOKhyIlwazbXterG1mMmS3UtIrfcl2+kOmrgNMb1REtLUnfx0Fn/cnlpKNzUaZuGQKRgF
s6KHcAhc011xx+RqmlBsFw3VpnSOjFKKDzO4PP6r48dMJLOeUFFHPEpPbIrmFSi/JDaKzY+D7gl/
0TDcweMfpHZmU5T2aVSsI4550pH6NDhyC4qU2Z40MCvVc8OMOGPGqWLM84bVx2uHxhzZa60Viung
j8i8FdlLlVtB/TjVXPoU2jlOhAhMslg8ikak/h0aFw5xeMOq+ItONXJJ9jBVSzLDnk2Uv/JcxVfI
7LfFIVlQv7ZfCb86j3y+BSQuAdLQWHDhofNmFiJSoYWPq1is2bfknUJRMj1CLKBGBzbeGzXHcupH
0MFOnsHvZWYy2Mxla4QtZlzWGp8uHB0Eb5FYFkhpUorW+haDSIjG/6t7yT4zOuI3pJQiaIdiwZLq
jCaYIQvKBywXA08ca5Gf/E4+nmjN01Ng/Cxj0vvEItF3jZ4M6QSiVEve/Rx62vySuyQ7fkUjkVXK
LEKpJRoJ+G7stimx1YtUkevj/9smkD5l7EmVNiw0QejBZ0credFakjITG4ilpmyQtL9v1jLS1Pyl
jxQqNcSN0o/ZnjAFIrhf3iMtI+0bxp0qPhdnd1sK1crRdVnroV3h1sUGKe8r3xDbXUbeBYDAht8k
Ci0zfJvpZAA7gW399+o3cF4e45gIhExvZLdTkSwMxrk83vEa6hV6EWY8XBFzkSQsdY18bhXIWWCz
SjHi6mfRovAWboL2+ck6GJLHA2xZPfAmSu8fFg6vG5/GIEMtxb5dDSSyJHK5nlVxKdAFtrXcP8bt
8ZVSIlE7PGZfg2X8CT5VnkONqzXUICIcnpoiA0B9FOy/L6tUQpb08cms2m8M4KCgJRshrVqu8gNb
dfb6ZLWJapoRxn53tkiA0hA8PLwwMu3SarYDl6RiupPR8mc/WKbrY60AMefM+zS8K2ETibLLGfzC
hHILfRTDK6kUUbqEwpr5LyT8cwDHVelFdi4M28YU+2Eo4MogoR9UFRmumFCWNPO5yNxbk9hAA9QK
jzDyBZ1bktZZq/6fms1s9ewJ13drfhC0juz56HWKeMcE5PRqrW7lp01UxeAqzeE3W7fIogjKRUDi
F1eS5tIbJQB296+xJjOHG670INsCICimAq8bCCHnmQQ0hbz09n6r16ArKmy3TaVZGO6MDxLRic5Q
mhoD/+dqMaJvHJVfpa6ozP0sFdaQbB1rkVBovty5vjyEzPBK+ejapAd3bnXNlDFIL7AjWpdz/2EQ
M9+ggPm5ANgXLxSzmsnJRBI0cTDHpH9tUco8ZYrtUPr5l80SkZh5KGFV/ejzJVa9hmQbvOxYcIKF
dko/cWtbTaOK2ZtqHhaNQUbFSspxQQd4anv36wODnCEI5gQR0YVCmJKCh5D+oVN/rw918qVgDf8w
u1zS4qhkrxdKNE6dxlZkHFhEX6suVPgKkEJDIM6Bn/Z3BGK2TniASuSZeynMbR4Z9ylVnJLmruYh
LnhAhHGFBs/TvdxvH9nwvcTrvXqP9v6bk4nsuOKLdToRL1b4NUsX6974eHkQWVGxG48Sudohy0FF
C15IzSQx4yH1SZVwU1W0KZajZSCD4qeGn1Kz0/hNfILXqUs+Lde3mqammoFE68LTINQbgWpXoHji
0mUf+yPYQR3PZvZSO03ZBaqWieltHDL5ODxnIeLlOs+xLZCUeZjsTFko1rD4EN0MySXGBRM+/QwF
lIfJiMCUr6uzpKEMKIcVC4I9PvOFAy3M7s83bCPJ8U6z6e3fbgTemUXLeZldn0D04gv/AN8bOJGf
HWzyYmLQqDj1Z3QoiIeodxi0xwlpO8YdcZQn5B44n9msvVTNjMPrl2sbpqFPK3wLMnr9+jBJoQfh
3xRXc+XPDviUYowA2bqD7s5aLnxJwfA1Ps70CZwFl+ZA2rFIKyyVm99sXna70UDytqglK81GOdiM
Y2lIcFP/wlLFBJqkbExzD4tBs7cwy2f73cWjfDuP8kDLNbRLd7K7a46xTDujmyCQyBTCsnmaqrIu
2i15/SrGw6T/eJ8nZt8t3nreGGEdduRbzHOV6BHx3o0/jSqOP9JM0kH/BhaM97VDfOBea+8a0GeD
sQcuiI3sJHbxbsdEl3p+iQzsjRSbEZ45RyUd2YjXw14wO4xC0skRlCus/l20USQ3h4F1zLEjFpog
OWl61N8dPle8l4jAcT4ivqNXPiTa1ep/+Tfb/mzli6CiuB2Dw7CY9B0OQcxKo6JmcHrsSzkrzXwF
sAjUjIH/7+NaQRN5cgmVYyJGtDstPNyLbRGb8JSQiG+z/t0NT0NMbCbWCj3dcLeGfpD7pUHPVctJ
A1zuBo5q/A7z2BYOrrcT23q8IcWB2vYw0lQviZXjR1F5U4o1K6R8sNkPQfTaZjAaZTW+W19m3VQf
V50lYR+0fuV+dW/3g17uDia4fxVXmq1Ct2cHgVEhq/tgTxxhb2hMg6j4yFFrjNoES7RszLzwtz15
dNH6FFMGB+Zdl0fJti2x2ub+vJ6u3g3YKVi5M5vMpseO1eRxqdRrH7y9hJXukOuP25n0sCcjH5Wh
uXcW8C+MQQyhK1PkYf4C204+IndQg09dA0ylyAust4m34HqO0ZqphhsatJlc9vp2LNfmssYZozLp
lUutkRFJ1BnWdR/6qgPz/N0NL+oU+6A1rGG1i/V7O+ODH5ChcOAX66kmDuF5340gsg2vQHJ2XxMN
rur6ewwuGmmxutaHOy7uRRjRO0oo0xJgM6Og1+Xmdi4amSA49oY42NG+F+2FHu7R27Qvlk7HdH8G
i4IOhNKGyEyKXnqjiQkC4iBMf9360r5e3J+Q8kkRkpTuAAXtK66YOF9mSiPJTEdVqeq1qmvtzwDe
j3wkw3NgxnORNManOCeYJNCnFnzsW53CWVSFxWMS2G/e+yqYeOIWF6o6QuCmCNsBkmaPvKxmj+Ag
Uiy9pbvjVJsGDzKPNN+4ea2BD2nQQnUVLyPbldVMwBP2+fuRWBZVCJbDEqCiFQ3zpPG819b+XSDX
nS8DXZOETFN+TUIqJL32ZyK+VWezdaoxj2/I+Axf8zpD22KabMowP99Yl9B2GnK0QkfdCz57jxo6
L+b7xIR3KmSIhRaZrwL9+ba9kZV9XZ6mdroW8aux5GidqT2SVMODi5EQUGE+WEw9mifIVtQ/7NPS
SD0VK/FdXzwyPiqeOZv1WPb3kZhhC9jlszeR47QzZDOB2n4FSMr/Xe2YyGHbkyDkDxGkkTq2B0M7
ASURzPt7JrtVagKEH/73Uubi2kSYk5g+TycH3AXzPYlOa5fyunPXVM4aqSquflUoqWMqAGGH4305
ROiT4qqVolKp8mt1MJNys5Hywz2+FsXtitUCI9FttH363tzFYyMUAcBfxZg/FyfAhDrTou3snDhT
rNErHdffDKHnggr/GnWToIAmC2SrP5HvUseqXuIEVn7dN5ITRFpxU+qkIanC0bZ2V0ClDzOwee6h
hf/gripqzdrrxTzUwauafVMJV1Yi0tknNnmN2PRoilJHmhU5mqm6h8fXXIoEr5XKhl4DJX2PNBg4
bujV8B7Fm6H2OpS/n30gurNqbOToU6EYcUK3R+TdK+ih/eT43QrvPROidgKX+MQBj5KQmuM0nckk
wsQzHwlksjZbUTrj4simNX4fLlJXRCZ6Ot5dDuBpoKV80wjQmCPNcYDAzhTtQXHVvJlSOvr+4HDk
t4Vgszxo9aAoJOXa71g0BE/vJXsp6JicbGFD4a95oU+WL44ONZO1W+UTDIfsDgrAfbEUqqf9AIoE
9CYh0WWHMLE3/WgOP1lPLSh0YXhT5RKPdaYv4eTKlAQh88pDBvr9oQfcyVd4muITXfekvjGxbnTK
7WreqM4kIoG0PuNz9hgoRKYnpOqFDMqrTtd78VibK6ZeTIidEZni9zBzVBR/j07KxM6cnrhl3sJm
e9s5k25D4kff5YsdehctrxyaWKJl2L7P+1UTN+sPI8DPo58JtKt3dIW39okoeoIsA6lF9H1cym+Q
HmAJiOr10YTp8ep5EF7IMLehoCMkdyq0dWeLs+XY7SyBjkxHNdWItxCSAo17ltURLd0bk7Vba8Ug
riG8PwKPI3ZIFi85EI2kJ2RdrEKptcGsMYnqRg8CctgQe6g2zOTMzLJk0ZWDBnUyTPh5ndNMQn3c
Qjm6KAp7O+Wt1ktH3GXAMlRKbk7IZtYn00xnu/mntvkB4NcRoPiXU+0Rk8oHH+1JG4yJ69N5btWx
nt9I6GMhMqCY7hE06ra7lJ3F8VGiPhnJJX+eqZvK0a92oSpT61hzurbJFR0kAPmRokbaxNM/4Dh9
jL81q+913PxOkuakbz4cNFLmEauNBEwkRIUOmK18XHhXa+pTQy7mp9qYWtICGX4HEDyq1aRUGqNL
PFzJ80hYj/ncDsfcc8oksLU05yEJbgIr+TRq4K2ASJ1RpjghLV8lA3vqdFlo3Bm+20Y8YwgQSBnB
IMA3Gm3fOzhJvYQ8Hh3ocFlapIwzOdzSMikeen8rNN+Y9BAWE9BMozxoPl+ds1lSb2tIJG6Jh0wq
JBiBsoRl5NNLlNPNn27h/5L1A2pXFMVOOPzUzmPDhZ2pskc6cNHMfSJQnGcrQCL8xT9a2iOo8ckq
jU04BWRvz2LGDJjeqgGMxpVAl1sF71SGcaNfa3RsOe26CeJ68wyOqP+VUEAS2Of9S1ToantTvhma
oZ9VqK5h2yABnloMqsSJT2l7JSbRwCd1Vjfv0NrtKO6pCnItygWW200ZAgVkp4i6eju32a0f6gEM
pdIJYkABU4eyonsfpTpY64+Pf/k4kWUgHuoZmiOJElP48nR2CkNi12bO0fvJ9sku0bn2+2enUkAU
T3fPKOO04j8zubAuIZg48BpqhNlc7eTN1iZDUq3c2J8u5bQm6ix5WQM9Fk//yNuSne09fSwq+QZo
bx+CdBSWBez+lad8IUfx+JS9Lb0t5ROq3FcV08ksJTGKMe81X00Xz0xV+GLXdb1t/65NiIzwh47e
mUrPboau/q7lwoytSUgawuiHPHP5gDXTVxodCUjKbcmusyMFelwMb7AehsrN+LAxqQtSs6dD1lFg
kjYup+A4dlhL6PT82rWW7jBvcY/7nhLmg/zqLcw1QLtDBXW+tHpEyYlrJFpBzO5tt5HnnWrHfh2x
0CaOef8XXGiqo97a3VER3cbH2GABf4IL5tO3gNYTyrZGWFdL+9tc6IKV5+6lV+m8glNpcJl4Lwtr
BOFdxcYgixNyEpsH3NQZn+uGiB7i8dZTO6SkA1F3WEj78DKzEM2tf0t2vQmBQd0rV+SiXMyA6iNb
fFDR7km4qwSuKY/nMbkxjuxZBU8o9J+rg+jYDPDzF1/V2LDvIY6gBGvfuM/nEnqQXr+AcLpnqMlc
7eBdbonhJclUFyMSTR8LK9iu5z4utAN+FV4nM431HG7GudqOF/r1o5VvagaS/hwSsKL3/IznMOXE
OLkE6XHO3lhXz+Anfxo8s2j4DDwfTXIKRzFdXD5p/KKCQPtg+vGq1L9Opx0eNCVo/jwra7jrO/C0
yZmOkuVVupN1766tKcnG8bJg5RkVIeQTemlbIdAfUFwDKrARp2xqdQJc1EhO5wz2Gt7VbgaK+btI
8wa6xT6YfKy8DTKGTDaUfLlGIAXVQ6Yq0WlC/ueFFWbJ0Jc/GxL0N4eJkg0bkd08yGVf9l3h9rju
XGIz4IHEUG1KuZ0gGlcygkWcgkbkaqQUv3B5n2DapbmdR2b4I7UzMXAVxJIHyEjwhcKQnK31O8J3
k89Fg3HwtO2Ukq9oS+BOtpW+DGwrW3i3WXHbd9m2ZxeWd31Pdoxm53E18JMMC2FIeGrAIsqHJek/
jIFTx7wTczm77685lkql16mR4g8TbYHjioZ/CKhHQhCoZi3lbBdWjUGGH9f/0YuL3ym8+bXn/SMb
OaLMYhzgrCWN1w+P6UTvO/lC/6Hf7nsgScncoCrTKlPTLdncgVpyLRVO6QjtL10Vk85Lps/i7JLW
qDivAgr8eSQT+Y+Zmjr34aPtKs+F1uINff1iH5BETj08xalaahMq0WLXzKfrtjKH8KB2HBdWByl6
/9m93xCb18yl1UgsYNgW2yQu4RJBDyhWH8lT2FWYeM3kDk5rxWLOKxQZpFx7LMGCBc82nMeNAE/Q
D0zWYAzpySkPiGre8BdLRplEdN+MaRe2Pk2eu+mSM25IqvbAb8wZYQ2w4qqSf6EI/HKba75XCoZT
6DyKdOS7s9F5r4dYVNvLRFAkfgnuQB+srwbOpKQPqXiw0ZfaF+WSlg2UPO0XPfUHvrvWNEB3IPck
5K9PP6Sr7uasCzwR1E/laFlqjigDIh/I1P+qLonlG/3usYtPULn8wv7NrSrHPPqczzO9d0gBOp/i
4wi263th7qsZgm73/Q5z3DHmM4pkjnhJFvUsv4gbjEw/LZZk+Sm5acczmXJICb9x+RAyKtF4wcLd
S4ogAiH8NcnAf7sMl0Tj+lRR3HdP5HBe1PETgLcg9or5K5JWQtT3PJ4OFgZsySaiRtTjklLR2xM0
L+2SvC1Y0bleIpyTDab+aHExqcbu60wE0VH8qo7DAa72+INWaRMIXAQlfIOXKSh6Kg7cEfSbFUx8
D13lbakcTJA3TwnvE9AeBv3AV2mAtPVVjRpsF90mzgqEQeBEM71pH5FSVJUktjdF7RAucR7vEiHS
yfL5NEGDpCETenAtkSPCiwWKc3Uz4FoG05+ZvyAPXa28ra0+eJGPrpWffqeQ3d7+yjvJp0DoX1t8
t2Z1p3h79kyVUQpl9jFs9XPWPgiIFCKa/lmmwVjl3yo9Uzl+zsvSAWmSvZ/UfcO07vW4y1JCZMTp
KtfvouxAEWrMUFf0UIfKW5nc6q2sZOMgXZfftaNPrTktI33EaXhmFinNeDBFqE3ydrBrf2p3gF9x
tjqcqcIsGH6wGvW7Ojkp/P4mbubGgZVGYNyWigyudJRF+rbVw9kBDFkOJXjgRle+4bxYD7f0F8ED
vrl/caPmXn69GCDUTjICkZXnqlAk+/NHplKHZoNBgffnfWNPJZoI8F+GcSIb7seRmCXPG0ViEBl7
DeS3xSco9cZvoZofcfwFFGR2kDIqRtfjXJ6DQtmwWWDCNeOeHRcxNP9gRaFRTnCFt9JpZxm2cNSv
03ffxUn/8JxoyfDv+ZL+0TdFIMMEeaSBVQ3oTJmSLX2B8zuPO/cW7+usZ9GsBhTlpp6QCMvW+zoX
i93nbemt+w81EsMi3vs97xKg7SqNfmPu8Jw3tIw2qVE3QoKCGQiYTUBSI89CCI2wb1zER8brOyed
Zla4cImTWCjEGDiefQddZlSqI1ghkRgGYy9A+JTc1t4jhulydt/87TziX8Se0RYYBjqzKM52mn+E
rYXNJ51d455BNsXonG3Z9PoFGDUygnIfJ0fZdnxDdQ4NdCMS6Z3j5v/G5xun9QamWDAHPYrgF7sO
DhwDqnUO2OOiGD5dQQMQxiz1nItwbt3xFWDYetoxX1XInnk1JPuImzx9CUkFDjoPj02IwM6lKWIv
70LXeUeyFjMO4ngY72YMIqFYI5A/STaSxw+QWtADz6V487PHPgMwmBCkg2aR5Qz3i8Lttw+/98Mf
AZ2VKM6n5uxahkXGmLnPvZl9j2ssPo5Q6mCPP3OxF2I1ccQw2auQAJ7YiMaJDUGllnGb/aRZwdZP
EXPJfpkfp6oq0Ol0JSWQiJ3FVMUryXM/OrPkaeUhyzHm/x7EwUBp58FHWy3rep2kvv3O/3Fp8pwe
2+N6oky5gILDdb1lmlFnbWuyLNi+8LJIU8ehnF2n0RRLKEjSULORJY2R5YqwFXRc3j6z+SlfzQXU
yrVGHf+0OxsrqifkwHAivG3IcdKwOBZWztyYdLluH8Dq/E8wZtgS3vO8mfjD8MSZcj333L0zxzTC
7c0Js+37sT82d4kTgJnExlmCSL7hPFfNYGh3G11m2QPKGB3owRY778TCA9vnHR7kunA/lL6FMDJn
bePYayDwGAN/UU4Qe8GFqsrI0K16pOODctYw/3Pim03voEJvmRgs/C0vQhtr1NbHDFDI7sqyz/sN
mT1ZrTJHyOlL/cjZ/qyRwtEtByK8KWjjaQYfbk4xoLGRas2Szlqi58310oaGBDMRRtjl8FMOSr/a
GDxFRd6EdbGIVncmJHuy/h/UZn+TyluSYTKlRQRI2xdHeb93jeCTkG2k0LRTjlmGsEjUR7phWW1g
78q6WhHO0FYb3JfCc5EkcyJ5Ng8+4mAsg8hiRSMdvLfrsYneGm/vpF2EshZwc4J1WfhpGz0JouCA
chPTt3MDMNCkz43xnb9ziYapXArCAyM3IoIQ8lZr3PvbWI+lGFMO+ffzPHmuWyGIWEwKvRKDXvfi
h/v8p4wC6CXF4rX037dRR0TZHY5wf57z3Y9oB3VCM6Y/ex130n168W+UBteSwxXHQkW4H+PsGNRg
HKIVrnewXH5BB/qZBVU9O5d7goiVmCmywJDmelYa5Ul1Lzn1X0uZa/tvMRg4/JNCF2hC5VNrDoEr
xmbO17+cuo5iW89zqEoOAlgIYWUZKOghZpyKHhGnUvoftI92hXz8I4cTdqcAXK0/ZWfbMQV8T6YA
jXORmR6bph7YiTUt47mILpT/pb4VSKVSZBFhO5+uHlk1TVP2aJ2dhYPSjMUo+bR5Bj+vrG8+Oz0l
J+DPKXfteb5SsmxwW4Eo32LDFxwoESB0V28uD1ep0o/TLB1Cl+53IVzhJh47i6tUDF7+EumKdM+D
2byY3bFbIdPprlbTH2DuxHexAYfTkteyGYloiytSd1xe4cnRnkX49GK3e4/cZomF7TJ8FMGiZaEY
3XsQw7mfhKBT+3i2oV7x6lKgLPnMjwVEkzqyysW0Y8ki5+y4Wgi8ww8OdM497k9XXeLbBn2Nc1nU
HGZ7QNSpTxP8PnELxqyqCWkVcFgPs9i4QQUeclnsXkbdXnmQhEQXS5tegfrQjaPzaeF2N51BiM65
CIyB9x2H4DxB7wob2AvSGMRBdyBDn3YevSv68Gb7WZZio8tZ8TspywK6TaeoX/NwGej+ikPTIhT8
1O3OXySEyB8uyOzn9cJIXd7wP0OoJWpBYgOKM/QPzH8RxMehf2I7Xtmu3XZosdYx4SetjMX46OVw
oqamIjCMpH+D/5Ww9K10dqxlMc4IwmVKmkl3HL62yYuMkWCOqKNjrM5nEqf2i4SQWED9GctXBjAY
HpxuoCSqMVnaficupsP0usZ/3hqweMI8nDrIxisFyQ7vhX4sTuDGh3vsYKC3TSgCf+E+PU3pLaW9
jmhHgoeRNZLiiwtTzR8PkUyc1iaZ3GN0JhFaBuHQaesIbpjxoyl1yTvwykW/cSoiI8KsTesOX3M+
u1C1Eh8MKcVtNRfF1Akbkvg8G4pIMELfmupf07d5iB5kykLJOSQ75iL/gg2xu9/CUcdOnUDHtOvp
7zv+4nOv9HtuUYNwmQt2US1aNUjzqMdWCmZG6Rx3yMf2+ehUM4wLF7ViDwG7qJ9GbQXcrkiufeX4
z1G19rLlzpj22Ko2RAaqnW1RG5cMr9OSlmnAggEHdQWUC4s0A/Wg2iVZyJMlX8Jwja42zZK2/LgN
L2v0RwVPIJsEe6xmhkjOFE4DGtTJbz2K7codwW9tKqgpJgcWBDNWr4v20YiQMsZx7pn1F3xnPiRA
z4uPyYF+FHjkXMK2aBrtw8dG88DL887LHqAxhTxypqsk/oTZVXaxItofcSHN5gOSamuuNxcos3eN
PpNEC1g3Tgv5qfT97wYVom22oKU+RFzI0/LspDDogrFREHWyE7HaUtLgZs7W5/s7vHHDu/NyYcWA
aXiJ8KlDj8iHnmLkkr3b+7Za+RxNELqzpX/qdpYW98J4enRuaUv5REM42ll4ZgyLUsmL9L2G7H/l
dlNQ5B+3X6Oaghs3tV5XyRu25PcoIriXCygMHcmNzRouyWIwsAiAquOi+Jo46ZAVTMafNgo+XAhz
9tcDZEvzdj5u8IqK4dLwfexugktK7FQVALQZFWPMPCg5JdGhHJV0hddg7pNnXSF+7pGfHy3GUo9e
7sY9WZp7NvZBkvf94YFjIFsd54yN5XFXFDuU6ebdO1nLZLTxxHtCBihIKCikB2IWeEv5WFqc39z3
C8Cle45mKd0b634MaFXp8kXtJLQMO+E63gU3oFqbwrwZDmzSoMDmjswgUT5aqIZgDUN8zXi37Q7M
CKBWbLEaDd+GqCEAm67uRHaqdtbOpCfPUYbX67WGUUWTL1AeuriRN8/XwcXNUf2655zV773dX/ZH
vrOwZWYRYIG6ZQTLi7TohNZ2s6Q4ns4Eo+fxq0ncduuxlGHyHgPRBQnyc+RoeJkyQNNo1i0EhM3F
euEW6+HTP8MbHcTqgrn3RDkDWYeqhJ2v2COdUSF5HLwS5g8zHtAMpINcx5NUSDZCMOfpu7b4yDjA
Ig8gRxs7UKFwAG2D0pluyIPq4q6YV80OL59qenkr7PRsG/Ytvrr+uBYzpPzCtkdqCZqr672Sc2LW
0tD+meaoqiU/UyhZkwUd92NDLOQhWDxSFwMQ9gf6j03QkvRb7k9tLJWTkfrsOKeV0QUUmnwvUdjS
k4vOly0JJSiWAZtjnD2Gh+cWeBAnqAwLhoLVG02IclzVPl0gfCvbPUPDmgZvIU1cvVI0g8d6eVIR
K/XJAsckNnLmXHUvK2eebpmSYoQI5hjrY0rAuRkrKgmT9sRBea4g/wGmd5gSushc18Ucxz2/okye
luTUafcCN9jRdp5I7Uhfj1YdZozLORaDH8FRkSvI/0hgNI1snv+wXhQLg1yxVIU0VTSiK3mdN38w
Ub/xyY0dj8uuf8nUfhcRk22vuvThpnZHXHvEmKaLdfJ/vYEqm1XEKcotTttaJJzaK6s4IRJ2ZtTL
NDjr+CAHmyRRlbsEAuHRWDqD8CyiCwmPFmSD2Ar9iHzs4FsTVKJskSvx5v/Gy2n49URjAxlKAL9I
/IC8O79nDAIQn77Otl7+D62J1N6zWXiT/nF9PVbLKJzGDDvxjly02qHwifjNayxqy7XNsP0TFNAF
o3X8M8Bo2qSjR1xnsA1GvFCrwBA/5xjuZ+Y67Xe/YDNvX9pxTz9pWBj5Lyl3Cp/CROOqG2aP6ErJ
DvNsWDpngrjXq4w6ShUOiVeGgb1hlpDa1XZpGPB1FYwAiilj8VBhYugenYUWMjROQAe0AbNkU5OG
SP8U2wqgnt+eQ6MAYXjajTcGTlD4z6VVIOzUQCWVcNr5s+CUB4QVwGev3WX+xUDoZByIVViPY8e7
1e8BV1u4mA/r5BUv2Wcr916lW3rvLhQE3Lb2WjQ574piGvCH5ffzV8r3BOTSzG1eIlxJArq6QKbi
Yo76ANPfu0VrMDBWgU+J35HoLH/YtqDwvztEyKID0mMWMa0h4BAKcN7MEks93mRkE6zr2rSBn3Fi
Z7/3q0i+8ezNTdoOWrePyj3YMd4RySSQIzwLedxqB6L7xhKAHWt0etkoqSUwS0fwo8q+DeWLL1Rk
kUnhIyLCTuF+ooorXvODDT15JfLvEdGO7RQCBp7n9PLDjhxoa9HrWlqexcSVsZxMJ7VX0EfGN5E5
ptoevz+p8o3m0QYtTmiNh5j9hKjhyOcUOKWfqI3qFXGS1znZLRmx5CdKS0F6iFSEXIR7WJfHbjzB
E8Ses2cMyV5K7TUunhNCtugFEr9U87X5/HPkemFGPh7nEzzqMfqMRA07mLr42b4DRRne6A1OtV0Z
JEgnhE20yX9ltnj1y8ksul4Mvapqe2pejINVr9in7PGeygXy3RJtsWG5y6bDPhcjVMFDrJ57iYb0
Wyw43j7XSGPQ6+ytpP+E0lWJdJWYaHi/PdKzc3otJYvl9y1HT8sCto0R3sA35kooD+UZe2NYyBks
P/o9ZTswS20xzuS8njf/Y3i6oSBgWB/CyeBB260B+lyzgmL//PJp6DOaY58R7eWgR8eHvTd0tTlY
PaMjAs2ve7TQqrvrqakw0Bcppz/KL9IOQdAF784Wls+HtCRR3PUsyRUzACIQp6pQXlkreAYZcf6X
06Gm0qwg+oqMkMeXklhtZ0HPhhhiUww2l/k/+6PPDfamlMT5ig6LNNg9X0uYdbyRW8O+KR2pieaG
0h3ML+4FChNPQb8DKAhshCf+IYoIO94HtY2xufZSEWpl8C0v20kCWRo6PQ8khPFJR5QE+2BJrxYY
NsGmPQPHv/b/0XpEJWP7UJRiysKuyRN7GKZQr4jqYZ9m7okFDRIwL72xfztN1mqB1xwXlb8aP9jg
LCVJWChICIUi8xWHRpwVHMnDcysnY8LjpjnINpWuQ7j7Uc6QO6XK+By5+GAGRJwU0AFRnLDjalvA
fM8Qrrtq22fMmcLxorlyWSrF5tHstdbf7dFRG7SaBpfcLriQePZm2NuLG/T+A98cJPcKYmzau3B9
LxaiPyKgrbLFfMTKSUvpcAMr/ql/SYSxN71cHHPWtbvxAG6G+Rmt8LUHOBTd3+Q+fwVCf5TfBwed
nN8U6PFt6g4JkhpuzlssYbWwmpavsiGRjyyTfWF5MyteuPwkmp9kcdXxn+bYjHrsAyDYu4IULWui
c2XOL4brJlfXOTw1SeMLe+Zei5313qyiqI58XVjYoHe8wfJWczb/gOzOyIbn5HtLuPQw93NZ7Weo
wmBPODSkAxi2vC6v/0Bn02mEdJrHt/obsEycFq6eAEsntRHh0m1GlbagOhc3f6r8d4X2bPM7ADhO
PPaEJ82TWAVyO9FqVT4r9bxtAwFw95H1NsVMyW3withN0q/DuiOgKBbiiBlgKVl9SWjjH+X99sTM
2sqPCSrge4DXX+xmyiUOSOE72w0E4QTv/vCsWmdUCGPSwcxVUrIeZDMWUp1zDtfjNbcRSqZOr1zy
lhTEX8hxFlitmf08WRN2PVd3fkH6CLFlire/Eg7X77UaeNog0PycG/T3ylgKiuBFt1VnE7JT8zZP
0veZHXFrQ8B7eCy3y3ep3w6bmNVtcEIR9tezWKSUz7nruX7W8Ir9p1MPO2Ue5ooHRnxFCFVcV4nA
U4LF8LSsjqKPRI6BDilUXTBP7LUTLxIA6QBGgU92N6DqQFbbpffQCQMi8gURbTOS7Hl7cE4VTSZv
+4ZF7KooGdTxz2o1uR6a0wEKisPcoewcg9Pjz4QZAt2RVDy6e8Q9Zhsozt3cUdiXr7XQZvhew+4k
rdqmIZgoHFnnDfSokkVPH0qzRupxR5Dltk2swmCjVzU7OVOCYon0JR1/MXOEYAUldPcH7OXI+jxY
xQzN+ojrpwTulsH8WFBU3NHn4/uhiUonP8yXVV0oUUj7bGwFazrqCEXyk+MI+/b3Le7Pf4bo/KMf
8LHBkW9VCscDqY0Ip0UVKcTQDh5OwxwM7Ywf7J/c3aKIB3m+KYBAKuMe2N8aUawhJDmSDl2nipPj
ntnWN4HDK9MqfHqWdUbDh+ptIqL5tnDPcx49FHe46LdmPvmUq1TYJGiY7VoR21g4jkvsGS6Vsc9G
Qs3xopCCfuv703mUETQJwbdOGFUOfBgYPwHR/uG2UGafuMMsiSPANaAMwKx+wnoE//jK/ulTc4e8
IP1eybur9HR3wi0jkleFVyjFwr6grbbqHX/Tbl4lu++LCplG9jH4+X0PyyG/1B5XLX4hxY1nrWLi
UKFu+CR9XrUQaJr0BWQ4dixcKH05uGlcMJ/l4ytf0fXCJ9K3ZBfLTyggGgztYsZo2ynlT0iDxji4
EJ+PAhMfiaiDRbbDJlSpRjJbhO59ucPfgS3oxSIkI9CobNEwiqJcZH1GnFEEF96aJWr10iATr1G6
QsYjRPUBqUMt2h9L7f+Y7Sc3tXzZ8K220fkS4BJE3WiwN5sBHYqDLjqDPJnJ0bGK+i2AKiMDXfC9
2oifksTAKdPOy0wZFt23evAtMqcp9N+c65Kxi4a/FYZSZNpA9YFaG2uf44CWHKwrqf/1HbSVYsbC
iLHgIBLBy8D4xBJfnIl3Bvy9UBN91HNK7jdOwG28FxBT4MsJMoUD6QIBOUTm4Dq2IgV15UT21Nv/
RvyldCl41dAMTsNbpjIRBToAaGtv2FJancmW+YPGLq/lmtrGIgqknoQLtXE9NCq1sr6B6KJjvlaB
o+FePPpDPsKFLXcEACnwgsAlN3KDQNG/vy66UBAz/wsDullh4SJMUPtMbmKTlehX3Oyho1Uk1d5J
J0gigkkM8vK5QgoBX+P7guA/tlWDBtWMv4hbjNR04JqyUzO8mQXlQDhyhjhUnUzIwRpi4jCfGB1p
O5XoZS3GhNe/7pvBWNJM6qK7mG87BCi/TAI5jsMTYn3VO14MhELDZAqVj4m3v6ksIP0dmO0b1zRp
pDDchRkBe07q3AR9wf3jJPRxUHisO45SovDtKfZuG2RaDdGy0wNBkN9i/r7LZH3yjCrxKT0Zkmrm
k6G3H6MqYCzwAztkdWq2jI1Dy2ilOgwdP1tGoysa3bgncWOH93eFfO9ekqedNrlG8ZO9actZRl05
btri7OqZRifaBmXcO1fsXxOJLvLjfynBTgRMxM85DYrqC44AlIFJa1aT5fQMj1itZAOQq1whHhaI
0nf2gM71UkwxJtdU3HpylqCF6ETfA+rSJbmeDs9KIxNXn3v4p9IWmsilS1dAcWyX8K+91M31JRTv
T0um55stqdtEYmgMAJPK1ner4aWiXS2ZN8mwbfwmriZBd7hvwkKQ/GGCJrFU4Xjri4t5GnhhK+wm
rkm1Y5XzNZjkfMERU3f7wC8w3Zl36Rh2G7Plc+CJ+AqdjhhB37cpejFBsQkGzzGiiEG6zHmxZ9TU
e9NtWGKz7orlCx1KOkFdhIwuPqE=
`protect end_protected
