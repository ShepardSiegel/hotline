`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oLYMuO3QbaPqvPo9lWdtLXs47ZD6oW85y1YgWUTRMKHsL/pBiVuMLbzsQAOzm2lfaiPpPQOvBiY1
JXjHaBxiKg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eSsYQjQ/8amMriWYax0+jNGLvtQgXbTUwshP7x/eJqGh+tTiMr3z2Gb9EuUHR/RG8eIN2Y6zRaLI
bXq76Sis09QU52elKCPTZaP34XJeM/6B5Mjy748jAyHAGMppwH9/630vNJMYrrN5TDKA+xNRxd1f
F/rQdqWM26WZ8iaZYr4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CgkhH6pIcCyP8qYyqU78Jby545qoI8zzTLpLubCDQU8zt/pD1whT5GixdFFS3ykeINY8dxYgeoCF
oKcqN7pGZhFwHiBjq1JOtf+pjPJ7st8oVHIOVJ5715gxg9eEQblDfNAsdUXhbH8N2/gWpVkicYD9
wbr3BnjFGcjyXPBiEMY3V63ZREdSqL8ASwQs/L/ixYFOLeLSu5wDUFy3wVVJKdhlHirGIX/IiPD4
D3QLK3St33raJUqYdyxU0Q+8Yj27PZN+e39zZNsszoffBXGVzzQdH5vHcml8ZIehVl97ua5pBqs0
5Cc+dDJos2IRdPoki6/NhCPDXaWniOJQxOBHQA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LSkjiliz1ZShAV7YZ3brkqeGIDxplunqNCf7tjw6U7zHzu3/kdV8wRUEgstT3nlU6JTs0ulaFMf4
UvdS7rDv65/D/JauunRWhwchZnYlJPQHndOkQn65/PGjsXkYT5y+EtWMmrx9lKoo3sVxnU+GeEAG
aoCzwTsExuxEqB53Whg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Skhg8AscuVeaFq8twTbyiZRoQwwBjjJhSTcH/vkzNvBvB43nqHacydB9fhEZuatMbi8VzOj0OUSQ
WtJGhkHqyqX6qpTdPV1UtG5ybXm96K6Xp5IHnO+XQjpHN13ZaxhgPppjluTpC+tvuV1fCXyPRfEg
GgVC2PkMPT8Kq4DIXREpo2rKya3PWOhzYFU5feCn2gfwqeZEhK8GOmC/85PHNMFuMvBCGJeci2if
IsIlOyq343NQdlr1axjCOE9yBcylb6ZXLDnYVoeHB4vg4AaQ56OnHn2N2jwO+Cj3rToaCrJ9lCuH
0vh8CvYfIO5hRoi0BInNk17of6BAs745dW6fAQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10384)
`protect data_block
gXhBte6vN7XcX4XWpQztML5JRO5x9KQ2DdBj7gzHskpnWOXvFTQOycb1A6HOZkM8jo/i6fwKdTLf
tCDyMGWuaUd9zy07gYX7XicX00HSu0MlIU41Kzj2Ovt9o+yRIuN2airdnkunU+vX0HY7IdV93uSO
EbvPkHezGxJpx/ODJigru1qPSa39u004FWnvaBPGz+V/B0CyIfWDTz2D7uT3dCw+FT96XddwNXoh
kp8GdK0ksI+tH65+fght/z4NEe8R3LL3NRANhrM42HvbZvIGLuxXpjImiJslGTYUwyaJxnzwX9Ed
Mn1tRE/T4N92+lPNcaftZD3yUgCaQHm6zaY1lwd8+SQ4U9wCiMc/rAUkMSLjELtp1GRvzNv0BkwJ
vV44NnMGtMPBYkb1EoEpc/qEdg/Scn3C4iue9wVAG9KoJBWDCzlmtow+N24Pk99lcY1uIGE5n8A+
++QVmsWDA4lbsG0klnyRPr92m0bLNMG/1H3Wta5WnZquuI4jTV8dyYgW/5ZYUV552tEoifVd68rM
guUQBe/U4MdPW7ufSfD6I2wt3AEFNqXMKH1ek6teeH87wyAUknF9q8fHXzM/+3tK9YPf3kzaZwIY
MHH1sl0cQx3AkfeHxYYChvnN3RCoqBTQUn+HCVu15mXh1mUtlYwM7jUBExyxDk2ICoNjoMmLI1JN
lxNg4dd6TW/x9VZoItdlsYBk6oSO0U7/fGAgMIhwOzg1yvmYJEsBg6n2+jBZIL6fzFhbWdtQGeh7
EgLrQVYzwmkTu5owOKN6JWYOyPgQQ/vwbjxzDj6H79rHc6DzWf1ib9qnIQSblsVRH34FmxdcImlb
U9gdL4y4IJ02sytETM2wKMd2gxtOUwqUG9L/yrLL8YCIXe9D0iuWDdtJIiTSgLsBss9T4mNY+EHt
Jx62rVcEWQn2rCc7nGzueCnbE36IaeZDtXOsOWeV7WQaa1MFugQSD2hYxlMPDOQo0IaZ2NAaYTfV
wStUfl/2u0JgK4nYCMjZq4tMVo29obEnP5gpyBhNMaOAV0mMYx756wCX/sNiYBbXt5cTISf4Dext
YPZy2sRooEF1C9Tc4AoqzQNPiebDCpYo75mIHahLYlqcMK/9Bop3IvDZBXADIpBT6LBe5Qfp84RR
WjyMbElYnAJsLylHNonSk5N9mJBhE8aw4ez0jrQbkBTLKJnsOpj3AfOQ29P0l7HmpNn/8rOM3QKa
9Jff8JzvwAVu7x7NrUyZYgs5pChCkGJiFjmTdQCI4clUI+FB+BMBf+vBPdQRhQlGQsvWN2FA8BeE
n98u/02vgqU27oz6YsAH3qSXTB1HfqjAApzxFlmHcF7UVkTajEQ4FJSudFpbMqVEra26w88cT704
aEtcg5rhtUwhOQp/+ZchUi6IvEtn368ARnMFf/OU4UoTpWQbrZO+D2wQDmA9yfqGFMULFGiK1Gdm
EmIVu+D5a60vLsRb1s/hG/b7JQyHS909XrIadiis6t8EapM46r7W0LodZUNlGj6j2rfmcyLEg1vw
f/GskeUfRfR5lR2KZCqxdyzWwRmP1pWtyxLEjaXB/h40LM38Ig4rOPUFp7HMVbPMcf23jXi/eMmd
7Fm8A0K+reFMWssa9zg6qE5ePGpb55VOulok8jpKgaXu4G/aPemlUsRJMjVwq+uno2yg0sUg58qS
eJq5aSNy28DZGWwhjzH24SHIt/zbUAa5qzL1jcPQXlQSsH+f4TOyi7xByC2TZ2TebPb6A26RZMp8
r0hOrtPq+hrRAlFw9TB8G0OSlzpbeFLUKEc9eSJnHX7f1gPTb7HcFrXyjXqy+WzSCPKb5bPX2LWI
iVXgpbdjzeAD5sCmncgH3Bc8RzqCMcUm079zonLGvIfu/itWJ69JQmk9bVsltTyKS9v1NTbTXOFl
qv/jxwUJBOFd9ZJKS+CH6gHXLyv5aiEmQA52avkhDZ1ibWT4Nmmd/n7BwiuQq1MR/zypc8WsS7jN
NHMAqDTJ9PTEdgEWjYXkz+5iCK7whstdtGznW0PRK042j/GMagHdKx/21apt33GU0p3A723dm7R0
ugopmZucE/b3j8Qw7ZyvaqhIyGutsX59B2jLn8y97KDCAEkTBq6xFKEdmQ+XfwZWUMIs5ktlVa1+
/BLs6GP6CPIkKik1pPKz9b8/qg4L8SEPA7YXTVlJpQFWk02t1RXaGxlNYmoHcpWgZa2K67pPem/j
Gloc2qg8jU5qvtvw4ixmqDoR72ppXq4MntZBMBUv94SgEXe3jFUZRySGAQsCFPp9oLkBuKDIfD5w
fclreNOlO4876cSwam4tjUi85gYlEKtNLZewXgv/wA4Bf1J3tDSu7FOii/OOk2OaWbaHAVPJ9EuX
ZaWqv0P4GGktpBGJwqsaF34k882JGUzsVFIDnX3kgTtuLQHmhCmVaD51cZclxN/h8qWB4VSd5g9I
s4+wuj6FW3qw06I8Bcuc/VAi5FLno1tJBPniDcLf+B2KQNVL1uJ9VYyzKyeLNzwdL1kyqN/6IcUI
C6UrFj+omU22PP4+Bw24CS94kkufEv89s9k9RYj9N/7amcbXxqNvdhldxYdzuMBlIn/MFqF8+jHr
7mcjTbEq2mLxCxHUeZLEP3WwY6q0bhHszGKdKmi18w9UJFt0goeVEi1bSDyuzhjz7nLmlnvrnVGJ
LnFrhQWmuEQSRs1VIcVQHHFVwMVQlzXpocAeIxJehqSjj3vUs/nOFWk+lmr8panO56B9TBXFG7dK
zTl/g+MpSH+Sf2bmbQKQ0Jxi1Mho9sj6Jp75B2ZzMfGo/lciVwDn9dNoS7JShg5i20+dUfI6OysG
Si/zAsIz7pAgI984KLyuYkGa1IQQebnQwD+uHa6SkKLct2SADiEfIPBwDznEhskdOxkLl6jojapi
saCpGzFQL/ZNczZzdfN6yp61dhgWZxivexgF+UjjaFy9ScF4qtZXfnTzEwdXdUBlNTCj5+BmvijW
kOrDGgfPtq6Yq2lT8DOAubkd1acQu1B72L6i1wbbRdbmqwfLa2Havlicql8sR6ww2LmDu64OEo8n
B5NriXZvq5UiKc+JSPmt5IFxglffWJA32FpEzQ8lhyBF0xfeBrcHbcFd2AJ+z4T3v/pOdr54Ra6s
yS5hHqJomG6rBmS4qG/G1Ny5T8IagtdBPHkLnHbi89/HU2bGs+B72Soze6efDOYSG2RJEWApHU5p
zDdN1CSKKIo/nLbwQFDkB5dsuxkgL10sXwBQCogEwkOlNIe4FFNA8sExwBT3PAPc4B5vB3ePL0D5
iYU7FP23XQsO9u4YQdFc70sQc8SaMWjPvItZ2LuRc0a/jGKh7ajxJL1m8y0gGuD4Qbt1LQcbmMvv
hVKPt88O6efQUgofOz3FNTNMPZq28j8r9twqY/nJOg92aGRoA5uS3OAkA69ShAEl/E7+oRRiOmLp
22mtgzJ5rv6SPEbWhVDJ3mmaD1LB4snf/5wY04KLXGtP9i5jlty+dtm3sGLheHUTLcY+WyxlXlY2
rBRdoG+SaQRYRwqqT/SKwI4QPR245ORW3Y9P3rpGUo2NYV71c5fp2wNh+jOf4TzmOLxc4rzkQFtn
eMxZdXf3CQd+v6XzUVoAFtedNNwGHljhKZotisxrZk9uKLPEInkERvkkATkoS4hm4n5NuGbbIVZp
f/g9ESfqA7oomW14VNe74bagp51uddvSpobihO43vROCguQydv6KZgZieTbcLMLWLGj32XwrPHng
5FA6voZzgm9tDPyAfmR4v/XY7sEFdMo2cDws0yhPTkZzw/MFKV4VTr33G9WKLCe+KC3EYk2GS2X5
TK4VJ11ROZObg2KDVOuJ0jKjtfcw3f8cjekJMyZowrputN7r1jC1C61c9gsTLe9EKMUupWfHva/W
7SOA2EiM4gbc6NRlC8NItAc3DR1YikBOo00iUXkdEzuDuCdCPj1k5g1/9EB2Ll9suY4FwtUpw+Zh
1PvDzxX1paVnuNtEiJpPuyVp60T1WC0/Lt3CfSKCNDPtXmyaXRdYoEKzQwfnAW2Acurkb8QGmDrI
36yS29AFvKOfS/QfKb3kJ5W0TewHWOycQtaAFa3akFqO/T/PZ+ejH0e8MI0zyhsSbK0azZMhZiVj
r0xNID46qQ64Xt7jrk0CQI7dpAks8+N1LocczBhJemXj8wkkPD19A5PuGT3B+Rs8YsvU+yyMWXY+
CzqEJ95oPyW3ihJ85sCDieFywsV3BLGPjJX+8eS4BOUrVbwtCY7JYbp/vaWIrgsncgIZoupd48Xa
5IvhNWknW7qykiHrkk3otLvEfEk9rSuAt6azJcnFhe99NmFb5xo5Yx1jkEYn759IRXXuQP8sJC+9
69/e02JNBuKgHmha3kjAFE+KAjWbplwXXf3kfiaSFVp1DUOQweG9WUODIRmntRI+eC43VSyYpaJy
z4DxOBWsv7ahb2EKwWq4d2pVbICoDsZTs8mBjrjJ503NXdlP9ga0MaLHjfGJlnWD5pjTN2/ZStvs
TyqJjKnCOgv4MVnCaxfH8tygytv8LK5WDwoHj9tKyeIsod5yXpkkguY5bwdco4ctAqBcLCjI9Mr0
nX3ROOs6XFI0IL0R0B9YvbByZQX0iBbPwVuAj4VHh4Txklcitv8NjOeHWqbt++ZBbU/SEhR81p5M
d8dQUOg03VaxSKYbs73uhmggqnjpFdz+EsPNwi2p6kCBV5rqdPTbuKXZkF3se9N9Tayae96WhiM5
N6T5V9LUsTSpLAwBCnWJQx5pLR31Doxfx+/RIV2nifZ8gK5E/JqgxXBdP7fNf0/mtZoaoj4M5KxK
dd3AgYHZG4fg4tblmECzLHYuIlhkqxVgD6c4xhs66MYKkghMizJi1qlS8TcM04FJ3X0Hv4DdohyE
1BixnIg6GTowp9p+9adwF22HhHZW8V+lOyw+aBFI9RTUBvFEOP1Xk6d0waIz66GpaszYJS9BUA6S
xARq1OUkHhI8bv5e6VT9s3uope6SaHopWg4OIZ7yOzkMpCYDqxLdPMXI+aVDEDG4bltfCRalafYN
SkPi/GDu/kZ0R6tCwOc+aglAbmojeyYDxTYI/lCdXYG14P07gptMcP7ZEPaUgapjIwkZ2+vxfrZ5
eWkdJ+2GXJcsWEz6ZXYcrhYk531we3LqSyx1QBG7bX28zqkB5wc67Mss//NlUQKzgGnjtGqr5dZU
8gRWf26RMMhL/OG1qlNy9vpr7k4Nu45lN3K1C2bGSCsqC4lZSfqor9fG4kzbnMUP9l5fZT6X4a29
2OFegJ1nOj3ys7liAQrXZsf9jTOYIaUiwMAOmJpTitDJdbPVItgmWdQs5fSRRhEv6H8Y9xfRQfzG
ovLl3y2EiPGdXBtGH2CE56nGLocTt8oX3IKl5gwxCjDuqsLfqdIkbbsc1HHi/aRPToRJsyszDas+
YJ5K+mWut1Pr2TLrMIY6eXeDvSTISjsxUmoAP7oVNAOdTX1VkGjlekjP25oC6S/Z5Qw9k52NCUtj
pvcQVVz34n8zxMBJkbHRmWEpOjjTRnE0e9nIxM1zuJOKGOfQVs404sy7G1vWLMLN39hw+0qUotcT
EUGtINuD8d4bfnOvev82qfCUrvcU38AwGc5Peak6tQX9yIofAkxhQWesFusjbAJ0vskUbPYlZ2j/
am7IY2o6x//PL/8vIuTdi5cVt5v6QPv6AI09fUu9cpEpt0MccL70BMdHsgHEoZ2f3O6HecO55vEx
AT+3xajYyE+PIATMO+do7d+1MUi6CqZh8HjucU2Usyq3o/AXWQqysUb0XxtsMYG5xnBzxjVuImN5
cYTmHDz0rEtBztFYBjFa5VMqCs6NG+KbncndFb7FwP1G9BStUFGcCtTqjJxL0Il6ZU/zsZrovbjq
v4gbNzVI9Yj5SxS7nMhvy5Lx+N7oi9PFcboemExvvVZgNl37CyqP3BhIK9FqXdG4mvxx3RXQsNzY
yDDTpSw3YfsfvzGlqE2Ru7STQQkQCq50VE5XNWaODtKgskcD1TVl/yuCmBwEXnUuHHpgKn+vAb6C
5n0s874YgM/QXeP7qMiE6Z8VkA8zj93k/eVDkfy0u7hSYUxxb07MHji0Zm6GfwQhX3oQlvYFGqyV
1mUXLrs1l7w6QVCo6abSGFCuA0LzWzOyusKOa8czzwiwcEnDycB2JF0K8uadS0RcteN9vfgdEMlF
TA1EcK+AciT3szphqTW+ZIBKWP4LiCi+3YLY4iEJafzcc72/MpWxlQeGXw1deOGtg8hos6lra4wu
L4jnArGIRoJ0fyUE7FTEpa5CCgzU/GT32ooz7rPDlGch2f8kTR0EjhZwj335MCBQq7Uq5i09ZvQq
oY8wprMw5S5FmHhpqvv5sXBm5NJqazNl9SvIZe0kym0kQMKk8u6Jqf0EAyygQWB2n44Uj3iPtzB6
YP83whsB84UsJD2PIOWomLO9Dc7sgZ6rypvVU9K+6Cklzqjz0ddep7H9pb+EbhcKF0Woveswi05l
kVXc8mpSv08f+CNSNoiOwJfMNx9KmvRgXOpC7zFSFK8YuPFeNiSqwoRe2jIN1xzETDd+AZV+kUae
i6g75mi6sCODABkfE6LG/75fEPgUH54uifAVqJ2fNA7Dr9PSVtHfffxaLRbBt+1OUH40Se74FeLW
552tEIqphqujurRxb8iBMKkXRyPmikty0WA+e2l1csV/9ZQPfzghY2/cf9muqaCktzSZkkorlCxL
VCQaE6DfOnAsfAeZnYCglPjjDGw7wjD1DchBfxbuQy1ZcKt0Mv+WbC44x+Fd1vE6S0hdlXp02zNR
QWn2/0qljR1zDfi9vkZV5AMAdwGzBSXV4wxekQeiOvpY8rolaX/V+oYs+SXLiM+AwzDBA/igor47
fqpZJ7NeuQWX3DCJJ8y29KJEhqWFwy62XU9nmptj1xiWjcNIMzTFS7ld+OCr+bo8RmUZ4cceFsum
ebrCbXF31+fI1kh8Ike1DXQpqlw8cnlZN6N2yuukjGPR8duw1X3rrYjI2vc/0t9yy+/M4vMpDwYf
AtkYqkkCJ8ciHI98KoWv5D9LQQnB7CQnTjG2Qs7YeK8EuAgAbyYRoYvIQZuf5OKSP7hJGSQ+2X8T
0CWRqQzl2jnUJF4s3TkPiKp4EvW2RLFWfZWgnF/yTzrDHwb3DFrh4Zx9l/S8giW5Xhxno0Yzoemm
kpiV+Zj+PtSkLHSpHMD+Uy+7E4jcNfYIOJpCKzeOm0wepIoPmjM2CojYtUL4BevqRXBV44kBMZIs
3OoNkiaa069PMdptUPTGffacQ7T7JFGAUyd6jGDP/+TJ0w5lXdDDh2tE0o9NDlomQbBEEGKwoR87
s0u/tKuldyYJMtV3L5ftlLLGrtZfoQGdDTpbTOGxzdp9hy0P1sKTmvJIKePs8GhgdruPfFBLBFLP
2BXv24NZsROWS+NKhSKWznVcOko0OkMsMj53n+BRp1CdEL+xcqQVaypZpVbz66fMmWM0aep8aFuM
84uvXqu5YGboJ4IYmVWLxOrcri4dzjm8XoOKj5Amu1EWpNAhsXB80KI1wDQ6e2CrYRZeL7iwMY2s
BbEEcsisA1cFdrAHfylKG1A49g7xceTghEXuz5MfbCCSrb48I/eCQo2MPYWkitbusGnkmnt3Av3+
KYr6JU+/DcKTYbZmFS1jzKM+bxAUoyyyUPaVmu0C++m6wMzIpGlSPb5UD5mxYtIun13P3LbqRqdz
OiGovDygOlMODlCZQAmN+Pj16J2rPo5sj04deBtQgg1VJKJ+7iYNL9MHdkruw36lsBkURJkTmOKn
uAs/A0BUd9Okrp9OhzD/veZePVY0qtQhRvil28jyJSTvlW+EjoLkskzUYfRasDjldOhBk9ofL+Lh
/YRO1PghWHwmuaCTXx0HvNih0ihBSM2c8vBX4hva5HmCTAPMsZKEAVMJIo9886zL1Y271+f9FDQ9
7U5muTaojcEgGvj19c3aVWowT6Q1Q4A2reu90ht+VT1tL0A8IIEB6RUsno8Tind21XV2zkEfyWz3
EH4qebh+pmNgqpUTO3fmHZcpncfeYgfTkqaokP+uQRJboKUYv3Il9fxkh/OxuAdQQABuKcCuTYrF
kLDUdTi7+cwgiVMPUItISkaM0WZ3sm/gaIOODIN6o9VXdssEQp+2u6clOLkFPTw2Tb4zqLt/bhtr
pRpOUrqqnhgUYI1ocokUupJnwB4UxtziuS8KqOMAFaMqc2987HyUcXKYPvYJdsU1bRGJBI0c1X6W
qh63nVNsRLCyqDlC1w2RujYce5DxGxDFmR6rxtwXWm2ecqEjnLbF49yxa0ZjaZ0i6wJ6uShs8A7n
P1PMyW/Ts1PfHNpLhL/qzU8TudrR/8B6NVacTXSEu8yy9CLF1XXUTz/cz5rK5pWS3OWNolgTGiKI
nKKSq/m7DHxKmhr/gTxYfulRXzHmfhm4TqoxeWPzQA/3bNi1Dovx0MlChSmxeTx81jWcdcUwlJq+
8YWBbztjJfZXFO+rhxUSwcmnPJD6YQhlniHllO7s7ORgjgQN+SIvzfIuhFKY49KRCd1cg+NfE8gZ
5aRDHQSkqi5+u9IwSxO8E7v0vOidfSfX2EgEGCzxhjBGPGgh3XC8lyOm1bMXNFFmx4lBLhOj/tCL
OCTqAoSpMSekIEbgWdiyTtFH7esDh/dDUWyn8/UIy4ynjJsUereItPuUbq2OmumVtRQnbMDXFeF6
O0q0DJUJmI28znGDwr7PoSCTtsLvwNLEmCRdH72x+KuN9e/sEmFS78/tf9W558nZOBvnZUO4dMs4
ryl44HO4BfRa5EbUXcTiQEAGvrvqzmTyzgJpRAHUo2kctio2QzgT4dZ1o4mUG2mAQq/nV6IxBUW3
bTnqa9GFthnaEjlQCe2epd2PtOGc6bkeMXHI7/XZ+L7wSX8iA6Y0RL0gWKAYL43eU+pADwNnvf9o
lAS42bF0vmMslfosL/hfINImIT7qca6h3THwF8Ni8Egd3X4W/B98E7yOKGBPlpsFd+7S97dN60TN
+/y7rMUMCcic6L36RF2ImlIpnrMXRM6qX4QIwkVWfrro808pMFL6ITpY3iUONwtbsVveUWkWDZ3/
51ttt+CjwSaCdOeZp6yPfNtCwbzWYwZLbHp5gWl66c3mjogS9Dc4sjcOOBuIMA9OOSQ0DX+NmJgH
IDYqVaNK11sWtFqBzO9Y3MpC+LaoFsAZEMwC/WcOcsLToZKlfjmylAMbgoQs8WxdBBlNCTRCHOLb
/uX518JdihRi9YOsXY0qqzzyZrErZtzymMnWKLTYVCfO85FvrbtZxuqNkuBDKPVXOniq0ck2mHaN
NNIfGnSmELbRd+XGezfV/mEgmA7grFEOo4OI60YJVqxeqirNTf6F5Gs6KToP+49TDiqtFzK2BwW1
K+SQ/6n4hFIuU9KbnpuZzULkSKg+AxCBNMqoNTD3MYRl5DHB5xUn/WIm2ufUFox5nxfWXdjeAQVZ
CxJXyzSrB8FOlfXIkc48oUwmhe7OE+hwjGcBBZ6dWE+GrCfKHCYHsVpqX/iEyicly2VMF2J7gXAF
qbSDiaH3YchHdLLu8JNVB4bcfOzJu1JEzrQUp76kH1I+FZpNB27yOyXuSOm3hvS4Rpf/lVXLLN8r
3sOEO5BWohPNfeWjnCAUyEojNTYZ3ZQ6owCGSPVBYqpQmFtuJ2e2zHp1vUsTGMnrlr8s5i+c3AiK
n7+DBUjNPNjHYvxTR42k330BSPUh7uU2tzB7fu5z+oT43H4mQqfPtziYMbzeVnvcFPidNAGqXQiF
DXWVzt+CH3XIaAcTgj+owrL+jxTbTo7Lj5NZKUh7ARsCnffm7NOq1VvkXhyJJylc0tCSAw/g1UGj
Ia+04+Jou6IZreVxLbCL/Qd+lHIi0kI8bfAUtIO/yHnlnr0RkfcHsTSEklWrKfFFfIU0s79K5qKU
mYurwIS/4G2xZQunmKpjHGYaF7H80yrxf/A/Jlp5NDFnBsPKs2uV5e+fcd6f2sww8h2uOUQqJhL1
8BaCAEOctpbSCznmkjuF5oqWvy6DSZnyq4JTqPkzQjddGV0MlmqlGpLWjhUl/Fhnhzrv4oo1r4BQ
40Kqykn4euaROtr19lke6iJsyZY5X3WOfAtZZlxfeVlAS2ExGonRYNDr1Cb/zQQhP3tvF96Zsh5e
fWGU5GGsg0kIth8hCHwkEtxmVJu/MkIcL1NA+uL3C3vHW9C+QgOoUFK+W8WhoOX26A4knJGc6G9D
dOjJQMs4O2/wdybi9WI4Ng6y/gM+BPdonl/urjajWmSA2vY536bZrp18/lCzfV7qp9oNno7tnzLL
aqpb3/Q8lrCkX4LU3l8b8cM+YpUfQm0cwRzVPhb3BSuZ4j7Vbo3CAIeu6Mu6GqFmR6+dAJLDmhBi
mpUbPjKf/0uEa0kccN3QDQtuis1/0aqLo5Kbdzw/3oEnt8++w+Y64WUsQot0Ot2dGBumE835iwPd
vRSa1PEZwqrzczdRjQXwSLEI1ZwA9dCh694HxK/x+uZFHrhfa0y6/oBwotGS6sIYkSRMXgF6YSJP
6N5rrw2m4rivp0mSYAUz04UNhCgc631HWadsDJA+dwf/j9+ilS8dsnnP3gizsZ4F+cdzVJn6gKkp
Z5waUWieXf7/hylxR3GG1AsvDQz/ro4zlU32C/PwrRVymogzEpjTXKK5Fbi2BkEttvwN0XAB0OUD
Ky1K7mh7xSHy2jEFUHmfw76o/1fFmD6wPxcsLmW5KDo84hDNpDhSj2yWluvGHOJ5lP47F5IXOGqv
5LyT9AuE/Mjkd7i3eDmFBHM/6VcbwL8D9b7d8lwgpSZwM8l5Psm/oRnvYpnbPHGfyF2UeqNkcPJ7
26n3y1IdafX81Y1fG+csSa2IbPmBqRVPuu5JqqDgLWuOCF00g36Fe+GS7A4jjhmVMHJpOAgU3lMO
96wW0zbAiKI6eVZohu2jGhU94X3/2PsZxAPK7vmy9mn0jwQKQdOKh6p0jIaJV2KD2KvqipFvdeYY
nUmL5ZHVlTe6RzCIDuMRsQ9yg2dNiPZyK1u1dEyw/wJWQhJXymres7yVUJxaUcLvMLY/xNDLJIQj
k8QEMN+ZRbaCQc7VloxrEVxjz3yYUlfTYUPtYXcIpCypxsCExKe3nmgmDLcjv/R7jKqy4beVTxPR
o7ocOhZrOsuwwER10BHT1IpLo3txIJvXhc4nH8jTfrwkksSbRb09OD/2wO8n/fb59N9pAnaMZMaq
7JVZLJRCX1Rn7NY+k4f1cQLj4AmZtAfNupW2DL/t0do81/2iTsoPJeYmHHMqqwSqK5NCp/rJ8gfG
1sYk6VBaXTL6K5/fo2nZTjgq31bQKlQCgfv4u7BkL5sqVrL+gRIxt5311lzd0tXybk2/DjjZrCtA
5O4XS3aA21CJIXqKd6kejZZZ6Dv4VJmM9qZ5me1IgjZSwaMAm7jZdM408TVyF8QIzoenTglGPdfS
bcE8zdBSXPVLZJr7iF4MXgDmDU5e7GOX11qbnfLDg/qhMs1UkBLPQymwCVtZ1kF8BKdF5HJ12rNI
6ivscw8fokIHZVGjTBCoc0x+liHjq9GDRICdi7j+FyAiG37/+P49nLL2UWZNqL3KlKLvmZLc2qde
L1j0Sr/23FV7rfTAgpXWySmzJuudoASBiCTysxdNewFuQGfBwfDPOvodvmlxedLVDLKMenz0Ov05
bZUwRQAtOr2yiEOXxNnKiONfEoLDI4MSmLpqNc+0Tj6UBC9dnG11i2a+sbhX3wN1pEtOmq2qvgV3
UieSoGHqe47KiziTy/hsX3UHs0PnWrBi0NRsNDFwSq6ynFPcT9y3qS7lfawW1tZO0bxnFrk80Lqc
me3+S62UN6EwScYnq0GR6rYoAlF4AapFEj6XZ7RhgeBskb30HAaZhMvyNv79uMLkRCbObs7Q4GOf
v8xEjyAH/2JyiXKJS+EG+4VKqaggTT+Nil8qsj9+FA3Z/YFln4gRJ6Zs26DMzptdjurR3j2V02vR
9A5nbBCce/QJTg8cCVCbCaRWZzj27mIV1rfZ/lZg0hKfQ585q+zmMGFHvTkBgUpivnnczKzmUCTC
EAniAwzsf9nBxHFqouFc5o+P3qRg+m06MgMjdPv34+jbaA1ZjKdNBWNsaQAttkqzaIlVDvLgxkGL
NfKFQ0RAjDwbxe5tqjDJs4gqkegaHeePxCxLi9wyLqsYycUBrfdmsN95RHL+UUPvcSJ8zteaCn7d
ydbW0jvDGdFK2vt9NSt3PrmmUgnh0hI2nk8xdVFZRRlb6EiXDsjCq3nNR6LZF55sK/+cGX2X4/BL
ZMZZqTxdGkC7jIK0iERYuEy8cYmfgLREc3o8lXj6jKDYUdBeYQhOjgNHzSDdy8AzHulEEfU8dDc4
AjmiCoCkbjvqjj7RGgOmFe4njHOM8Y/3XtmZlmGA95NQw+usRs4Ryif6bMf/GmaMOj6heQ4UjpQe
/6/ry6SGo8w9c/dL38VgJ45NOQ58UMb9x1qiaR/wtltDSFcW5GylRJlv8XARYrzTvkyn7/bDo7s0
eOvdKU/j24MAqgQtgL2yXZnFqj1xw+XQIEwuZmsl14LSFVDCIm+ICogBRsBbLsFab7Kc2FFCekBU
6cVgaP2tksejcYlxgTm7bwHsWIpahGXqaUD/blorD/Be6h5SqEZoCRrG0Cg7qM8o1mllVUMh4VHT
O2xTwYms87I1SGgvo0qWWBFkdaaz0Ke4uLz0aTfY3P56s76zZ+glsh7Fuc/KGPzhZk2oAQjh20wd
6ezjqgz+HQqnaHeklGAHDkk4lFUFffFC83YaK1rvs2XAYrWc2k7gllvXqWkcW9F3tWItKnQNUJZG
t4MdRK/3XgOm2rNni/6mCw3bTxdc/SSo7/FHJZlpkst+80vaYUwo+k8cwPrTN5sB9UnsYve3nNwp
Bq0UGGL0jEYAIdZ7HTmbj084YcQddUpfeCL5uX5HVlx72hjUi0XaChVPOH/ppasIhUgI8k/67BEs
l0BFQwRecLUz0+eLnzM6NS4hpMDAn290NCZugp+cV8Zml3hVWEefFTpXx+xcfCFg9TXgOuPILLS1
5JlNzU3zV89fRIjcLxPmNIoa3Zl4fTBdKIbhnlb81VPQoDfwovSAjVjQtCJphEtI/wWqKg+DO9dS
B5cglKi6t0+191wQxW7jEmMp7o0cZmWP8BqTNqsJcWTsmlhJBVQeNfNlP9LZTrcYcI2BzwuwkjUh
f7DID+IdjU/qQWmHW+4Ku7y4uyaz0YdH2AtD5+XkO66N143wsT+B0ljWTMnHdX67ZeayT8BtdbgT
w7r27m5js6NgaJDcflGxXMCNdbMjklQZVhfSU+8wbCbRCmjHJ1w1HQx4fiN/GdJsm8OBCLSMgHwZ
H6PULaBJO1KUG/Rsks5EPk+BsSnUInf6aHVW7ReP/2NpNKfWqPCn0NoGAnGlb0KCooZVDdrV/A3T
vSo4XEbSM6BEtuVu+mhKbrDk8ffcM+cNE1yi+/lk7KHIDI67BBfISFzTroGjvDkYNXBTyRTHpWun
THe+LalLnLjspGwC7sbpvVMGn10xgIkl7u+L4/HhaLfYFSBL2IW9K8X0iiiJOhL3ZxYKP0JuFks3
+Aq9fdNtwEYKkAcft9BsKfiCqhsmYpb4QHQz3+EertRU5ZsC7/OuU81cMZ/jtDBSI0Dz0dd8TcD/
Zul0hpwoyZKPtD01lqlOA/lReS0jg0zKmh1wExumIV3y77Q2aDpPNJtLEy88TqV1E2hHP5TNStib
pC6fC+G50MtyR+AVmUWOgU4Hw+3e4POWlrvedkQlae6udzCxS3mv9zf7R+BnJrQ3ve20ZpsZG3ZI
6y75Qte0v6cBRpy+iqo9WDIKGch1ND3ujInwjz3/XlYY92W3aEsYZpvM3WH8UI6mzZ4+wsmbXWav
68HXUcor56Un6w==
`protect end_protected
