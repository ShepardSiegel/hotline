`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
I9oj4uT8JgCSXq7nW6SPXllL9U28vzGr3qJeGedJHtNIBDfD7wp5xe4WvKGcnzAR+NeexQIxEMFo
XT/xn7eAiw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WIWZmY2QtI67jm50OGy2VP9355T95KO6QsGFFAA7YUz2f6+4qivHd5OjAtC63oJKt9GxRdJ31Qg5
nJCglbykcMgZYtV8nGESIu3KTbqLDk1irn5zXJLFnp+Q73fhysdGLwzyQNqkv7jYu3E1HuPCxQTJ
1lwCsglUu7suqoXzklg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RTg4ALjUw2vYxYx7cBbEEihK8jE+W+INSv6UC+vZNPa60nQLGIwxJ/4HMmRDcWKdIVPjUoc2Pp1Y
+luqvhYE2W+3vc13HGWuiesmdNVBmkiHay8JUsZlRR1s9GDVtI1p//V1aBTcg6gKOo9h4pR4oUmN
Vn7LuBBbV2r7yLCEv/R4wluYoZMNhSTnUVIcVipNtDd96y+G7yWt2c0LVzzssPkET7Nyu1HBpSGn
nwGIFpkUeUIX/PRTNeh6/m/jZkL3jHdYO6At804D20BiIMnHa3/53Ax0kmQeFqLsTIygzBO7kKmb
HoUClt+wI8wjKLLXmgKUoTcpFzW2hfYNLva8eQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DcjM8snalm/bzzjyBsEEL0i9qSKijRKlmd4uAHDByrDa9pKfoLa1CLXMcJZ4nGQ/V9MHXqkRDWHN
yfOWeCv2us0uYyo0rXp+Uhw6c/U6sxH/IYLq05O1A9JAbOQryLgwQUn8Z5wp1RvpmvIjF6kfIBKo
UpF7z0ZVwnWK/naFEJ4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P1BriXwyD0OlvYADfd721Lffo07QTi0eSBJWJ3TkA5KK4etSPop6aILZmH3s9jzWoUOsyn1VuO+n
TuHjzXfkYdsIuyOY2yE95w5gmmYY0NhoAk8KR3XcGRDHelImO2Uk5sArFzxhmlSigFXm5K9JPj6N
46l3lJe6x4QSVu0IR97h6NsU5TytSlsvBq5XJf8JVophN31EyeMUBNryYCKKhutAPX/hoq+Pr89s
PwK+vQ/WhM7phhxfcjDApVWT7X+NWHWfT2a0AAF2pky6AD4dEnPlJM15S3tXCBFb4FamQrqxeC/h
I8gskKiJ9O5LGkit07zhZpZY+XRpgm71Nh0uiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13296)
`protect data_block
VQg6y32pmzKSXm01BUY+4dk0Nage88ggws2ptU4qrasNRBEymIh4AMmYDG+zTuAd5m8UnkUB1Gw5
s6QQMlV4DbsqQnYiz8AWY/Y1n6J8DAmc7+wscqiUNaiDvpvo5Wc80XIvosjiTRNjt+LaVy0rcoKR
K5VYmSnvtsiG/usAlGDzu0KiP5nmVEAnSEU2VFTWaC/S2y8vmT8aYWgiE0NUNk/T4d/67S6PrjeN
AVv4nZddwcFgIkRsF5h3kE2eWZb4aRNgtKQHxTNTnjVCbtfQ+ZlKYEUnuC3RS84u73ZDJthvkmiW
BgAFv4YYXVlOoFAu4Z8zuxFE612Mnig7TVbiRBMoG678Jy6NTPV9tkS6Ig1NcbAR+EsMrOsdSNWU
fYQO9/iJxy2FvD21PV1n9lyMjRp+3lKWtT3QI0AAyV2YwCoi1xOIBqakS86Cpv4OMX0ohbGb/Co6
H/R69xeMhC4UkKf9LPcpCkUcWM/i57IP35vMnn9RmtHIr6HKjU0VmVZJ7C+gNbZ7T0QIcA2UeNz0
pp83ZUpBuKKeOj3N6UtQn734BIonOehDdQCz4vfW1N6wzjAmYTkysIPjP670/36o0AQ11/rcS1LY
PjCCadr9btfhStdNDLS9nPyaMGAplVrLBqr4Jm/AUTfMBZNmurqgjINq5uLsnhWDvEu42s14UMRy
DtJ+MWO/I2LcKa5lCFTElHCMg69K3mUA4FNAVSehFW7xm5Ins6DDAzOHndHPaiArfUtIJYV6GdaM
LbKwNdCxJG1F08d9Yq1bClOuYL+A7TVescea/7QPw2o+e5Cxm7L+SDr2SNFgKHRJzSTEKkD1NEoe
RhKRQpaKTrdVElygJIGIYEpnVxOg4OBrlOAHILndM/OX96Hb5RDvzdUO+zAD9gJtXq9d3dIgAQyI
iYl8XbefZwjzGS+Hsx1Zj6CsUUxQIZLv7pg8kw/G6Vm0BBLTRv0cAbKOBpkkDrQyvfj7KhZ1Xuhm
YDZdPTTcl09/vI5uwIzAyYO2KJ2fDGKJ6u/gOt5rc4Dqby6g4YREuc/tj3gniv9EJNH7PTZylONh
wDMaMw5ungk5JWSHaAt2rgvncjqt82taF9Jthk2Yc7EBdP7Wz2il6xJo0o66Acv2XEqjukGv2CNo
6xOueF6vvjxsHUexycp4FhygAvcoBeVpGtHs3EbsSbw1IQ8N3qBHjjqbc4fjTWONYM1uX0aKzjhp
DMQ3+LxyfuST05poQNuDTAX4exFpP9zCTe78eSQB9XV/VYu3fAkL+OYcAWvsx9A8y3cz6LuCwlEG
qycRiYrmbAy66zNVEHRHmzUltrbQ7Ldc3vGK2K07R3IafzTbNVAMWW8LJ6dZeILRLw/P6fwSzthO
i2jec6etQJY5Sbnt/OvgeVk0om70eB6HbVjgX6C4s3DeKaDiEf4EfZ0uql5KhjKVCDGlDZ0xy9Nf
QQiiAE4Du5X10kBBiycKkueiv24wro++3G9b8U09ZQFPewmJW22gk7/Hh023hC66vZ+Lx3izMryB
OdweljzQJDKH+a/kNImm5Q50C3JzcKvNw19L2BzTx0lEDQ0iGpDW2kMYLkZmUXMrZfONim5Coh+f
hWpuh7rLECkEfj3jTYAdkPP1cKgItEN014as1lH3RSzjNyAHZFt5FrWdswOXRSMK07wa6GxIawto
fb7bKaXXGi2K8bGGPUywZW9T1cj2BBC27elFX47OYdQTzvVs3tbcjYjpejz8i/DTO5aEhor1yzCd
EtKkSjQ/TGyZmY6xBLM2pURR8KQMu5wtgzwh9DcIRLGec83+5lX3DfBgYdp63WC8t7Vq1AOXsu24
XJt8EAcDDYArDgOZ1P/4sGCj8nN+v7KWzZr99bphqGimfsTCidYejiuCDTi3dcvgj+EYSkEL/zjJ
UAHBeo4K8Omc0cmubmH+2WHPkZ3N+6+kDpYXr6jlZPU0PRrCWfGuabn4K4R/Ix5aq0um5GtzJB9e
OY0/7Jsvnj3+ghtjt4+pfsArlCm2DrJqAhAaV0zYCb+833WFd29Gyh/TrLPGgSihO9tgm6GGBsW9
ad9nq3xUz4okWctTHN2rIrOi0R6S4LDodicY3Y9nPPXs8xJ0Qtef0H3VqwBC/1vZ5lrzvGO4+5wQ
jJiAXEDj2mJfbCt+fAXnATdXLVpc8jn9DPIT35j7tWAx2sLo8UACG8TT8C9Ws8/DHJJzaOFXDcyM
NSHJlH9xzssHU76gGRTYwgl82tYgDQO6Fip5C5D2NDmJg060xcK3ul611jk+4WO9K/sogZ9D8w/+
PKMvTnrYoat1u/651kbrKuZbhArNetUBOQkSL8H44jw2acbCgS+mxkzfpw9Yzckv0LJ9mOROyxHy
+ac3GWwt72K2xNrF+XoFiEttespb9d2ijgKd1x+CgKHEooAuchbkFooxmNYFWoa5KIdGgroPeoru
4ilYEcLT2EN4wJfdmRMPklyhKmrkNgIaeXsU/Z1QguyTwd4s5925jhdoM89ObJ6qsZURnOJ6zTrK
3jz63E84/GeP2vnW3wngbVJv4yzaesLaxjnz5TaRztIg4jIPV9XWcMf/X/nGK32yiTIaOkm9ETCc
hauHyV2hCnHmzGYVH8eAAxITcYQr2L0DA5WH0zGdr+X43Jq7s2W5JeuMo08yU6rBY34/Dluz+XQS
5W026Wo2h+ePBkB7loGzQG0IdTawrj3eifBhy4gCClgXM7z4prxNg6vep9gsf926EGIPZVqtFHgv
khU75ZK441AjYRQvZKAYg2gbsHwK0teWn8bp8KEVKQI3FD0GeIPjGtkhVfFIagUGNAjzNS+PawzS
D1osV4OD6JdHxErWQnFC6mUdCB/SBz/HxkFQ9KtJwaxYIj+RylFLM1vTHH1PdBjOCtOmLMSQnELI
pIOmrTZg8FAioInx75SRipF6nVJeyC3++rNLr7w8nZuIOeaWOU7Gyi37IZ3RcKN6bykf8Y5KdTqf
Vcx9tsxDX6ZCPWNW45vwRojLj+Rr4JbGXT/zSe/vv8Cf3GIH2ktiPnfcqscghlXOu3C5ljRVo6od
o9gztiwnXRAhxXVvOgKG7ap2DSln/xa5A36DIjDj7dP1+VOxJNHSg8NtnVaqrx1DU93O9h5s3nxh
5c4EXXN0Jg9kbfuQNDaaI62eeRrISzKnWcCfhshTQ6E+JtiEVWU3U87h6rI5Am5YyOA1tbp1sBks
p7hILWdiHDrs9kmEy9R8I/DDuzZ1uVXOTuS/s3ANwicFTqiAZwic0dDu6IMQVTbXWPvYq763J1Ak
4i/DpyxyNEcPvhYHOWa5mJuMdMLo8O4uG4y4eBNLmGkXLEY/p4jkJP0Cu7IRv4NBa6R2NXPFsfuq
a5LuMCmP2pR027jdQFvNDI5cre3DTAhH2Bc/4JkFLyNMKzqv0uk76IteeF+5LAJYzRf6VAdgwmGE
wPw76Rf+Q0eUgWjZPbozj1F7QqsbuzDEC0cXgWN7goft+Rruk4mkn0J+BU5rdI73MW0aUGAvGF9I
3GbB18fG8WHWQGCzgn0VSqfSp9M/T7lQODLixlam05KW9DueD9U9AJDtcbtk5sn5l6HxPHEWoN71
1Qu9PtQZUIAqDcuqUrTnkDB7fAaUbzv/458vzQJVMNA1QVrjazwd2K9XtgSKtzzLA2T+Agq0D091
pHZn6tFRN0LuRktlgxDsXIvgOSeb/SJ+OUHnvOKB8wyzoFMrklXD+034Z4h/sEZd6LcpwBtuuYWD
0n744MmPwwQ3fpIXwAsqYkVRCY3VnQPQ5VxLvlqxwL86dwurZiobHKRWh3Ojca+B3oI5q7iOvdDY
n4xOEFkgq98PTl/PjAnDFgps//5Rtv+QTjPoTs0U2YmBs9LXoE4MQWJFOOBjbmrNZuVTqHl6HEoQ
eSoI5QRgqV8rK4Z5iTY9PWrfR8tY6w+0o5BsxVfZ3RfX4OWL8Wn9VAZlJrf6lnDTdAJ8vR4f+2OJ
Ncuaf+vjvM1CZir7NUfTT/okn8etzpKE7Tq5Z9f9dpyXCs40ggbxJishsKNvE7o1dWspegf0xMqM
CJx1EaCRjZvIsm7DpjHdZ2nbth50FHVJ4bZK/ESeQ7GFsM5U6UZn1lpYbDkJM38Fx8IHTLN1BVZn
0kY/+2fE9ODsiynwLpJcbN2dkS9EEGsqAN/3w/VTS4J/DN8T7vo5xNTBYt6Ssg5jivKik8ZA7pib
uKNhtDwSRrZjanO2Cee9Q5EtRcALLkncU2vuJZ2yr6xA7ep9+gvwCwEPp3ZWldz5Hwk0jBEqLptS
MKEATQGi5OuRhR2micE1txVRJJlEii/rSC5dIDVtUtQ2J1jwKQ5+cWGAgchclfjqe3Dn08dARsWR
OjG8WYJnpwjh8daMyd/tXOvwTF6c2Wgzm/KQkeQRBpvMZS99RjJ3Wzh09RUZ2QkksrdL02/whOJh
xsf02OHBwe7lB5Xtz5AlXiz91plzc9XClagxXSUlDVko3GQlwQGBoH4j5/ujSytU2WRCIOrGhofN
UDochriF2Z9IKqXtLKotS491nIN7sqE9bnK1vbhVs6fLBKqutHXyEb/Wb3/fLWPhk+Z2tJcvwYUF
NbR7y8/onYmTnXgby+vBldLT1mtw7EdAFYnKDeYzxxZcR740D1p13vQWBfhnNm8oDGklsnJUsbPm
d3yxpfIa7xQCCl8NYc17OKMZzjfYBe4fTLGfIK91kZBgMtndvWLZeRAp9O+qTRIoneG1U0V22AWg
PQ+lsmOAkqaKX6Mii+fuS+i/YvqLi8c2NlRQ0P+j9FpELGhm3Q1crKNgZ6iPG9UmFW7lnKsZsSlx
lHQllRRFd/2ToCRf+S9ICfY7Ukbn8+8JXZESF0v9VYa1eQi75WUfgD+VjaWaV+naxqYC6kTpYWe3
Vkdz8FlHfZR8R7QzMCh6Xo5JCZ91jCF2H6eZTrxocIpvc7pnIMIIlB9LI1T0ZepWw393Sk5P7tP4
+ANl3WjmujB1kjiyk5D9t0LXDFXwPLwjZeZtWyXEGvF69K3+FdpOvqVv/HP2rRAIKPhi2LxZq5vf
V4LXnJc9Vpd+bzAsF0XIBtGRkDwS3OoK0NedPhtS+lvPsD1clqbzCAllEH/lecMRYxGi27gCKS/6
4kXiuPrXiu2Uu2akVk9aJ/ZsNujVU3nTjgjoBIcso7XErlXLdWF5GsymN5PMF10RuJ/M+sveQgD3
4mx4CoZR+P7ysOV7R3G9iwRILe95MwsNQlS4Si5lDp0OorSQRJREmOQliD0eWXjYdkd5qNbg0cmD
06qgTA1VxVuFZUH5zWe4605EV9L78ZOzk4LGgh5+fhPXTdF3CE1VuwXxeb0LvNUW6ZcIoJr6bqPA
inPjTDWTO6B5iVeIRCK/xI0j6NHOgJDAObNBTytTxEJNCM6oNahMsThJVQDxIZrmCvceTzmCud3b
J1QpPfsbiH0fWyKaasqvHN/oJmFgx9BYz4kEOCS+C1vjyNL4EeRKWmmq1mHfxjlxJglk0lPI2Sn2
n/YLRBHQ5zbGlocfXv9hsBx2DaYiatF7PehL2g6iQ/gQt5feZ7n0vZSobJZzhrHRv5IPMlWD30Kw
IcuMSWbi2AvCVLoiw/a3LEfmgMz/UyAYVh4s9klXgsdg5GaM3dym/OtGBsP/SN/aN9T6iq2boAHJ
y9KnCBFFN8DAENyOmEU9ghH8UYX4va5Qv8nX8aa27hrDijh9nDGJb0Q/hmuo1Z4zFOaKiWMjXBCu
EDqdRytDxlBd9BkN9WXQfdG2Qqs8f2a7gkGUuelEHwKEfNx3uE06K811KxfWvFpELkRIKb2JrZ6b
lTnwoR7t+205KQBTMgnD0piTxtu2tb3v0XMRJnNgK/qxgcT21GqAyDG4eGmo4d2zltmwgIMALL3s
KCQGitK17c5SsrQd5JSUYmjvwZkD2papA3FeHUV4ub+klH+1n4lpHIsOND7eXP0BnoncWxqp/GuC
0wyjsdTZxWWngUaEr4Tacq4PMZ7YDbsDRAUDZc8leP11nBE+L/NIHqknfG3ia0CXedgykSJagwu9
KpMFtk3hJvH29TlpK1ufBCO5KjKg8ikMZPQyApF6p31NBaywuIKRja1066r58TzSn25XhcVs8x8D
4xI6mPyR2aJ7FOcuskiCFz/2bNv6j52sc0G9jaaIbgEANs2PNvxTi4wIA0+s9w0rU2yqILYvHo4g
G1FYTWkPf/lR2DnuGjeGuv+US6CY0kz17tts+FdN/fvIm556McF11EFVEz/OfUd6sH3hFG6QldQV
LUcUvIWDKOvFcF9iVvgvcCmuEzQ5kt3OCCW7sNWIcMj1CjnITSDL4Ayr6bmG83+akfeALUmcawVU
QEPRXGqy2hq8NSBbF2e6+yssN8brun4JLInhc/hG2yeesmZgTH+Hb5Cjgb0sgyT6JHBeI3wJfvOp
9LyMRQTYmOZF64kXNrbI0+Up0MhgCX+GLfeGJuu6lqPYShXyOoOG+R5qXwuZgxY6me9iLCGzm0I8
4jfYQIW9WOIJaPY4L4rCL5DIahbpVuOEr+2UJ2Q1Mt2PSSehMWKRrMmPhEZMYGrpuy2eTqs89FQH
yHmAFi7yp+6DsbUL4qq/V4MPwGRv5iJt7kF3YOGvprHH5cMRTSjGyWLtUt6qPZ7riwADcnnuuDb1
2vqG1/Uw/+lQROm2k5SPa5sFU70bGhqa270BJkTylT39OMe9V6FIGSfisd5BZh72iTAKCad0Gxxt
uKVsCqJ2XYGaY2EWIeVU8I4jaWQtJBKk4W0bahJwgk0AP/TE1Or9467fI761P1U4H2wNDpz7N9oR
E2mFRyyOzL64Y9uz3WFZom/eBuHiiB5dZAar3oZVYkEQ1yX+1bMXiEtcBzRRrWmZVw9SU1UAvQx9
OtLKddSc85/47M2s/vW4T85ITnnZXgbROx9+TveOJfspN0slyfGrfSvOLddofdl4VLyjthaAnQjr
996/KPccn3h/9OECXE4z5NkeEdoo8zHviAdlsd7Si2E9S2A0kcgbgCi0GZO61pv2nO2Vh1aqz9ms
fWBw2r0CLhF93wwEvxTmFhPeJynUtzaZpI3TBFQPRWkhYcuQCRGQbQ1fm5hRkXHWBINhSJAbZnCh
dTRHqogOG4+4N/nTQFJ00RtBJyQfAbGKiSfQDxD0YSPxgcIcPOvNeqSs+Y4CzS8W5KP/Kf/s7oto
sF6EXf648Xcjk/aWyIes70rI1/gs+fRielgo1FR2uPMeLdSU6d2ZMvN8Vdv8TXpqUBZmLB/q0kwP
8UKR2Vs0BaUCPkWBQTjwobmQ5xumX1Q7r4SU2eXIX+jQZMzJsWxdlDQ9X4q77WudGPxosLqlDse7
QTJxgrxh+un7K8lVKB7W1UXsLuDndzpS/X0e5EENbcibfA2f0OWABxpPFz5oUJdf8CyZEVL71o4y
fBDxPhgCi4C1EBPJ/ASDel2xeAQwjA1fXBvaJZVgrsHU0crTKcBdZL12+xm/y9OTVl+n69aDDDK6
ht8Z+A1MlnHK5EAH9fwfkQc+YVxTRP96dtya/QXPG7AuuWFjQOcbZat/kWuQmvqqfXV1C0mpcvBD
FpFCg2PoEuZp8Xw4k0Beq83Jl0f30X3UeHxsU7Z65DQyUV+eqJaoemCsxFuGqZHioxt5Ja90Kq0K
6IGqbErPspvW2K0NAqdtZ9/kNgWWq+Knvn1hCdud6Z76XludAxsacIkA4MRSLvqpjgjNZy3eGbAp
AeXFs5Jm97Q98cNtwgu1alX0hXnuv5Vc66RGkUxka5379SoaEzrkGZvx5dhlY6WqpjeDbQJX19H1
UuCy1+YD/Qo5mdkTsagyYyX2fZgBa9uVP0zpHyxTwOYPnUjpa+1EA3i77LS6ZS4/+MNpkIPITbpE
Vb4/w4lVsnxkfO3g4g6dCtMR5b0J8cW2G9bgE37TuYI4PN0B84dDFqTMgrR4RryhxaOYY+WCxmTn
nD6shh0qnjREyZAY4tOsnoNPmvr9Py2RY7gWE6I8wAl9nhFbhqnEpe2L1ZO9gIc5Ay4W2E5T1ElK
Bb6XsSVdFoKRgPtyUnXa8Xt2b/h+wUnvM1gULFW0j/XlR1bEKYmDf7itjVaPOOvyol1+qWy2NzaC
f6/yRM+wofqFRJnZmkRp1x8k92UQyLiRL3xTnHwXio6YFE6h1rTwBQR/NwMQLPlmTXOfSD2jSt4e
dRJywoayieCQewepDbMvtPs0PXtjrLwIIRPvD4EyYcYDdrSbmSz/4I5+ARxVbYrcDpJq05Sja0CQ
pe3O9ibnXvokK5ksrkn6apC7sGYLFb5TM36fuOA7SNCvIf1x6p5UQTX4+Edd9zkXceArqCrfo++y
Bs4aQn49lc/P+NHMJtWdxDgxUIfl4BcNC4lG1OyvUT3XMdsHOT+C6CSu2An8Rdp6O6HbSrhc9CDt
eTm6JynBP9ov6JUVVeDXZZlE6RuE3ARuo6Y9KW2vaz2g9ToLOlmx1G597KuPK4m5YXkzzCAcQNsG
IBF8nEGRuJ84DnhJYMM+KYyNHeer22o0BlsHYP2Yn/Rv55WiOK0JieHwglAoBYsYFJ35vXvUTmSG
RRcS1i1yw+pB6ipDDgjznGk9hLBordjS/7/8VNy4C+nmLmQVe2DDpV3reI44VbMMeHe3bDc72p9l
HuZ5i03/8zCYN6s+fZBUsCpfAAYwfe4nOkVh3Wc2NXWNS72mc9AgJIVFEXXB70sXHbTMmGsv5T99
H/kfc1kNpgofIi67lY3etTpE8pqTiY6vl7mr7x/xaQKn0eGAzC9POnFbotyeYpMiB6DNtDaFDdxd
4y07cak5BV4kg42mop4O6cm76EInsD+LgfTrfQp6yKkVWBtDXMpySJj4qc6OVINPvXBQtSO7GIuD
tx6YG30LLpSRB1Bj+3WnJJ0/No2tML7psNpr/XoN1Gkzb4zzHMu7W1qV6LZwEWPP22zSY07UaUYi
xy/8C0KZGFsA0AASl1DMoEzZTBXe5d2oea3jgxPZ04vUCKkz7AuXQOxZ3Q3N5lte9UNVzXHQy7pt
2DVOkw+C0log0OajKBTuA8VI/Fg8DJ4TgbtuWXR0VQEKES0T1nTCUMeZ2oQ++LANdQ1h/gxF9+6m
S137L2BTRFjA7csVl5OXeQc9KXHGqf3u+tzXUIHDLIUyqdjhomSxBknWqIfE8w6YtJ3acuyTNSIL
8Tu5X2vEEqQWeQt5pzVxpsmJWaZAoaNnFyYY+umov7SjIU7tV/Bh0fqbC0i2KXbQSVqoZVY/qQxC
JNneUsatNziv465HHRDiZP7x9PKlMmRqTU9ahAVN+af2SagiruAsLLMjcWch8V9PdQh6nsPjlD/B
qHnQ65PMbd7Kj2xqP7DP1DY+lXs6MbIkAelpYYzqAq0yRZKlmvTgK6FHCvunH8umfXu2B3yeEICy
4dFguu6eDBOOfIk/BEg9VovFO4TuWHGN63HCWOeclR+ZiCOYuMxr8ieMlIIyx9x8zIJ/67LreD1X
bZp/84Dw4keVS9TUpyapwyDibjaoLFHQdiUS2RIaFigsLc+WfP+KB5FOct133qHRQDqVGkrI/rVV
3JWnZexSSsUMzg88mnkBdaUeRpxcHZzK2XDw0svvEqYj2j7CvVe2TPI42wemxGjhGMkvrIrCEzwP
zAJBSGCtBhqItXBWKUmvuT7laOkHvdyL7SpNgYu/KKm/22hGhq9kC7v3B+rIHGrMnN7zYJP6eyOA
vZXY3yv6nbnPI9oBNaujGkG20Eejqk52B21TtKWvoZSTzFF2XK7UJueMMKBO3VmbEY7HG3Hk8kNL
x3Yy1qiO21R8E2qN+wlv5sjCn4MuFOnyy6Qh5rhaURGMd4c+7DpVXzk4O6JEQIE/g5XP4Hb/By7d
2hxHqpKPVDb+pDhbVvKaEsk9VkV4JnSTBHdSeKn7R6q31ImSdc+Ogsp5E9xriFEhgqUglK2rsCNW
WNDNbh9XkXUjnWbL37NM1UlwxkbD9I7mi1e5AePPRKPnyvYbdKebMk9vEQxzmIg2O2DRJXLH/Wpd
mpq5ZBTm6LoK9zDl7vsNoh+5NTLYhklo7/6TBlnfM5LtwUl7xBntr5tmWKVFgmDblsIg47z2PZqK
Bt9bTc7niHBQZ15SwRXTzw0QLNqvbu/pxO+ib0tyRjURier7ENNxrz1HkLkgEXbws2BKXuuzWThw
/tcB5qFfH1w1OVINtTBr+ccakDkI1XHOQ4dvwFae2FCIJLRGbu7QkNHbGB1OzEXc+C0MLIY2bhLT
ittn+Z8XXqQasCPXWSNsCcgVwHmfm1iHRVCZyzZ8JJRrSgb60ST4MvshbuNNBVNWVtOSKFR2sseY
s7D4gcz/fxc9dV/LG8LoGoY46oFmv3YDBP7g88RS/fX4NOsiLw0DMaahuACUzB6O5egTzQhvJByi
4sjsfh3NjHhVjSq0tAYbz0BAKdxo+L4ynj3OHDZthfL3IO+vbeiCSKaHqn86zLQ3ImnVjK6QMBjf
03fhXLAex9b+2mMR36NXclHx4iKi4mo5EQTZy+n1k95ochLu45/dqgXroLJ9L8EegQ1VFF4GFHn3
/fvlHFzVde6pnxr0axaJKguExcHNAeEMeXYqcXIRrpiR8sSantbMv5+dMPLpNCsfIsGh9lIVkJ9j
H/7AdFRgoqjtqcrW98ejkrP+eHCc7Guy7il9HBnC0P7O0W6FvqFIUw1sl/454291sjuwufpaLVOd
qHDYnV1RhCj1NwBmo7r9SVw5pNRyH0+tbiMaMntFwfHWRi12jPtoi871rGHPLww4QJ43CfkLap6G
dgX87Z+J3y8hWGZXDnSP2fK75OCoLdNukRgvo3TeO4Gt3DtymOMR8BfsXU6DYU/ijxv2k9ssCoP/
oCcSshmPbCP23L/GZxjmj9TFLucDHocJ5F/KaDpJzW8NwIz+EKG0lUivcJt6HdZ6W+2To5/lI3Ft
DDlJBMpBP/d7zUQJhr9BhKjGezqyW4v9Cjb2BSxI+g+ysHbwAgm7Id6dDAQz/K4EOykwl4erFmBs
4tB3AKregZzbkUcE0bqP6fwluUCgEO10NaIP/14V9AbViGsAQCzRn0lyRxGbzGImr3IHOln5M+uS
S8wNAJbsNER5RBQhOHoCkTAJhB8yKP5VohGEY0jVHOl8SwsDKzgHshoITYfQVMXrJccNLOmVbq5D
gr/k6ClR6rM1vbGBNUb0ezeqg6+1vF0KJHfgmerfXEFIk5q+4jSr+hYq1k5UntWzGyZ5yJ0hgSHn
benFkmBonThahxSCUq5qlnDicJipAlZc07Plts5pI/ttZxHKQ1ksxkNS64F20WmRJLP88TeicAzA
FiTkO+awe+sSgqgZsIR0llicHqF3dK2ITL3O+NNPZOXt2P0acZQtrzf4vDh8AKGpgqeugE0Jcny0
KmnALIT39xaXyZAbDihn6QPD0H7/neliSFFwDDQgeNKjoQbZwA5HxEt/CfFJ+xmZMeX0s7kf9l7b
KLEiiVyoug2CI/i5neHzAIw7Klkbi7K80pQEiMJ46W7z6VJZ5VG8UiL/ITW/f+p16TPFxp/zUmzL
i+lG/gV2AmhEVEHVtnN+hYMUbXf2fjlB2P3ZoeEqvrtbKGL3AQhF9ONgvb3/Cc6wpV4GSmDYsCcM
ovGwSCatWDvohOp5gCq71FFv1UqnPdri4p0qMLQOyw/q6kJW6xiBSMlqtBd0OZFnzeZ8geshsSP9
aHgDUmTp7yGBlu6hjO9hFdmKnj0KkWfgyXH2pwGNjcy/Mi809b8Yg5N/OZXKsKQScYDj3hsrNja6
Fa7aZ61iH1KTRVnd0WNCBI9tZWU1zTXI17me7lrkHUqyj8dszqx4uA75JaxSMn+JNhe/2MTBl1IO
OuvxMMkC4ucmdYsuoQauTUH560pz2sNRbgsXzjzV6SHFus/m43US2pY/NtvMFMpSYENqAhY+0aSb
XVORmDqujvZu/x0OsqCe1C/JpZRdqcVqAf7XmyBCKkPdscRXnBe1q5FQD8whi3Z8ltfIfZQYeqP4
wNDIBMA8FBQvD/BgWXPa8vsOktfEG2IydIRktzOXmoHikR3WRwlh1XYUZqHC3GfnzcN3nFL8hSu/
xpHsCPp04bPKkI7b+W5xZ1g50BZp8kaKFX/+t8vQpTvoNTOkWcwgOy96r00fTkzi/+Emjl1JGYcF
ynSU2VYUg3FItEGCG23F9oXejg1wJm6/PkKGinwteWZ0TsahGbl15S3bKsn+Khu23WyOAq47/Pky
kmi0cgnOVtlsSkU0Jh8Op0z64QE+1HxLBIJ+cCaNlTFmO3te5hEm3yvL1cLUXi93KFOBENBiTLhZ
Ej4pFgSa1zVMG2E2vde9d9zI/UgfeeqtDjSUYDnsw5UxEeS0c4uXzmfyt0/CtpKfiOhF0CtgSFO9
lF8fux0csVcuI4Cae44/gFerAGxYgAJjeqRdYAVmGX6GtQFjAmucN+t/40EgcJfm0ZqFMMKrrt2M
MZQtW4miTrLbJb1zw+YpWibhmukQtku4vTynRviqwnsrge2xFXhXZQ5S5Dh+ggq+U1SoLs4HLc+g
Axqp26P/rTQPhSmOR8mGrxUNeVNLqw0K98ewNEYilCM3OfYIEuq22NYIRixQfEbtN8xLjpqbX9Zv
6esaAbGQHMrJEQFHfntF7kVIDjP5eRLXzfpDhI0+0S9cOia1+xwI8E+2uBjfGMfBKGT+hj47TtgP
8AOEAd3zPu/OwnmoVS6RpZ5nUgZCiOgPek1pBWmBDz9eCt//SFroi6Na4FgGoep1O/5BzQSdRPyZ
+DDwi6ijnzBlTD7ys9CWWT4ys5e5GDgvKssn7xLH65Ks0I7EXwnya6R/zrMqthjsKGBwLvDJKL5W
+koC5PdA4pmzvwSHyyzHFFx23xu9STOBfivwpVir92P6OWnRK1ITL5GRnEBYcDa5yOPZ9icD9aam
Gurt4c9BNflZhk6v+1F3hGdRdtImpA1tdAe8cVPIQ4LVXU/yiWps25xoYneUMuIZ31mGBz8WslKe
Rn1+dqTXD5GXuzT+KEydEyoamxxXrwQeJa3cUQmynGsBC7AWZQJK361CdOQmEosi2/S1KzcVK/wL
DusdqdWpq1gl/qhdNRO/Znyi6D0Coe0gT7zH0loGjz9G/+kJuGQF642z6CqFO7COl2ZfmhFgPiiq
a+9XFnUNvPk2+yKiZVKbZiemjtqyruTzvFbAw9JzY9UGiej5TWwb2IQ3p8Y+Pyp5RKxsec1TI++p
SMEYaS/uSA4jdC0ZCFsCS3jefCLHFl8EYGYKWD0FO9pc1PSTeNDK1T1LWwapbnD6tOcH1USqRy6m
c/xDN/5IZzSlH0CGaRtL6Jh52pfijVcXfOWNaCHG6AoNxfmZVBYvBajYsawzYUC9OcJvtaY+5xqs
rAyuY8LeVhJBiZxwaWQGOyvzjcN+3X3a5NGOyqlabiU+ivVWdyk0YFv4SHaR3nTLTadIWhFK0SOH
Pdf8UHzf1kDWJImG++2yMSyWGN1EwUWtA0QA9Whx5AOTpCwVOLcS9DMHcdW+KVtYYojRP8i25vjI
Pc1MVbsb0C8yf4L7exh4gAH2kn7PwGmzRHJrPvyD8SxLcW/iH+W3Z6lQIMNlRFtsUw9TswR9607r
EGseLzrmMR42ZVPV0poq/XnTDC0LZsAYXOQrgMFcEhISP1hi3kLE6MoqqvdpDNibEExZAmJuIN9X
MWAuPS0jnJT6K6T5tqF1yqxDc1Z/2vFSfNFZSWT+U/14obVdBPnHYYIXO8ap0mkbC/kQo5j7cq0N
Gu5ke689FgSOWsptMhxzjgWty5hQjH/1YtA7KEWm/04DcxlUsG2IBOuqoQgsabYQbuMdk9LOD7qO
I6rtPDBq/D9pmnDli90Zm55DyUbCfwPMZftmmUia1fUOapj1DKC1QnLwSuGFd/5MkI1WlZuw06mT
sAVdQ7sfyY7qzIhMPBew4ZN6emww3C7yTDiOXhn3cN8OHQoaPyd8hDELNiqT/bvc17Ijif3nfDYU
PdbpqWtNOIi6CDykNPYEwH8u5xq4I2z4ZvBx0K9AJgie8zPpr+jzTmw7yZPBNIzPgVpCoKid7S2M
TOshV1Zw/NX7lPkqdzA034t8qcrbLdFVIcg5wI2Hiuj7tD8dxHJOnyVXRZO5CAU7mi2++aQowf5d
KRbOfii3wgBKJdQZe6DNWdoIIIsahXsrLMWBbd9Kv0IiL4JJECY8XjhmFL0T+TM79i4BaGxpEa9a
BRxZ95RrwgCn3rdQdakdSxT0wMfli1magVc+J+zpOWk3k+p+QOvktiNcVh7+RH1fJEhpF8gzID7Y
ifZJcE60f99mNo2g1Z2i6BYXQDWSSwc8PH0/Ru6pHwhxjGojg+VYdTsPCf50xSkO6A+82A9j+xAu
wr1db9FfmdgHwePDlDX0B/JNIC7hEUzYIcV1DwNCKun6wtBJ7a/6bmhdmbQgI5T7VlR7WU57S2E7
AcTMu8I7+trPfxIwqXFqlcePXGnFbWYfRpl/QMFKy0VKS37NTUXbaOd01kWD8WKosdMh9ztRa0KA
Q3oejtyjid/qwMaTAjPH0RYQ36R3y9+zoqFDezoOKYM18GDaMU3z5M9ZFRJFi9wNRiqeVHGrcvng
wAftBacjbP0f+W+onc5ODL4P+bkBBuw83VUks4hkfgBqWxeCWI9cR0p8CdeJHxCHajPeM5h6NGXu
jQU4jOMNlJIjz/k0dVGs5hgP+k2qPhItqAXtdriH9aZHo9kbjTY4oGeMaAitFvBy0bFshj6DsZZ9
0EK2nFTiLa9Wbu8+CA9E6oEJkK2GaoMMKYMbhxxIj95ucFsnvs5wxctAk7NS0yDeglbsjO1yMcgk
cEi7POXTD2xcAZjTzQbtU0jchZqoMx86hcq6Fc6Rw7q8EGIo9/RbSEaogO6EGHX/qjM47RHtDstz
YFh+HKbKoMv5HHMh/flImRjTLv8nkTzICLBl7GhxROj7Ne0fCppqv792SHaEt4lyzz3GCueQJ1nr
aJ74jjsgI3TkSh+wNPeoIdOgvJ/x5qDhcEcdu0VMT8A4s7JPxtD629sPbhd+wx16I0KeikYmRTEJ
PUDebL+XtRcrrDFXbSAqA3GGaDIGkP9UpPlj7Q55giUu4RSQwVIWuAJTz+mhwNnfrYUVo+fwTBHE
ojkkBJShYOYIqsyGApv++frKi1UDne5g7ERBqayX6WcwSpFW6rX86FXhXSECHnkNUA+Qg9pEsjrB
Ybv8SgmRi1MGyC4REr0W7JMkIzdoyQs3FZdSb/nYxvJXFUlIlAea1EnzuW79P4i8yIXhn1CNgjNN
kjH+Zvg65C+n2w/GaBc/qm0WrWtnENFNSye1f7fEEhwYY8tYh3TDLygiBhtVOZTQp7t8SC/AnRUB
hQO/CUv9FMEBkYGncmD9d3jm89RT7VDt53uPxrpSQKpCkq/3cHPI8AyjNCPlG0BIoTJDxsJLM9Uc
yx0nh/z7XL60f26tgpy30kS2vBKJXDxkVjodWN9OR8dFXQfPzC/DtXiX/437Gy7tPSG9oVbfmsEd
clRTAadFUJOuvSlXAtQnePAfgTq4Z907zijJEO2jkmh6u8xMWi7CX5CPniaik6wgfXOZWsjfdY97
zRGJTNufbpVwk8i5Z0GxxvuhKB8OSAB5CQKPSqQEDs6GwXPnBZW21LVOX3tdELHX5IW+I4dXZ1uJ
kjV4gSR2fIfeJlNnM55/bXIHCAi7jxCkt1yjbGxgtaR1jBm25kB/vRtaid5DO9oUOyZGe+ksGGiM
cOL0lYqVrVRDCSNUHySEzhqnI3Xq8b+Nupx3tKWKPwbCYQzQamLltsTRiJXP0TsJmG8UaePqBsUt
PtN7nc93cNgI4ZIKRYkUdT42tKtS2aMAZf83QOBwKtjKeZ4bxSgZFbcuvR4YE4Rjh6hC8U3jzmYH
/2wqZN72it9oGeOgARVnaUyv/0AowtZacj4Z5h02A+JjaW8YyJSuuLVv9af6I0attBbPG6zpc7md
KqQKbukMTdqR+HsbfivN82lHfLcmwIQNL3GAjjHWwq3rEnTYPRarlNVKCuE37pVH0snxqQ4GBsFJ
T9wvve2+oSbmth4ogVGbkWU8P7rafLCcukyqMUKv3yhTyUfXbWcwldwcXHQxEuifuyiBrkvp4Fjv
kcVxBTVgb3XEQjV+UVV/hp1BjhlSU/oHBFhso1tBUiuNnq2zr6NW9Th2eeoe5Y9FZ6nr+OxELAtI
LLbFGY+D9oJ9SfeiFF4I5e5SpBCPPAyYPTwybOPxBodCwZD1k2vvs4rchDEFSISf9Gq/ntKgn7gV
L3Qnx5V6KDP5W2x+KyPHCEyB/V/GaZ5FUW6qP7T2tX8kgqiPAUdorEBYPv2Rn6Ty60XT0J698rq/
/k8v5cbaEIdNzKcsHMJEdBqtjFjtVLIhJ653jHM178dH3bp2Wtorn6Ut3x3kEqSZaVD3nx3PIVBF
hYW/7v5dvTekcky2nX99w2ItXeoUIZJ/J0qjO1a+mjlwWtP35tIkdpqVr8KjU0i30tXBqrn+PqmQ
tGxwl5XUGCM4gNLQrAt6MH7C6168n2uz04ghhdiy90cg3dwFtWD4wVWV9RaFRltbTM8mCOYOfIKN
A2HArOcq2NBa/fNNFUUnClEqTC4kdZT9NHFwiowMfoIH8qi8BMiiM3DDeqQ/EtSIjcfccAOko+fb
Q+HVQyMbubSYDieXsg0z6evdppxDQQQdxtqvkuYubt1XhgN7BdOqtErfWFdI9jlxvPKdEgvRROKA
D2OKPmAf8Kg1wPtEpzxLkYFPFBro0TyL8il+eu63jw2v0Xb2aB3KNpWmwqhSJpQ/ATJ+TVC+DC5n
ntqX2Ccx9Ei1nA9t8mTWpr1zJQJX42DGupvmbyjhvnUVA6ShiJQaXeBsSVzU0+ILN2pG73DeAXD7
t5jj0F0bpZM0xIKBmQAkRSQNU49stXsjmRhPDkaNzXuZLhhOtMRteASkD7XHSGIDFr7u+1oNEHy8
mZkwllXf0unyW5h8t2q04nZUGdifORl6n68kC9oUY5w4QyEaTRYvbDGIrTytnkLlmsuaf5Qugwsg
tmaTySc3qng50GwjvB80PBVrz0O1rKZNyTCdfBFG/Hid8LjpnHjFoI7QAIaBMwOcNOFHemKXqX5S
f4dXdaYOiXhvd5AY829HubORXtfjKn+dagi+sx+OZne96Km7g/ZOJnvjqWFtgO89NfZxdyfaSVkd
YlO4cPvlkG1RNChVDCDLVpwwWV2SJbpXmjz5+CcAhLsX1oVjRAZX4mxh1ruCyS8nS4poLqfFfqhM
aK2cFQshtUzyUn/hh7TXDDg4oi9gnOnoyGSyP4DlAu6nCnJOBEXgk/gI3m4MwDpITA3b5iNNzryr
P0ynrKBxlGh3hiQzTvHKtBG8Qkdzh1y9QZdetjS4cskKRFtI89EqLQBtfUwi3zA9V1e8HLZSEVFs
QEGzTMbTxAHki4/XZ83R6VCvppaE7c4WGUS55xDefSTMyzi4t1Eqk0N7NPq6itBCBDKBjsDs+p4f
ieflkZjH4fzDPBPTEsGLvrsn9vWKiInb6Jx8RwMg1SkNhIe/oBXtVFvGmg4bPbjpJhlVT6/APZQ3
z5fNK/UNvECsF50gNE50xq69TXRudU7/CYQzs3IOLjLQ53TbFs5d0SfjLQ8/677SKTeUH5jSpNLj
A4v01udDv0Jr150jdUco1iiGfRKUM86gZanPNl9WR/4rakemHMSv+pIz94EyyHRNSycLINZz1sXO
gG8mzqQz4XTOVceEqdXIEHt2gx12UoXQ6VVZRKdE+XkBg0D1VtGcYxiBMapaKH+Sw7rYeFxI9aMZ
hel5Vedk+zVUbPJJ+6ls
`protect end_protected
