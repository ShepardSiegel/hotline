`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NmnhK+y/hJIlU5n3kv+qXds8eGDZ/aEYuYHDJr9XXmuSnCIXGjst8dewOkIPemd5GARpIVrTOLJ5
PfLMaN5eJA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ERnSok5BNvNf8m/lmB7iobgg/c5M3/EjvlzkMjXni0WEMZWMauzCFE29M9fkC9AFW6p7H6GU2Arf
Covq3FSP9JiTPGWmjq2A+iv9q51DeY+l97r3OhkoTgUaApshwLSuUfX1LCsZ5d6Q4+xEyN9R3NMY
hQRrBMPqbr/NmrpN2fA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
p15u81s9hx/I/IKCI1Y1ahjOyIaP2bIj37FcKuVtXIuLc7UE/Hn9FTj8VfJHC7pXm/WFpMHYpMAh
VRzFIl4z+ECJGkyqGR+kpQghXpE+C8M/WuFwGoK3WNlZ0NuTsMiT6sYaY/Z7N8bKY7hY0zy+snj8
U4sfy/KEXmINyaSwYbtKHN9jSv0GMZb2mtP6g41u6TLO5sojy8QurMtOHOKfoLOQNN9AIlbFTbMy
VCythvh0NmFviT7lysD5AKnYLXS4a9OXUvWal2ig90QCbeBvG5Py+TWBJlDzMZbK7w9rO3qgnEL6
8kuQWHLlNNHcky2Owvt926Ic1o8bep2+ofxyWg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
37ryxVRsOaRlxX5Ia/YXYI3UIyoeY8I6A/OqDua/MNI6g0XItW/BuLDRKWJbR5SkLtNm1blkC3gd
L1XONu439WGKGY4B+1bEQCDRBT3jGaduJOy7QO4p0+ytsIgUMfFv/0LyDOfDeCg7xYKgj4xwkR2r
QHriIHG/0pPYF3pu3Rw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BY9we6vxALjK6Z7b08NNLHzDYtwS20b6yltVQXhkexV7zTJVZSdAB5M5rfz923LLOBEWSQfXYuEM
Xtz18zalJTQxA+zy2uYWoi4dP2TcQAV+7eE3y1d6O7uYR0kpxm1y+DeiDwEPSweHspGFf6Rt3c4f
9hSzKRCx50lehJSceC0u2c2wmEmOMPhkLq5uNczrrMabcyUDouTIeQ7z1DhMfw35HB+zAr+g2hX7
DIdj4HY//m8TttshfKQ2Ux4jzNidQk13foZr5p/XOyDyzfV8iHNIhVL1sx/k/UF4nBxcs69zAq5I
2rcjftRxaMA1rcQOHJ8bMV/dwJxeonrvi2lOSQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30912)
`protect data_block
v2MnwiTPcvpRvxGFlCE9fkvfG9AkSZTOWhjYw1g8uwyLXImq3TezY0xtyLKMwBnbRMbCBQgq8NB9
8uWRMME6DjWFZa3BuIOczLDVGOlfbz/r7qlb4F1N0j55VkOnD/GAJX4pUaGTAwoPf05Px3BcfD9V
SrXSGQxQ9whkEYdizyrpyv9skktZZwg73UJmdxLCn481kh2YEaJF711wIvwzqmQP6u+dLF1Oa9Vv
fedd8La1B3fVbFI+MYllLHmKqCzFFXWcqpEpN9rM1yIlD+GkUGcuZzXnIODrYxViGJclqF6/vGj+
7u4pO8qBD9/obmmNeMJIY1h0rvLhWtKKqhOHb14190n6rKl7AN2ViqclybBTtTsO3YoppXPcbIQu
MlmXkVp1k9h5XaQvivo2ZJSYpTDoMfGc86theoyY9vDImeY+62iq1OCOPN2VDZ/jOalFu4+G1OdK
FQCmwYD7arwrLGUQmJqVnWbo/T4S9BHXEDlfMbA1fENoo9WerCsRWmhJLazHh5CebpvDDoESRvAB
lU+x8/u9yChfWaczFkHApUWLjcBZYk3f/GUSyiyB1HuXlVLLUrOHUel+d2lY/qO71vS+UaW3Zwrz
ER10D6rdXVPBzRPHVGX+4JYdZn9JnjgPNMRal6D0bDefrzFjqV2Sf4Xzfkd9to3Tw6FjKAqU63lR
RboaCnIGRmOmgGagxu1I2sni8Q2R2po6ExkDws2Ux+ON23bJePfnMsLGFYZ0M1M2ZbX61be3mbpG
UL8HlaQSrBj3Ig6dduCFx4opcYc5L3i5VU/Hx1wpLIgpmLrXplzlo1Ro61QBh/EdFllVj2X7K8CP
SL36xk1tbVfsViTf9wirI3i7z71VKSxEkfOEE3UBN94WeD+v6vO6yUbnZ+qbIFLOTGWMZ843xxMx
ildUcUrHbPpLxcc5uwzc/EQ7e9xS93u43cxLIFUIZmKSQtvMBTyrP3AnP8eJ3cbhE0MGlvLpZla5
K25MDg2amNx7yb5x5OYdB5qpqUkxGgapEFg+y4dAfoi+V9yrjz3YXmJrA02Nok6gaGHZmw9vwLWM
Eev2b1t4zfQ+53obDG2h0MQGjHmC3jGB/Y2Pw1+Om+R+5IComtdD3MBF8Mw7uArcbqovIQfCBFhS
luAgjY3pSJ9UmkMvGhZ+ZXTMwpJDmSS769fZsD/i5uSpScJuwgna4rw1fCNqnr9lQcJLvSV9ULJq
7Q9RqVzV/5sj3nmSk8OVVvyTrZceKzKj9XRupUNEK+c5gkNTtAQXNkuJoaY5IRG1wvX2s+FkYxEO
rDpeH8tGCDIcihW0ZNoXlkPLfXN2lm9uhqFuQX05qm6hdcdLXgTLIBM5cMWCednB9BlWkFVvnfRD
UMbG+USpgi4ROAvEGGvYgDdK3LHWq07LKrM4qiRvOl98fOrO5YshnMgAK3BI46jKvAtKQkQmVrAV
6U4WgReRmCjEbx4+IV55p3z65PZpqfxKxjfg0xHx+sElXUj90MNHHBRFHHzwtWFJ86Y73vAJPeaw
e2/goN4MasNX1ECExQT/jX7op1kYuW3+9jh1gxcNNK9n6MpCaaGLPbDqXisaLq9qihWdrcaAZ/nt
Wif5V7JPMlx+BJONGXUFWkyobM0INdEgsG+1WoMVfrrUgLbHGes1JmBAhUSB+gE59fYauoiHfGX+
FPfih2PAUmSWArE3gUulA2TPxWlSLISDAdV4gQlwZj2sqiFo9+D3zKqysNigdYJd2ku/cIL72y41
8bJcn3tmzYbyd8eYvCpkJu7VQTkOdcn8M8hVQlx4yBWuITgIaxvo9W6qc+FAQOavI5LTHG9ds/0c
L+NGZ3T0JvNbIt8OdW+vOaclABDu+wdPEflzzTDAiXXCi3XpWVrXTy73IoSAa5wM+127JN1jh6mx
q/+9tRRudyA2g938BkHuMpXJ8D8BOb97tMQoXlXi6IcU7ikRmunR2ofxfiorQSUWPIpPkdkyQYuA
W+aIYLbXuwV76Y3T7H6TmNpI6BD/I39RCERSDPwONcF4hxlmNwJuO3/iU9wYz9zUV8LVHQ29wNpw
uCLdu7+tpXxASZwO9srbp5Mw9+cSd+mUo5Fp0QR8ROb5KYNcXyTRl5VUBqKBdgJ3WwNNdU0mq+nY
caprWwaOsUplx2FXzg0M9k7knBvgoVkcTS0fNkJk9jb6vXJzCSyzmayvF3tiuhLEm4Q0RqObOP34
23hpdyOjNoJLfchUUBXor4EFrdkvi3PPI04Q37IDuLPleW/i4msWpT1/DoCbRVewgoM4/bSzym74
g9FVLn/4DF2yT63PTQJXb5Mnd3YjQQRerwzoVd/1oAgjqSNsVPNmT+DAo1ZvNJtDRN1TvJffw+iK
mDiGUS8uy/oW6qOoeP0pJFKmpqPkbrA1PRuRWDOU8C+wxtA9cR61+Qf3MKgGNHvkTOrbDfeb8dmb
cYsnloXSsd4hwiSxOYtweLHVgb7lmQSl6fKXPLrnmB08tCg/pm+s/Z5W9OZUz7SMmqHpM+H6YFLY
BWIAXnnFe/+Hhs6FGcbmDqelI6kt6iwjQJbcEiYEjMSOSu8/H8+R7YJbev+LVpsdELoo70OVFV00
y9tFcQLpGP0HuhcRpZ7xEAbJUR1bnrNjr5YNYSLSTJoIijoSDj96CoZuhfQsewRKSUXVdEBEcanG
kLuFMX7+DHlpmfDzfWYa8x99DJOsrURyI2hWjSOSVfMpoAuKAoBPjVUutmmemoU4Op/LVlTfG5ON
5ZEo+7AM+eh4P8v9i2L9KFGOEx/pGx5YjlfAS5AbRkSKmcp2+kqDLbtQ9RwLfBII3j9Ju7r0P2/g
vcdsVVGLnDV9sR25VbNlAhVukolPbLFJQPGVWMmq05uLHPVMrtY+Xfm6nCYfv1QJRnryJTAOuARw
0yjaPnrp3dE144LKwlunVlLQvu3eLDMu4fP+5COHnkRbePqWoVEuKIkkGMT+E9UbMm5JVxx4suZP
H1XtwV2Rd5qmcoA3WtnxveWqNYKalR+iwS1Xxdka4gOmKfy64Dwp5UZf8cgshQoMu2flQbC1DJn0
8YhRzchBxTCTHw/hVQQ9ePbLncN9VSAzn4tUr2kt8CJGWYEHkzx/fZkVHacQYGB3fn7oqeYh4PwR
zCGD4C6b2OqwiIF0Imw9nsfAp11I7jo1aotat0u8UWagAYK+/GALCLZrkSraznKMBXzF6m/GNhSz
U3bjFz+Yk9QUmIRmeFiJ4DHEp9mgmNPxZt1IQLE3L6o4trbVO4vlvD/pElO7iEQdcbxhIyA0W9G/
QJoWUhPXGN+AxHRs0bp7oUSWQzvYF7iAzOGg6/BGO6cb/HIIdAcj55/I467LTqZtGMrvnca44Xvq
ykKP0VEhx1j8YGgsucdN6jquhwoRBLeLAGuUw8QXQ9PNdhi2U77vr+3X0sHGn38OP8zo1yTLkC/Y
k9CQQp+/dgBZnMIGKTvYOiQWKJcEsqbtmCsX3gIjTLU1Y8A7rElh6sBCKHcrPPj6cGjaKSHG680n
8Mnm+VKgiWfLMgBAM5NXokqAvGKBavzVfvhiikSKs5UclcAErYJokDNA9psy9LmilDFj5XXw451i
a5zVNRhnmGvJua8nM7NXbFps+VqpcSiE1uM+ITvhIAfdWfcYrR+FdefqeZ1VnvlEpeGnLSMVOvsb
T5cTVPlxbdF5wtDFZyGvwJGT5ZgIrzID6sVMjuJp6KGsASCqdl5CI6BVK1IaSfSnZnRkFzmrc7zX
BQwM2vT7QSAojQ8b0KfWpFX80sifuLVGnafcYIkgk9+mxF2LyJQSO4RdgfT8iY2TofWnT0jgQT7N
JxrgRWsutdiqoKU4pr2fXSwNzdLBktB0m5KQ9VZg9OFii2DZd3m2dfIMlLgMUWK2h9JY0QmlLae6
UDcuox8QJAtqz+9o8Xs1SlSBes9s9JJ8SImswmq+8UuPqtZSkYYFZlL3QD/Um53PhSAI44pNKxaw
KhSud2BRarq3SzrdgwPhpfpEsoGDelajVTs+tW2AIQXVFutkk/tnSyD+ocuoAXodFq3LFZPdQ0P/
P7a3ZsHAyCsd3eba2Ptu52nTiCI9KVSCYc9/22K5NMVmy7bvzakzJv1kciQxyUO0RIa7++e/fbRV
r04gnB2nJZjV3BOmALZZGr+os20nEZi/b8pwET0aRKuAXM/BWZiav52OVUWPu70jUCLi4jV1EUnM
g9mhHEnermZSoeNTo55IKPq2l8jocEiW0PXH4yNBkF0tKtcOEhtqSuGY79y9O+pjlG+ZKSnAx+xa
Lrybp+TjWlZqzlRIhdx6qhvSgQk5Yfd6nUQz3GwsGxdhho3lxfzeUnVWNeKKSc4WPqlbHl3RDX9J
LnOKK1KkBCxCtPToSbyFL2AbLjhyUFPqLwtocyuJijyULD2fr+UwOPYrpkWIwQQWZZAd5XPz1baD
6QbU58+Wzri6RP5IhW2wgR/8JMTEC14aMU6cEMO85UUW4yxDCGTZaKAd0pbb1491OXz8nChkYEw9
BxfMYlpwfSHkN9tVAJddXWqSMIvMAru4am9W5Jrv59+Trjrg4vyw9ba2ReUae+4gwCdHCP85c3Fo
bZrf1HyAwwqviN7RQ1Fu4BbBfhunjGa9UOMkW/e6tItdcWrjzUg/hptZ/4QxKS4wv5ubfkF5ZfVD
EvkY+SbOwV3rdiyzwPorqB9yUMw14NrQFcpu4tYDJVvoYb06HROZY0Bdc7mj2hKAWsQWc8KTiGpQ
yo2H/v9d+jQuzHUuPKK2QOfhT9wEmz3JP8VLS9cIGpn+5o98dsOCl7+He16BTbPc9tPZ9niCLpQg
CeTrLnlOq3gPiONHm8dkLDZ2fsdXBHllmrKTIVQkC47mrjU4APzOM8X26oqww6GYa49hJecmcD1+
bgozMqcy+CvarawVwiIuVVZlLyRa5044AB4McQNeuTaV6mjo3engX/sdHYg4CETsc/AcI4GsNpFW
t/XpXQ0SzNvZ6RvcZCD+rH5T22lG5QLtYOfRnK64YoxVmj/Iq+a534R1ntrI2JvSWZUMZ1Jlfb4I
9A/nAXMt9KdFtj7tNg7IC3q8T/MdNrnD8FSn5bI1gbqleBcn+XFSopWsApia17AagIkZ8FgtsoX3
EJCRekwnX+1NRzfGZGwAPAn3yLPaUV9/VppNUeTDmm741IigiCTCTQg6k/aDMKc5SuQbDGdJGfxk
HjEJw58/KIDsIzRS33Cnq85imRM6UFB3Q7a+dcJuHK7EEdTVK6WtWC8eyIrebxOr8a7toLIO2AjQ
CMjW+c3KGSOhz9CGpSG03HlALGrsq/TyKoZoa57sMUamdt7HzYvCVCHfUc8iicBBFD6L+2ikjk7T
k8xmAwEKZxB1VBISPISn9I8+M1rJcB/FvlM5KQ0P3GfdMNGv+ytUHLrR/AGPI7iN6IUJ8O19NfvS
Kygkv1n1LFoGxDUZkPz9gE1umSbOD3SgCqSrREWJ6xpTwOM7CWeJvGw347NgUMFPzEsIszpS9O+J
tC6THprnd/YbBMjzs2aAG4RKxg23tGW37L4lnYY9Wc123RKt3neKYEuKlINKRoZRvLxBvd94m1Xq
hDPD4lYL7jqiw3PM6FcS4E/US8W8jgZR2nT4krqom5mZgfygrOXuxGUQykJ48l5IN2ReM4tlV6eP
zJwZuzp5Y7AL3GXheJfUhI93hAIGSSqGL/QZSaA8BhBxT0Q4nlHD53kcbhSoO3Zudl7/jc9RXJQW
Yp+sWjR+ltzfD5kx5URODf4SA+zuiBR5X6AnNr0ndqRS4lH7TvPvuRmvQz77+mvYH5HW6KXqkycB
gK9rXqlmiZhcc83GSzn3EduVe0XN5ZhDUXyWj2pvRZXEjXpb8B1DFNeJQZ1ppWhPav5GChb9bXcQ
/BtnUeCKtD9pgTeaqm1Tm/ng2R1r6Qy8AXd8WwchZPSKZTpNQfeDBUF5kUHFjPKgi+GJ6yAf1Arm
ICp9e8wn5uki9+tCIdLg1JSYCbcF9WFjDWKg7VJPq8nRUjg202UsHTqQs8BTBVcE973L4D5BClH7
dzHV2ittyClH+brRqZXrkSb486++P56li3a/++SNeXx/76dqCld7Jc3o09GLxWZo+PrEzmAeVPda
gx8Bh5nEweCSPiG5vvF0bB1lKUK4YZAC2si+wOF/r23jgj03Kq3p+B8OK5vyrCCW4Swh6DwlWg/A
oqb+VnkqcqEhCsR4RiG/zc5WfCmhtdZanadUzXPzy5ZdhegbOz1xYgUvm9HrHKCBog+j5BNH9GKs
C/nOqByKfGtl4L3qLZElUi3ztJOjG7/bdcZx8Er6QqfUoW3pEQyTEw2Or38/zBDO/mjnEY1qQ6Cf
psbZCesK9AxkarAF2PxHKi69fvklGmK2CcJtg6JdGrwJUXc/uM3FwrwMHzfvmXXps6fE9KMMfIUI
q8i9pz1RAN69Vqm7AEjgf4AXwnRSKXfl+ERT3Qp9iWuPrm+F+UvCxnNoEIffsx0YkGrn0Ps2manu
exevqrFbC1Y3pcyRi07rvSxO/dPfkZX2zZpQHlS4y98xuvZ4/2kbXcpibS4mF6kt5F/eEei9/VzE
HFnj32oWLy9MjYZ53UDm23n9TFHUj+SoRTeqftrH1yeNP+sS3f+OH/+xmZTh/0FsDa30m9aQDa/S
6N20P7otUjyjTzshRCPbHiHKxnEvvSBYP+hhRWL4DBHORMl5Va5VgdRAkF5arAb9valCUToCl2y5
yl92vTSuJjou70j3XMWP2Vxq4wBm/VFM5hnpv7m4zFKm5iyB0wSr+FDnAKmdVLlB1N8KfVWwruta
4CxS6aO07mLW4A/TDIgRan54+vHWnFgWcNMR9Cg4csV9SrMUiJvEOjXZWRfOrCfEuccQU8gWoEea
LllsYAOYh4jfF6v8pwl9hc6GkEaUrSr4HhSBbu1EIn6vOO7D/KEQA83ZtUefUzfz1vFGOJz+lcIC
NxN9L6PmlvXFpQrsseSpoFaCjqL7cLklQoCCKPqIl2HN1yAqO3YvOgerbrWFQPx67PxhgXMq+IDK
QB23Fv67TSyWYUQHknxlCC4XohR39v/efcnG0KW1QQieuEuJJP9H7WWvEj08AsApwS6EDlmc5Ir1
plZG4+Y9cm69ynb1Gx7O59fo1cc/8/xwEOi0bA5u+JgBIr9V00Jz9wRYwLLLqgxS/DcC4KbNHeTV
ZoMtTgtD1Ga4GQ7EMnrsbZOG+gHAmXe9/dGUw7cLIFqFp+RlI2RtZqq3HYqzMWPW90eU66QowNxw
9sP4RX4dzebiHLtoUbeDqmlTBs5i92z6DbZmlHDmPxhm0ngpDH9h9ak4xydORGkKWTVdkglvRJXC
9MfFnWiaFfrZyTtG3IdpwefxPBGcNsHu094jBHohJitwa9AGw4PBdCJbV/qgJLVbf4unNvbQcSzB
tQGpnGxL9PoPKw7WfbJHBME2iQ8K+DbRTeW7so3c7j8eZhTTqPNMn6kwKgopb693snS2Gf8tiHhn
ytpp/2bDN7qmV6DQn/UVcBfICyvqC2RkpqGTFsQ0JvjgF1Nx7wrCagn4k11WcU+XcEi0wxgtSJ6F
xY8bCnPxMkyEf2WwM44vXK+6XsXB4eqZw10+2P3RO4Urrq8N1Artts2ZUrDJo9pbZIvu3ENFKqTg
VMs/er2qJf/9k16sUVqQGfC28KRNV+9diUB9BJz3SfD7gTbRunpPb2Zxh3Ie3uW/3GlxWKDA+cBs
INu08S0S02pcSdgjlT1ocpmVS7fIsvCawZM8wX7maHE4DUECmgOetWN/1uMk6EJwHmQcmx+bshGD
QZApbB231pZ9u95xBt/XSEoiaaKQDZUixz4UekxhbK7BL+vAx1Brgsz3Q+YucF840uPb9p5lF4Jp
dP/zFzgmGDr3qSaNvQXlkgd/0xnJLiLBhzZkXaSM7yGZVaLw4+G5l56CZkeC7rBlPODJNo0luRaK
eMZchkP10kRJTjzPbX7CxYqNVgLsGziXXJ4oLXQgVEdnEi0/gW5vE3Do6RMUTClhS7VJk+Xykd6c
Mi5YAv9CPsOkY4xshGwubkG5yJbMUqANcqMrUjhLUtTZ19KBQssnVnrPKu4m4KIPFMB30MroTkH2
+KZ5BPzfvVUx53bImydFIZYTmb6rD4i2gvXc4eAWQLmVYA2kAl50psB16NVFQnSqC1RtA4muCy6H
AOBxjAWKt0+8SWr7PDh/NSFq3+zbFvVQ3k76om2UykLd6g7m6nyAZLRQ7ridQklfnQEXVvJxQPFS
XUhWZubyFXdFRMRmGgYrVSZCjmpUyO0A7sgKwONif4UAY5arB98Au9U5HVBJXKG761xmjrPLy2Rx
TlYedQpwjEph8kyG+57XEgy6uUrhWEl5JXxNHm6GceWi283J4KS0AiXQwCwG9OftTq54nK1aJQ+4
hJOs9n61Ijv+DaWiekEKlVilvagyRckbch5LU/UIIAGQMjjQY2vtRDZ8i9RTqrbUgWT9m0uNzNSe
vzfZDqr4d9NOOXgQ4IFT/C1IBqsBZSM3Si8lMA79wRb2CkT4itwumur5WLFB2Hozv4uJo3/bcuCV
vUNk2ioXid/p92iYWiPG68+v0cw1ypBl+hbijT7GkbBWpM14kFOdubkHkMLiGfPGqoMsRW4Vt139
aq7zXdSxJVO0f4pWtymqECY84nr61HBrkuQ68e5mF1exZU2XHRpxuOrlxH4DkPE7O2J2pt5dp1/1
RPnOBgG9wXYa9AJb19AMgZjwiVkgP/dd3QrbXOb+CVcpRWarJ7rG6ARHnIkMzk9zFtL6ZuuaoB1+
3XZpQVrmbyqcbpekfHr5T4sMJ0lhTYEm1ezINAKYKRqePDoLD2KXv7RxwMPsvaR7g+3tycyGcmMu
MmSscZN6wkw9CRO1GVoeNNrG/TxmCWd+yeKV8D6XA6DdfBnJbc6IA6ta6DBIZtKbIyP5N/9QYPBD
JDD+5WdH8boi83A4ujBTybby3BTZ0Zd7l+PQhnuS/cWNt3nQ8mnjTYtS1J+FAfe1xmdfBpTdsLT9
+F/m02hPvOAG2796wEv7fH7+UGKAqi4+Gt428/inTSdCgzZ8e5BDH8Q6+9e+L3Go7S86BNAQpdfA
wHGel5unmEglljiPdHC10x0SAA02WEU9PeTFx+4QAiXoJInowiyQdZI7Q5nEfeYW5vidcESzeUTG
pDNg1T2W9fl7DsOm77sX1Siac+W0eUVIMaFpt+eUSA8H3AUtQ58T/lFNJb9Dk7ianRpcZuImsjqk
Gw+QauY4r+brydERjVFNUoyFYSl7FxDX6n+7M/2zcMC4qGpMl/TRVISx+TzS4f5Pg49+0ZnoHaZk
ommJe5lo8wLMnT78zEwgwd8G1qVZukGKqSJABmMyyqt1vly+Ff0fFGoWJHLajLt5ojnQNIPS4QQ+
WeScUC6ye/HqXzI+wM0aHeHwXjYdyA/2gaL5zDb2OgmZ+OndDOyfkVujKy17+QC7PJ/kOLBo2xzx
sVMKU/2mh/MEmYhVtU+ZjN62HXBO9vSx93pKJbr1xbSWK1Wy0ITlPY3LG6BDsoO3zKrVSuemwv+F
O6M66GDchSjARMPBco0NGgU/5bO0tepK9qBqBLAoNvj1jW8t5zyUApFI5XmCzKh0ETArryzVe+QH
DUWrzUnYdgacT10G/0UcdeP81sGSF0JzP9ml4iyLE7jIfC9lEXwAXLRt8Bzdl5vFX6rGHUjwO/jq
LgwDKLfOdj1vKCNBbvahAPBJCSey/pKL+rmKlbWChJvUJ47b7bbPGhl1H60bb0ksvnVPr7Tavh/w
LugtrTNkDgSQWha9bzR/EDq2nkFVDQ0wkzLuB97WNq+9iN31amKS/qB8E4wP8ZCYpQVurfGk7Tsp
du6+A4TSm8aOl5tQ0OQNSSeWCUJqXePnO3hJwZcakVpOjHkew6mawtDIackGA50WdrZYTFdnjDFi
eO8NuBDLiXPJAeukTI1/r9qhSjOLpAJlymASfNERmPT6pza92px05P0LddhsRBMPhVSLyZihWAJT
LmxaeqQ1W1vZTLRwQigyLcGGsK3qMV/ZnwuT9Z5CO2rmSSw5qYFtGd2LF8lOP1w3+6zLGpxBLXuP
5BI1dW02PmvcI6L2j8Xb1LGOKUc3a2JbB0tU1H2eUsUn1LfABt6sRVrFC4MWleWaJxpVw8CVml6i
SW4UktF1SeSmln6uOk3gvPM/nKxz6y0kzZPxaZD1FRuFQjy/ZBityNf24x/fIKqNypPVDT80y2HD
d/An7bb+P4qs+1wFuAqGq3LgKJuLEOWoUivc8TpAJwUr3+6XP5mUxvHqxSXcaI/SrX7i/OKt720k
O0lA9IH4cDMVGd8GIFnwM/1SgYgkAkkh7iT2VVTSqUqKSQozOYBsSEPcx6hyZX8g8PGJji/MD3L8
/W0UY5EMd8crZma8tpv+Tysy/hPZ7Ut0THewDzj7BZr2kZqTEqNcOkKHOMPMOOEkyWftf0N+Ej8y
0RD5Sae6Wsn5m6qC9oUETrOVKDDyrVWlIFfDuEP3B0VrC642RwZ8KbnzrRulM6lh/Z/fm+x4du54
yDnOUfmrumaV1DwFGYNe0n4sAb+NQ2XquovVkMi2rc1l6nM87zzpQOKT9dGkV9+iADMSp6tih6JQ
Yl8SNhShmfVeF2ItiuHCY4Q01A7/pSk3Zvm21xaPHjRDMKiXh4xSTX+3qF/bsGfqoIrBa/3xkbBV
3CumyrbZ+jNBRqbiMzRabTb5kCYhp6rt54V0WARDY20+F2Wh9dLq+WySmvrzCiVye4Pp9Fz2SVWR
MvIv2lmACh1l24j8pqXtcpcxyNGr3u+4xrRbYx3djTbXuN+Dmpa8du3ldovF7g/gCk2z9YKzg48l
0NsRXAZMBHPHhudV8a+a2n7MwxBnTPmv/ivi6rKvIeISXFxPLwt7w7AqNMKJTzFvKyRfq3VnpX1j
ncAvk0Xrgul1mDEtFIJU1dbcSJfpxdwQd7iG9AWr6nMQ5Jr608ifVkJWU1XgUHsOcidwjhF65m3P
BsTxSsOcmwIFcA3L44i+i2+NotRnwIyCWl3RK7IRP1xt1TxKPj40HCcrDkngUTJRGr14soWvEmYi
hu06CW6/uIG5p5yblHqqmHWzMjdX79xHGp1Jez1wHqmcl3siQJ8Ax8IZcqpTLZBQSj79PzVjaPKZ
sSR3HlXZoVTH6Nfh4N8IjchYW9ovpkcIxGovnlWy8YR/f/IX9K5rqOSfQPy72j++sK/9FBU4AQuY
e00cpoB7yQ0kBFMBUCCPPq/bKNxze8aTorxd1XwYjujEvJylR/xZi6LuN4C1C7O8rR9g2qXqLpLC
fR6OmLWt4zIdJ83hiY9usCThM68bDS/uquQ2u1//bJjSS+RQa3iXAULN1u2Kg86cth0getFPxzmT
nT2zQKxXNHQWUqo/ORoWEDsZ7/eICFplSRkY7aIFuCl02Q6Yu+lNqpavIiWYw+9uoPgTBCoo7AVc
CcBd4KytUpOk56Mh0qtbpNdgmMORX02UDbYl6FzSOq83SZs0aFUMeAgFyToqimhNHOTGO3FK484N
Kd3KxTvEMKhZeHv27FdRoEPT4G2BL6oxMBoB1zUEytKUEFFrxPA8pJBx/FI9CBzWl/3zIhMjTvyz
CaXW68bQlDetC/FpZ0q/NDDfaSAYmORvT4y698Hd4B26kp2kQ3mTKU+daCUStcN2ipIJaCr6967y
JdAV2Eo33XBYOEuqpLNshoc/p93vcZCCrH7DFKMy2HbGpQMml+Sx1jOv8m1J3KnHzuvDU7y6vCGY
AeRwXpAWYtLJTOtdn/Ux9FDav2M8u6wnKMx4n9FpEUchdI2SjQ+1LREKpuo/RSGMKa1eUHMwMyZb
UM7f9DTi1RbyhFNMatd4zOMqlmREIyGNAjj/rCiX1wNVl5JykMgL/Vf18tty5dG/YsGHgu5Gf4N5
7sV2Poe+xx1+e6TXinV/pXrt5wHtbdGKgo4r+Vh+oMyRLHfpl3hjtivkmq1JOrP6tf2ZPR86XzIO
Iu5FL1c5LoUYm5b8QhVPQyqNEDh6HnXvbLwiJovyHpoR50/Py4WFbLSyyX6+SBEpyZUbS8vwr0UZ
WOeTuSjJY8yosoRiNTGZl7A6+OpHDc4O6fByRrY175Pdtnn/tZ7aWkClQOkrIMbOMj/HUm7K3gyH
X/bJxgt7TNi5LMOdDSClHGrrUVmKjACnUrU/JDGKsI1gZ5qeexQywtYbaktUKlcvQliGAzFj9M7y
5Pt+i+Udu0ENGzNBU4gUfVnteQQuPvgBZ008PyNvT9TKlZry+eoiw5N1kiGq8ud41nAoIDJv1k4i
rKHlVfIge2NLK3/7OJqYI77+ON2y36frTlbiXrPY/ZhghdkroeKfq1nqXZ5ivZMpZ9Q6XDTGaE6u
9QiB9JsA+1e7T2ZZVdcxhaLiqdm1L59EquV+gZi4uCP4CR8qDgHafi0sgLEtkHDMp6bNuViuSCuo
D0wKkQCt5K+/hVgZBpcOzpm3DHHkFRDZnijFXLtV6lVL5H4cD8ttCxjfDqxa7Fbh9mGQGmG3K+/2
TVmZjclxloU40GyqUyxHPlmyXSLw6NQeQO+BN5867tHs72cxvnRlfUOIqDddgO1z+Em7O57xUpg+
1E5vYZe6tH7SsMa0LFJ0QJwg53/P+p+unwCDuQj/YOfWNCLlfx8jaWS279B9EAfwHJ1egSKQntYv
wEi+Qiy0A7ZAG9n/FaOzCb9I7FZDMIgnhz8UmgQpVpTQtJj7OF/YjQMJlryTMzXD4IfQRAYcp7xA
ge4lae7D7gJW42O/G/TblfvJOqfg3ozto+o+gMJA8DZ2SAn1iXlJ/JHS1wBPGQoM6bYHHRj+5Ceb
qwtOTwJMkxbcv6YPgCWDpV0WeZiGjo1SFXROiMBBBzDP26bOi2+cD0a8gpWnMT2Shoi1QTAEwtjQ
4a6tUEGM3YbBZyyYxGBtxM1Mxj9bAeyC9zIUlm/fMBQWlHVrhlOGyuKjXdG7cgaG6A8ubW/UseJd
cWRj4plbxFw1T88C+MT7XSW4MxkavGTKxFnDORzTBNiq1f3++U/4Pa/XJ43hoHVt3ZBQMswNuq1T
01LGNMHARjkM/Eq+nDXt7WvV4XF8QwAnYBbsryLWBYCNSlHidws3z3uSdfZ0w1RglVldPgy04RPs
l6tq5OrzXrhiDkoas+nTb08yIJrc5FVhrD1GTfrDrNO4wasMnKYOVkNBVaQOexoMUkiigLBu8Q1n
xgNHoBKkWU7HWAb+ZzoVlSOKJo1bJOWKl4CVV3UVo9roh/fHhDAYlex5QxMxSxgsRahsUYVRyiCw
9Fo6IHTH7GIyUlUxuFRgMQBC07fTJBC+6bjWXkZzhknwhIXo8RoRkemcjtc8EyMJF1yH1pSLKImU
iymFEAjB0qKIcIYyCbqUo7ltCDXWine3N1BBxAu3BxvPSXg3rRVpObxF4pSNFQfqzndIuq9TPl/L
Jm8dgiWiV0G5qN4e21ZWoFqv+R9bXQn4c/XXNstzmYPLUMyAW1Mw8GKT1XAgXMktAwHaDCpeXbnx
NLDwA71Yp6fJ23ZdhgIHKGYRf4BPJwQUvdYky7bdneU1byvwCEtk+IGO7WnOgT/atDWCm2ELCdAq
m38Omw5TWUhXyHp+KOyfuSKCglbyvt2pr6XZpgeWQwqmUiCwpynX/qiDyuVi5xZEk0N6UBlCVx/x
TU9QeoLmTf4ESlLd32cij5xfG5eD3ddcBrh4Eelnv4aOTG+2e1IhZt6ewi497NeA0n7cbx4wRlKB
yb19evoPKfDYSV2hrYcnsqtQpCgjBiLSjjWzMoieiWUIyHn6X0lcGz+svlQafuWuqFFDel9jBKzQ
0nqUVRhhwwkDWr55k3rs4l7YLpusYn62JoKyYKIhr+WxI4Wed1gP5f8Eq/xHOWIX9SloX+D5dd3e
iaKZansmD+ptNf1fiDwhLCXq2Y/r/ghgu7j+7nxXNEmE9lIg5UmSwdt4u+joC2eCnSu10vIHLeIV
Yb+spKW+8YNZYuHSS4EhQrMFYlJxVPMQzQwNjI8sngurvZY9aVhjnZ8jq3nqvzzqiRJbL7ddifsH
3TI9erAEJHGHAcpcihVsjVK/8/5PODZVCW+9jFVyynTokkfxzMaRdG7rwfRr0gogQ81dGVGR3Vt7
iZd6LSrBIfdo/gmMK8lXZAmGo8TC8KmOBtKKkabBgMJVnVEgyX3uSEhMXeYoQOiaBW1tjqU/vPkg
f3trBXbU2gL7NBWsVtz5ptJZFLP94QTx8kwKX/t1Bo/QApyMK+/yCDXS33uFkaykJsGMQE9gBoyr
8dSP+aqwtPBLtsaPJIEW3IDCrQVn/M29EjGX62mo1CLTzQgw4bBHE3+Yh4cfdXSShTkaOZabIkAD
lqzojItf4gAnamqmLLm/RoNSNGoo2LH3bpRZlXsomrIZMxJHqdkYWCnRs8H7Xwlbp86ww4B90PmN
9HU8zfUyLdgxBZGwvI6BUsPpjwHtPe5Qp3R8FXWvn47pTcSTMGQK08sH8itDir27pRHbeU/ZXGHd
VOWzuIlMX3Ib7Id5qiO34pIVs3ri48VlixFasyt5ECI34V8Yy5FSTuMsraPTdAeYw50+9ghrk9hK
AWZj9dUMBN3gnUfLAFbpe+N0wINNzk0h85f9uN7MTLEy6u9GxeOHttJcFVys/ciNKECKA3ADRW0w
ZpGR4v+B7KaSPS0Y/xjTzI1acE88mYW6nDmKWnyvPT6GKK2oQIZ3OL5nkSgcBCu4PbBXoVWkxdfu
3nGRckfxJW9Jly0XLHXYPR4e51XmaGSjQFQX+X71jvqINkU/cY4iayZnrHUaIgF7weBxMdxhs/pl
bXpz5fh/5fYlM3lyKTJJPDD77LYarghbYAoT4ME2shsVVRGom6evdXK/dfqj3HVPVjuCg5+hkHYD
7/DUM13bOp96afE9quw/p/Ur1pXEcErjCNZjfUhEx+m6yfiTOobXzAnwrWRzE3dOw7KzmmggLs6/
wK95QmWnL11S2QwY4sIZ1vgSJyPnUcbLSxGeeNkrmKDxU4sldfwBeikoroFuJv+UcfC4n55cwXK5
jo+sBhBcF/0PL/AfQo4Ld4P4A+ImgNSCHx9igoFnu0BXQs8vkY5ff7eogRfjiX0pbcU4CDu6EIeo
aklywYkcq98iSAQhfAL1pvtD6wvGrdQJYxrqpD0/bpEXpWfpZMOrRMNtlaEEhpoIDsk0TS6b8xw1
zU7pPbvse4W6h39BtHPJvzhx+zU2qjELEDJTxo9YlpnAZl98/F6qGfWWce5sZXodfinq4CfW0Nwp
JDDeI/7LP1aOCa1RWMwIH0bgGSgQeMnCqsW7NLeqAEhZIog34hPG/RdOmEDQzdsBSGeeqFH1ZWu6
umthFb335onPGolg3zvRe3UJAHJ8u/ZuGaxOK8aKzlQVFYxAmkPRoRD/2g4rEJr4E+hK+95MZjP1
w/U24nKnzCKgsd5q4yhFRO92468DE36HXgbNpHzOAh2najSOqYROOFz0wfPQF8hnw2nmu5jJmPhJ
JNARssjsBwkSQMKMOvDlTw2oRp24Ak0BcQ4sfR30sv0CPRud+urg72mwqU0EmDvn8+V+Ctw+x57i
4ZEXokeBNRlkhI7Va2xEuLDojzp+kMKMv42eEgBx/k1xnpNm+uUF+4GVP3daa/e/d0UK2eVajR2M
4l4X9Zl4Y4JYCA0bETFur3Aza+qBjJj3HFGw1V70B8Uix6e2hQWtWBBtW3fIcMnl5f/x6ugQSrT2
/NZG1Gn7V8I6Id2bG8yUK3Ot1R5C0/R4YqskvvNhax3g/JAKbXH/iV/zmdwOiQWN9RjkRVtmME6h
KFSviGsVndA/PGGZsedaPMYmo1RRC3XehMgpdTBXn5AlmU2F7GhHoUhIVNE5zXZIv9FnT4nBhPNn
UPb7TIvI0VfI0e91fn7N1hxqu9o1cnR5M1ddQ5AfQbCxj9YjLW15G/ySrmoC31tMDWlmoGYBu4le
FaXGA4rqGv/Rfea7kzMW+XZ8J9v9vRhjP4VGFfkBuhdJrlyECskg39La7lkrn1WEmDq3EjvVsLNB
g49IWmCu2o1YXo5lYxmo9TN/ytLG37bcy583ksMZknD0uaVV1XbYNbW6yAfrBzRP6DGFRB/gINSg
gZVk/qayNok6mzO91GmT2ncnWXhFNAZbZ3qiIxwl6y+noosEp4Bno4wYGoukZFIJ26sCXioSxgkX
tSJzOVpmVzXwg8Wo8ycMa8KxgUAo+X1n2ewtYGa3pBND46oJCDUiQNlTIc5XbZfnWN+0NBf5rqiW
zi9ZkVsSraFBchzqLmCXsQiYMpAyIm/sIeN/s80dxwOed331X/iIzheOHgqX4jGW2oPhCTyFSrXp
9M23ainuLQ6PaUamXv8OtDv2VfTkgJPTcCjeC82SPbdDFpkzZ/ktMgvPAFg4yREh8S0l/mhFdOnG
Th7cTcuXckMDSB2hPnrGze97bnj5SVPzwSec3B00GYyqrUVLlNm/KkhMYLlh5xbW93J2sfmOJaHi
k567+mbExrCxmzACB1K7fH1NU04VC/4NXWCImN4qIWcEYLCMollfuq2IE6kUhL6lZoYRpuAsqDc/
hAcXu+AeWMQDWEQ0SJ/ml27dMrdK0ivRVNeiI5+E7jXUmB9bYgZ6WpGm6kRADyViXLCP/9/cmMFo
IvkdrzSj5ZvykgIbHfNBCQ++OPFxpO7+GSFJbYYqwOnp3KJngGyKdM/A18divFK1rBG5jovQg9d1
jVZ70ukSLHxJEAtw/5aRSaw89PEnvMF8igw2i20Q28Bu6cQgx19cPwn18pWJi4xHIRklmGWt0njJ
4yE6ivS6AnwveILE+R3Yz8RE4kTk0HSLE44yWRKX16ohGSb+Yf5ACnLiMrkruWxoiqmYy2TzRdCc
mtqggDYdhkjUPclSvfYHnHMZDcgFsGdvRb83suZnSe/yF01HfDOEqMKTbqkygqovdF89YhkIkSzO
u8rAMzaHzxE6JgML3dEI7CMVvs9M5r6dJ84GGhlV5nGeb0DQTRXQyh4weyywbdn1PUJNBzTx9dGd
ml6ywSObks+c5+TGb7+7RkloC98Uzkh1aS+ja8kkqOuFWp+qmomwGCMQHk447nHSBOPoTNo0/n4G
0zi45p3aDMMTSxm33qQT7SQjq2IqyA7uh0XOrIehuwGZvTFHJ0+HfziOVoEYsvbpp0zGjV3nKLX9
xdY2S6dyDvfStADreIGiYio58yb1DMS19dLHLDfry0EydZl8pT5vPEb2MK1xEWrT6+Xxf4/ufE7H
kt6dhsfl4mzO+Jjn6Lzrvlq+bBaFYp8Av1Yv7E4xJ/FVfXiruP0wFAJbwyrBIh14Azk98prd2rcW
Ylz4UCH2GGpUTZ4vu+Yrtp/xnlyd71DL5nGfAfO7dOjXThxZ1qdN39F0Re3plmge9YWGq85WKEAP
HUTICEMhu5dMynBefof6VNpMWAXhvZn0C5kFFZN/5Bl0duTiuNdAxdjK4VSxO/DWE1bp3O9Km1J+
t19eCSaEhyXCkB8S3q+Wfyyt2JeJkr4rL9zWCkw21wlrnSgsq6eA1SbFRdYUfsUvc3xcfNcigGZA
ucgfZIx398WqPlPNBi9CrcEzkXLV69X76ClHurja+sE5oD1On0q/KIPwvNYVCY1aU/KXTgH7/z8m
MBmQ+ERdx0vG+Z4NKz9ybQdCu6km0zHRQZplQLlRmqBTmtay+r+VhT2eBmaojPT/SokUWYqdlx2Q
IBgOBVETauohfa45QEFWLyLSoYM4FD7m7aKxSMx7wetT8Wbtmz4ufQxqWf+PjKwxvQPIHieMxxtE
BNQQoabawpRdGT9o+a9gv51olsC7Dw/d6BknJgve6z7zzR35M/ZtIrumdrP+gsMJMqk4U1jUy4Hf
QNk2o+BvZlVttDiv8vqiAY569Z6IftySStTi9TyyN07Jkfcx7+3fEC3QGMQVCYMsBDRDsYYsMypB
KWbPoyMlztAPcDgIpjI3/8ZwJBYxZKS8YW4UhQnPPzIADizJi5jnt2mJjybYsNVHNsPv/Y81guvP
apOzWq5WDolFTrsCM6XOKVjEXY4d4en+Mfb4UT2O4wwW/REz52rhzP4LJZQGVHflqr2QED3BiFaC
5csXPy07Kw3GBz3CBwMZtIT69V/JwrvwBLqZuFNMd34eeXK8vg+ZZO5w+VSJXb4CQq1jsVuijQp5
poEbj6qZvzG+XierF8ebQ7cxaSgCpq2TYfjSW+2q8iJOsKfk4puymGc3tQ7uBeCD+SIJWHpoEByz
BajATl5pqk2fFywiRWIh+ibICxoVeh5pybP1Y2IsRskgulcO+jxbYW2Ej7fyHsrp0W+/hAG6hPv4
OfMJ6UCFcIMywAo1vR3XkU080/ARp5gJAZATWptFKtO/mCIn3jK5rygyH7RW8JiiUSwYx7HMyxfo
yGSd2wy1TJqkSMbdPVTaZsbTXCF3tzF4jCnb+Xgp4ERhnZW5C+cXwUaoTB5ZLjf2+L0mGtTUJ15N
jq4tGniD3+Q4REyFAg5mY3jstZD23Zd1RCwXV7GHG9yPI5thzOvQMw+GgRUlRPY0uQiCHsZXLW6u
qr/5EVf2bUTgBnHYvXBUyV8jfoe+bVq3aOM0IWMI+9Mnh3JIXT2n+438gKr4BiA28jWdoNi8UWNO
M6+ltXDt2oTUPCuq4LDNJCzfh3WL7Cs9KWG4y4H0oTacWktn9tn13vlTQMcdZ65/FzadGXL/wI9x
32i0zhiRupENrdsY5Vd4xwCRJkBORFe13w/qBi5u6CIZaFC5xX5v+3Kf7CbArnFdYA7Qp2ckIVas
o8quzM6eSUBanA8N/kvrhiYvgGpW3DG34LuG3fwK2V9ysjuyCfFAyEg/z4GoE1e5zDtbIEe8XoZP
TUHRnf61AugOLU7jCkkOqj7OfJSKejUxqA+O184ZDLd9HO1dPcy130yn4L6FvjwQeKwfC+nk93qT
zn+Jv2Uhj5cm4J6ZJyecenLm3CtCfyX9aB2O6MgmnQU7tEsjrpFmzDcz6KWJluE+suJlGlAylUOK
4i84K5SNpc189cuiGqxsaDsZ0hpfO9l0TsX2ssma4HzuCCxRAkQBptuRjVrk6Y72vy0kZ+9wgoMZ
dvZ0FU0J3AXSEbb3MXVJAe3+aZ+7Pz4TJT9iEWzHPpQKruIBF9jPlvXbs0lBps4jkJ+3IH7W/bsa
QtXOQeJ8pwDaTimr6O0KSUnEnf26UE0fydCYa7u67FaYUppxHgYTR6WarscKwlIMvZN+vQAwAKuK
PUU6vHN1pz2sxWg21uHZNiPfP1cYRezoU/qawTgkbnWtqNa5AjFXDYxuaKYv2KtlWD55udxvLBYz
sP0Y0PKM93DwbY4Ml6g6xw/mvixoF5AjGDs4eylbzsJqB/Cbs8Dmo6cLrf6ykmwIYP4quEvjUvVG
g8jvMTViaQLbuvQdsIR3rBGUX1BFMhQ2o4Dj4ylkuLaDb49qhVDcjDhQbqeSJT7gG+hq+Z5FGpaw
siJrIk5ZSzGOjjvOwT8L6rFaWRlvYSgzVwHDZ/r+p+EgjTRYCDqX/0gC7mEWmfsXrYHFTVX0v+ZS
pBizYYzqvd+ygLq3vRSk1Koa7E9t+UutbMMc2+a8fbAWkaMgSAFuuq3KlFU0BnhVoDRKeFmx13Pz
uwVVzJQyTq3u2IYUbJzNDxmLlg7AnBfG7hrz1GuAmqN34SYhawIRU4qjFauTMPNFySVDH3Ze/R/o
O4Ra1yySiqX2GjVmPS9tDhsjt+Lu1keFaHjXkb4moWMjP3Z5IUkNScuzr/OcaM3LomvP3yyAeVN1
wJc2QpD92ovJE1nXLo1rBBKR5/cscGGLHab3FFGTlMAp222P8DBbE0Ong46Nzes/ZA8ardQ+2As7
L9ckIOFG0PXgrfNYErUCHrwG8xfLX9HMYPcIILUC3BUazn5S51trL54BU1CaqVIINgv5ndFXAs7v
ZMzamPQ/8rhwehuWRuFrB5rslVf4br9C9yv6A5MLIhJEkLwSXrGlldAc05mt8pj+8Tncn3NXGJZK
hZMepE31ISBqFUOJxgIt+FbOU5+aZl86NnAn6udgNBJsHF3beHIV45AmpF8HjrlR0L7hE2nFsb9v
pvYreFvufM0X+dTLQjXmAXqaNk5Z1Ww8ZMP3GuYofnVEolG52jaRNd1B6RYIDOnjLVezR4F1llEm
qGhsL5rW9hk29vJb1t9UpjjKr3ZQXmyuCj58C1dznkeVxZs8YivhqKKLMwfbp6tFE+pE7tHWbfce
LSXWg3Jyu8YH+oYKN0DoHEE1FINAbFTIHy3UZRGRn3HcWaDfLAOWTIB1qfo2X68u+s5HmN2UJVKo
YQAnXE6U1SvFlUXK7cNyKo7xj1x6C/1nXD165ejkXX7jZYveZNQ163Hjl8j1+Yj8Y4UXjWRmt9Cu
KmaT36w7rQXvL1cjUhPvgX75qABlT4kAPlTism+aqvYzUXrXVqjLTOjnNvXvy6cyzUj00c34ExPa
hPwCnPqtP5xiuYrjrmeNnS0KTDTfyLhWlycRrpAQ+SFvlZ+XheJbT07Wu7O7Wq6hFJQ/dgKGAvuU
0FHpBxebPStVukM9n3DJp8BCUH+kw+aApI8tu4+4KuCvzI09YKQlllUwnO94I46onb/k1zWDE9VR
wi+FkBMRXrx0O6zy3d0W/YF43r4FxZ7IRMPoRY3cAtG0xeV/FXzDXY+v03JgJ1ejX2WsiRm/aeFY
lN16JBGV/3fV4G/hUKV3HznjIhfaOborbxOaUGTqdTnLth7OaVLJ3YWnPW3sUVK1tr0tiNZa48an
Woh8xNqsLx0TRhmzfWdO40Jis1AqvEUozfDsQazPGwPRxGzGgxpuzKYyrL6tzvqpjb2iMr5OwPbt
Q2PAyU7GMvm7z9OpgLI077dQCH9xH3tvjWYTG6TkGPmN2QI2PWMK16lE78xK+/I7ihMMJjuOgke0
i1oaCteuGCcLiH5UXmrhInkmzgWd6kWC09uQPc+2pI5oP2lSQGuNz7kEBnEMH/5grZFWmSLs5ugN
kbJ8iyZ+oosKqfZU6FI/wp9MQYuioiP/m37Zq/7i4vpV/DDiPKgXJxZvpqg2WaudTMv2W4jXO/q/
1gB9rsTNIET07wyCRtZpWK/37ZCeVW06AXOfpp1WTlX5fbKg4+6THVGkB0YQMfHCvdEXJOhi+oJG
EPE95QbObUv7vCsxbFYTMxnjrWOmOujXYQWei5tkxPy/GAQ2jF62Oit9/Gs2l5j/ywf4nAnzR3zO
45vEaiXpZHfJfKSdPsV/ybJ/BQH1G2na9/K8eaIL34b+8EUVCn180vEtdLFn4oCGW/qI+Qyw3Dn0
wE4puANVJUIpoEhtoMohW5ywYuSukkMvm4nC/PoTrKqi4pwGoaFd5uZKn7Znwn+HF5gBJ3stM1jE
wi+77B1bNs1bpDtujNw5O4b7z4RykJ3JkEHn4u49QAcyxEURccWeUyIcmJ/DsOhY/bG+0eU3WQpj
o1RL3dgcvHbgB1kLYDm4pyspBfGHx/TR+xQIs4NUR9nOy5hb54MRfbIYzZwL63ZiSDBNohvTxARA
Jz+7lXM0yBaIJx9g6RWnnm1h9FR5xqnZxEMeL6H7uuD+Kd+C3bTJM+mlj1YJTCXMDghI+JXxgNS+
2m5ZdV1Ub4T9RI8ZocrAMb+zTJ/SfY2LU/I1ud8yE4lDXtru7O6Iy6OHCMvlMGeyghnrOS7hz5HU
Ssk7V7KAPdkVCcWPnfadC8qPTIzRfIuNoI2oJXd7dkB5/9MJmymLordXsg3kOQLC3aE0JjaRhWme
DTF0hDin33NeDMJOPLhpZmaO8fBasu1o5Ouj7nZT4DUN57NBkQOykduKpZpxrA3CdtFpwBV5UwQA
Dxc92UxGjbL44OHq4ZREX4ZD0WGebyk1TnXYRyImq/0NB1NbtyFzPFtIcz//ekthbj39HjH1zD5G
yNetySYpnxCSGj5K7acfKE/dPQY+NAAPYT6qr33aCFIlPH+PmX78SLNjwhB5SDWd1wdzPxLaras7
q0LE4k+3Mw1cZu8QYciv8pTHws6a+lDEfPpHVpRnQ+belZAWOxYvO8amKsF34iMm8JTgCuFckhST
FgWyAc9WxVNAAWhPrwjO15LZtpW5/bHv3jXSUscE647gN9E06T6HIaJXL8BO3AO6ootSfHnBsmCN
FF4hB2wwKBG8Yu0JyeyxTmSKJQ9X1cMzp/Ah8/IyfFRVJSAXsxMHnwCLRPknOwBD5YbEawk4xlta
8DIbhL092C41DXR/xxHBir7xH7MmsSSbENHO68fpeOXl0HaGtYxwRnlr1D7oPffQ/NPEnsQreJOf
66+uxdrZofQwE4K79fTNUNEfU1qTq4ctWNi5RmvuA4rMorCrpvZ1m9BcshaxwRE3nUDlO3LH/gMH
N0QdoizOJ17Gwmod0/dCyra6uC0/i2a5sR2sY6qO8t8FdPXlnQrLYLctCIMDGsjW9jL6TNPuxGJ+
E4Wxdi2oGYNeomn4QpglWSVrUS6XnRhrDKT8EqmRZ15+SyQnRkzS4p0aM0FWY7xoMfE3cNuyGDKv
27wHVpFrMuk5ddhWM3K1NXtHNXUVdBJ+YU6EvmCV1TYvGiLnVCi6h+tZOXEBNKGbplUm9XLtAUvK
6x6kwQhCtH6K6NMyi4PRmoRdXUIwLnQTJ2ev4bVqcGSgiVcGRe3Dbke4zfYewHQ2Jh/1dJUu9HRu
cAoCci+MEAM2S4S7a8zRR7C+pJrFblNFyuj4h3mTBrdzDRHq0FskoRc+REqHQYXIqk5z3G9xjedZ
njdE1os1ph+CuHbSYLcupf3uaDgfbMYCaoPRtkDGZYoU2GwhWmPfverZdzd1yCHVgsako7PA4NcO
YkXN6/48hQgOU8PQvOKYUSxyfZipU4049fYQh/z8EIsmhmHHvyUipaa45xE1AlyQv3YO1vXUNbph
neoYavyEHLBEsAdt8Tnsysv8Cr+0RlyMzAmYzgnZqoBdWO898fG5UBxSHJ0qwjONK18DqEtH9yYf
gOJg64jvIulDvI930343ZGM9Ei+amwcHmM54vUnQaUosqjanKyrSVuEnMp/BCJF0tNBEs5/fkxt4
vyyhO4VcTeshvnvwwKRfSBRCulSYIFjv+uK6QtGby9O50cetiKIU152qnMVuzSaCbOgshiVW7llQ
VZkzfHBb+5EjwYF0oMebo+0jrNgtvn7t0RG+E9QjJZG3hzQIgtwYmPXieQazTf+QaT8eb18SKFf+
8zDv2RVwvDSybOJ5xRAGx+KCqjz+YAkD5mzSyajzplEZejEC9pzwzsIfgmMIBg1OWEI3eC0EobRb
4CWzW9zH3oSuKs/Xfd1aAJCfKIo/IJ8J9/J1qoN7zjgNusKjxz6bZ/EZTbZaYeuBfrafvEdfMVYM
MhJVfCZEg2S4NYQUhlcz5D/3a+kRIB636cNpvU962wiNiRjzmTAMZWDt5ybVhuH4obgyFZEM9jKJ
4O90/UURxikrcUxB39nwM9kbmIK2l5ccnkmFdFawT5baTv6OO/zUimyZaaJ/tTF5Cm2jEhajYGvE
0JnTzGWWRxQy2GQtea9hsu5LoVBMzNtdO2ZFO7E9Oq7I4LWOotK0EWSH9wltYeHzbb069EcrutiD
6slKR2BD081+6yam/hgH785oHdyZfo0nqFhiPcv4kg2OyjY7YM/nGptUfF9fkyMPEefz7rwQmghf
ok2pkxmx9kXQIjzWCPw4PGz6gSq65RikiQgCAA4VvaWLkTTHryxo2GF3h96MqeNRO3DboKRC7p+Q
JW5pl239DWKhtybY/9flb93Hl9+YGe7HbO8FWR+HEPef0vtPz9nSfHoSq3zWCciYN02Ra8z0dD0x
EoTvP9fjQcuyy5g/A0D72WLGODO0Q4lJm2XT5eLlND+670JWqFyRMjHlkcWRUkWH0RWcdOUf1JBF
QnNUFz8lQr4Ojex5Gq3Lou+Mfaigvnq6HNzxzRWcSrxgv69x+/bIK49JJTUOlJlJRsD08V0lTou6
cQ/5xSrY+Uw9dWCL65LL06hBIqFHtS+kIEGgP37v9e+W7F/eRsnVYBz/iIFJoCB8vi9SDjSyl9LW
zGt9YeKERK0/vmaZWvxC74Y/rizB5SV767BtXzSavv1WKuC3THe8JF0kd451+xlxPAPyyKCowPr+
ki3WFZRN5u4IJ6LwsMRaEy5zE96Bm/TMS8zyRD77TRHQhAex4orWfMGixZxgWu/wR+oWKZ8df9fm
YtEmrWVcyn48f2XjXVOj8j1mn//SWbS8vMfMEjHlbSuLuWhDIY3v5EM5zsVbdFXw+OLftS3CoySc
XIcsYSbGbHGsKT37JCt4kYwdOrIOWxQyxW9NJzuLehJqT5En+tXLc5Ql5MravJFYVUpg0hkTIk2G
aI5mEfstn4d718Xaqh9BPlymzL/V/2pN3aNYHQyzM2jGsz7LahFuUdGBJZZcNEpKLHUANpwovkaP
5hHh2+KTw73KQQbYVc9KSu56OZ6tO5MBdacoD9HaW+zEVHkTEG2Bwv/ASsm4zkRYdhPN9aGyWZCW
s4B62bUPE5i/1YNlCw77ix/Y4B+6pdCpRlrHnGM6CnqtMkO7T+SBNxXmlHby4EsUMt9tpy16XACK
SDo5UM/309Af4VR4pjg04MYGMiNGHoHC0mXZhBQ2SeWqZqhCgCe8N0mhxF5zmQxBptc8r+k+7OT8
Y2qXW3WeZN6WnKkh0NlELIzFhWHS8Q6XxV+1DT1WnYm3l2wzEnEjA+9HOlI3315d6dyRClsC7jvV
ZZiKsH243RhQQDeuypO3T0aMY8KN+Q9Y9S1ssTlMzfnKPGSR2PHVrIWBZQ/4wLvgHPSufiAm0zaW
itEPRz8RPks38f3cXL1U5yrZFfvpNqJ9X8vUX1LSEHdgewf+rFZi2IVDXnuiOS7+yrpf04CPx9pP
Xwucs2KwyIEFdgP+BL8nybNa7OttDkQoTxcScmdRsD3H6qfpcywgbgPf7ySl2lstgbbtUFt/QtEO
p2GsEN7bQ06e2doreqQ6w6U87lRR71WHeDwKfGF7+YSIPDTmC7CE/5nw8ZBWzP2P9yFXJrDAjGVz
ntQyaW0d84qjr9+EeDfChXrHuDh7FPqAC48ujCO1b2nTye7A9huMKDM01Ku9nCmhypQXq55P7m0T
x2bXYE0KPuaXPFSGYmqpFPm6vyDLjJYf5ulWO3EXYUCx2seKwncfVLje/WtOolrmz+3tk61palMi
qNOnNg6EifyKXCRDzaGkPhv8E94QnFgC9rg5uf+X2MEnAvSY7C1xvjWY9uh3+gqH7V2Z0cUz2Qlx
o4RbZEwFRlDwgJlzd94hkx2JiHJMTjazRjgpTwyhleCpgPSnGRtzWavlu36ky0+ayBgg3SOvD8Fg
/zqgGvkqgOw7WggL5ulzkDnDqqGCNSjT/zAlr7A3lRLXMIFKiSZ0g8fUDbAFetTKTkHCkdljwmqS
uba+iRfdT+TIMJxLedVbrrgM3TUGwQxIBDX+y7/27CW+1ncK+2lRkpeHUqSgwoQLXAy3B1ljdp1L
q5ypcMRzydetjgCQmANHUApaJGlWCSM3Lfwd0F9I+APdGiqQFDmi361jdkmhq4mOXRwfVbAiYu1O
15mQjTuhETiomUzLPZxKHX5f6wCwaDAEGZMJVPPrxEK8DDVALODS8y08i6oXaBlGU2vpqBFCqgk2
WJEFkRQ7Vd3Xz9MubI4f/93O8MgwMIl+3UKHosonhHTcJ8LJXDaSwBTtoufw/P2zD5lZpLoIVJpb
/OZLYfSWGRrrPz14LR6s0JfXOkopDhW3pvIGtpf+/rFjJi2NjEGQfW0EeWtx4Tns8CbSk9sYX/JQ
ZOumMSVF2AFFEw+8uXn3KDfPGDBLPJUAlym4Hd+ndX6dByBJhIm44n+rtKMjwc5hDh354p5DXiKC
GcIJeSnEA5xRP8BBA6sXNgqNfCP9bGZW1+1Hr5A+KesbNnuPqlyUahNIg7Yq4YgnYB+Ni1YT7Xjw
aJCN5vdPeunQTKGhSSBod/jMJb+HUhfMVSGBKQPL7u12eYiEB5nycbdagM5IB5lj+xBjXyzIRa3L
xjE8lXIsBY9WNrIK5ykRZIOrf6JdltJgT2gcrNMgvwbDRQukTcrWZLrVx9nwb+5ks6EjR0BbHb8q
R3AA+58WVJIaAkArHof8wRY5FZ2OUkFYpKgA69EBj1Ccts0vjg2bAviSitK7MBpRERLppDgJ7so5
Ta/+2rvxITXCLhq/jQvn/oeTNpTlPu+CLUsZ/YWuNk+ABoO2Uz3lzEQ8QEiQ4yMX72ibvgJejUw+
TQTo/Pm+gKRv1NcVvrK/sK4VZ6kl+eY0h34es3wOlUZsVld3WsKbm9jWVTgqn8aEaADQdDrzPvrE
ReyPumweZ1owSBGmWMazMQBQbMCWOueehQyi1GTgAaaoqM3kS82gBK5PK7C0eT1AkDPADM2lGjh+
gXlgc4+6mubA7UqVSxbCHG6GFm/FDLhiqDBeoKW3wVOp7/mI9f/FOU2IR/uUNCRMexdqSmXbnogn
OGSB3QqhGaFCsruw7DNBlDL5OYXEtpTCeb2q94rRXeGGLek8UJo9oIuPw/mz7n8aRb0rYML3WQXS
fiBke61tRD6iezx21TKdMkaWXmqvq6C6qs+ezbANddUhQ+KBYB1r8y+bkkdSeYlQZWfTlIfH/4X8
V6FGBOTogBjXjrSY+GsiV8BMvrgq94g3p760aV6qoQmH31gcR4iDw4YgrjoGJWJLt3SwrrSfOkK5
ia6cJj0TIAFKLNN1DiXobC2Hx1ps7uLzX7NlTn9bGxvcz5RwRbFlk/4/w2jeP+EBJKqyvMGmE58E
xbSpr/xi2JeKJbK+IMpnGAzx5/iyfOEKKzU1bt+CqYuxc571ZL/2A5Wd3TUro/NaiqL+9j6MwLpE
ox6rTe7klo6xXDjBcAwNievY46u7FqMyZ5OiQHnQVknLpKbTbq1Gsd6ADae8W4vImSoLbL4qhsQR
/yqPOfkLfY/wcmSWDnMU0CY+Li4jt81uIQy5Ja8FCWyHc5ovUXtJYKzQ55cHvL63CgBGBNkBMc4d
BZJ4X+W+vqyuFLQkwT8D94cB5voJ5smlLzhclhLzvpUC/peOzPasR//gOMOBAOp8az/aH50Lm09l
QkV2fVkXEdN8C3E85gbskdebkonvR4DRCiTT856D6FjuMss9DkvwX4Kqy5Y/kL7K7dR6WbcKvOIC
Y5vfyflDm4u1pbzQcVNLYiM09BUPdzSeqS3iHu+ROzbW+gSzexiQYuMuTQPTFhXPcV6WDzHswMMA
v1Iy5I/S4jpLyEVdIgnXop/fFrjif/7ebXCFnJKH0d+I5nBlnQV5ZcwLIH8otEm+XEh1C9lA4y+C
5jGZeAM6XKeEbBmISgG4EU2K3P1WIw7m8zYb+Pu8zrLOPzpGg+Yh9trnQ/WS/yvrQAyRwkgRG8Uv
p6V/En1iqs7PUW/J84EtmZ/Tdsig+YDIBawa/9ZQdmZNcmzg7za3mTz0m5v1cMV1yhmh0glqcyW/
7MOjdhj9Uu5EhzUcLdvxwvO6RDzyTzAkE4Yqw2Ua5C3Pa3Pq/jfKesG8LKaQBlezjVWs6lhBiHdN
jHXrDfNtcjXdWclT7b37mLFfEiw+oHuzlvBzlzUu6xjCahfyN17ywD2LEx4xOkP1bmZDQnL03zOf
2+P2DkKoCItI6TCGrWFEgywbwHA2K5xbBsjeCup9LoPNiua3m1hcqCMepn8ZEyE7jVH/IxZ4Kj0q
IfTZxQLntHrK+CUAKB7xnZNU1n4tgFTPdQVG5a3rFUHaxt/erbl9eu20URJ2TxIB2gxcBb7EI7wI
hmkQr6GJf7oEnleJluF7NNJzbEG7cvb1Yr6aF2qAhq4MChlITCzqk+TOaIiZzNTJUSM9YUaOZnfp
vCJ0inXSnu1CJwdRJSGvYZWjK6KAasHAUQa3uTAgk+pCZjZKl/ERjqh2Z7M7MC7EegNdwaKhqCA4
sbuXMfj0ukUGy5RK3RNPtszYfaqKUMQVplFfjnHTY6i+o66rOjVcQBu6Rk6d/tljrG4S0PQdysQD
Pi8w3/oFUmc4txI4d60bndXefEOfni/zGv1v/bRgNmANoqiZQF2BsZY91aS82zZXCbvYPDRVCVx/
DbvaGc6eFoYkRTbOHqWVc24SBJCwLJ3C2hrXoAd6E95JLzjlxoMPPMDlvnrDCH9/79LQuj0JQ56K
wix4ft+PDSmga6fZ5c1lFHWp7A5HNuOY7q6ahIgf4RQijaZorh0md51L2r99MulcYSqxFJlcS1yE
rQbXFsdNCCntGBVeIWCH6iqOr3TmenF2CZUXiYVAvRjc0B9oqS7BkKbS59IEhrzq5/HJX1ozqXo7
HJYRvKWjuBgFibN/KUQNy+0Viaika1b2igAqbrKQG5EdGRzYnokrl64HZEEL7JzKmMMvgpF3wcsv
ACYGrsNPWfX9gyo5kCNDWYZwj492DsXOU1wBxPdF5/onOuDd8iApAlwjJ7dwfR3KX1HaZp2vwgQH
5IkuQt1Etw49LIZU1eR9VPoAEkY3XD2yhc/VbjzWYw9GaqeJPd2w/D0Rmllsr4wj8BsbSOn+y5od
V3z5gGennqGlAuZTw/x+Bv4ooXayGVM+xH2T3YeYpljns4nWU8ZYQGGgykWHkWKmkOTxnDCdS1Nb
zoBvfWpmLl9HJD5jf2wnb+E9h09HUpa92lFTxegEfSLKc7IBiwOCbT4XE7ICSUZ7SusaQ/HgsYv1
pGaAvm2G4j0oX5FSsjuvRaycJf18e1WJtTAb4s+MBZuBVU9xp1LyIwxw/jYAaNyoPPk7fIrcKMXf
g3u6CZgPXN8SY45aBG3BwUU3Actu1roEE7CqmEwevCAHG2qZilAs8fQLyNAgAWY0H+d+Da1KC8+Q
oZBvdXFSCai3aPPTo9rBNuaRUsx4eNY24j8kY3fhkM+7/sae77GIx0aC7fmxaqeWHV9vdDIjYtf3
VeFXuUL2QGNduBy2uKiX/7t2eHXIlefQzr6xdyxEgCLf9Q1E6rJ8tKZqQ837fKNh/1RKxI7EhWHz
Tfu0NnW4zJObpJGltlUqVy1TOyVmXXDRkDBRgIaJV/d3P5tY2iHYCugNyln4UorhpgvhcJgzz458
mtDOiiWwZ7whv09Ryj6Sa5OYfmix+OuWGWYBTa+2RQTdSjbeO9e2Q0Vc+3DQ8r9Szi4gNp/ixi5b
IVi0guUvJh3eWF4oT3krZZ4cdwnv8ndp7fA4WMN2jpgdTvZBVYkzbgBFBvrsR1HE2tagHGLzplpC
IDwpgbuDyUDHNIiYrk6vwwHCs2etze9xf7ndAHCHHsPqVS5m+QpPiOnbIBFmKWJSVUGKLUArfxtI
UxFSypqN9ug5X3yNhPzWFq8xUlRZjz757BWIECFayMO4DhmyaNqdFLChSY8PQ26oco0Powvt+8ta
0AzMjAu5A7Mgce4Slb7tptsxn1cFEm/E3sTMr6ySoDsBxfbLVIDgRmiEU72FtkIf8qBeDy866vlS
1Ey8q1+YhM4YovyTbDko9z68BWbsaGhkrlHNBddJgw43WPRGNguzO/TVp9WNgFnZhXwdM7eoWgQJ
xTvU+6NXFOKpTkIJMzLJDwhiVzg21q+UoG87/2jghUeOFm4tHnjIsTXgAccAuFZMTinWsuyMeEPk
mPjH/LgvoZCAw4K4xA0E7LMgOpUJiexRYT6HFpsG5+H7STHoMlB4wBQYAWYKpRHTkooCDnSomsyY
q6bBIuZXhF8dn2CK94LPg9MlomPCZbkIXRnt5bGM8ee+tPlfKapRWw/KpcVO+JMXhuP4iGolkHiN
MEuQBeDr8jQJeNOaphTFacrvJQe6F75AcGFp6FMpAMPCBck3cZ4YgfEMr6jZH8AXUtRiWytvc29W
t734w/f7x3npiPDvBzNZzwcZqdu4/bXghXFKnCBh2e0db6uql/b2mc3hmcGmrmy8fzOx3/w3sWnz
O88ePw5fvXzWw6dlAsUqFPogdVxjRnaxSQEdbl5SZy0C71moIvtACLFma5bMzNwHFvccDcZTfgUr
C/32LSMumU7G7xNqSmuy1luqj+krovyNLZjEslpq4yB0SeUqMFvRbn4S918HuFdvRw0xPFhoKSsi
3YP+uBsbitUwFpGxEOn58wtVyngtl5NlSHCk7fZH9MsjEI0ISZ1mPZUyoi+u/PPhth+trRSkcbeu
zZyJcRa1lAo14GQTjMh5Pow1PC6liJ3QSmOsktihH/NzNyjH+wxTsxQZpMK7PasT9CsxzHSA/m8F
LOvyAHtVJlnGyy9Fhn30G7uZ2Y0/rIgA5nsY/fdZkAqmgrz1KLFHWEiUDXHKm/YqJmZ605tTyECo
DcVDnPSV7UduhmWicuUykKZMnxj2U11bk7xJx5Uvu1pqpuWPeFldK/NOsvk0B6cIP8S9SII0OrT0
PmX53ylSQEtAY7/lkz7WRa4bg+MMd59hiO3KlNkNyE5D7eggdtCsRjSwhtmxEW5s5jjW5FxNt1T4
RqwFpp4lxxL7AMPmBuv2di/V3hK0xnqWdi85HQ0OdYj9SFRPwoaJKLbbJ0Q9nc3EbcfAQmVqFArI
/6M7IU52vNDAcjGrmFqzF7mvwryxQUS/y/LxgWMPyAO0I2x28qyP/nC5Y2p7XcIsGjyywYvGmFZf
pRerFE/b/oCY8OD4Pno49DMGEyFOC+Yq1yV9aVlHskJqPlduVYfK1kFsVXXea+SB5Aa/Rmz/PJdd
Y8f1yJWgQ23IxFHiHqD6eqcB/l2e+qD9v7YG96Fg7bgi0k5BffzuiplG2PWiLgOLx+UwK3kQuDbV
wOfSYEaCUsmmKwFLaIvc/++RHSakNmquNYel/zJpNXTrdXn/BOvtRoeg7hXWmYa7Le6qYyFclIs1
8aO5DA4XIIYalRhdwGoPjWVIkBt9spr3TUsYeWh5oMaVZzOcRoB1bKQl0l2I72x9mQ9XQMrjPyT5
sjIYdhHmgYPJQDBOMBt29GyZ6wFigCKyh6OCW+cYhuRy+B8EkkJac/AnRPuQYDUCnPbWzyRv2pEu
bWrTyIU2RhsmsIO+asclgk/ZYgpLspeHFakibp4HMOJT04GXyMBFVnLqEP16Je8ihwsy6YkeOCRI
7F4XCLkheTJeMunfGp5+EH1YQI5jaL+1SNon3Zq3cPgBrDAZJEwIMwRhHCm1m1CbXrueoffDQw4s
8vMFChGdh3CEbo0e6FEQBFEYOjgyisPb1qT+iBhdANfrLQr2Su8e1fA00g6fponMVtHgn31siMx5
zvkjZREbGTEJR/gDpK5RW/NS7TO/vKgeIeLWzRcnRaIuq5JnYsqsgiq5S3X/y+6tWcaQDJJiO78p
JFWM/Pojbv89FuiMdRA6IAb2ktTNNavvj5sAZd3jki7Csai2Klesu6xAtVE9DiJkTvoSTLjMoPeQ
sGRxAtlpBKR5cRsw7qRtJm494CVbCMENU9nbeDfMom4nzRLAI7lLAE38an+/E2Wlxs/8R5hteARD
Gamfwu8FYLLsvAaTMaOBUCrTw+ptulNlxZ305nmCgwxJoCwrwzODuo9gXGJY6sujceIVobUbmk3P
4gRzcHbp96I44ENfLA8T0jVyrEYgaB59npK6YXG6F2HjDZT7mF0HO6Ypx69Q5ww8Wt/wDgt8MVyL
IJ4ALayQat4A10O9r31CRw/Nz37rwWY0OKUCduSVSAqzxljH8zJ0nDIC2tDLScWtiF4H8WDJfodR
0DDtWg1h5/tTWtaAi2U1xR3S5lyUXdX1XAmAOQl6uUh8Ex0MUC7OG3t5RpgmIVfHPjzmr/ii5Wb5
Y31BDLe1xtbl7VGcN1cEgDXpr+MelrtxgVs/ZQURua4DguekZGLHWPMnEfKYXCDVdnBKqCafXm6f
Dyl2wEZzmO1UQxXWSU8AFk5BiFRHF9myHX4aHFe0hqV2xOHbKRun9d8F0+8TydaJalRSrr3g3TdT
hxze5NWPtTGMnijZlixde7yMi/3F9G40PK6xRMzDYqP8i16AVatO87LYUOLB9eYLIe/Kku3LKZ+7
xW3PJdiaLnwfXY/6pfH1YpdiFWq3V0Q9HaAprdjFp+MYUlYQsgo1EfALqpLKjO9XDHuqeYRdwmFu
3OJzM+35gKlpOmOjL+F9sS9AmZwaHF+hWxrWtpnDvU8HcH5zlWhfDy2plvFwiFV/M27nfe8WzyUn
G4hO7mEEHgcORMh3Y2SVO3PHUsTKuwEllVFdJFDMValE/OKhvoUmLzBLuDj+rCk7s2HkKZl5sRte
avteAaZhOmTiV3zxRCUQecCGuyfTVuVE8VMLcJNl/C0aTaBs3jiiAjDgGtkKmN98CAyt1r/zvX4F
dH5B3mWIBn/0jRIBN1tnK7h/Lj0DicfrIdlN7W/tGcccgH68/cxi4KUtb1FYTj9Tasw7d4pBOqc1
K/B8Q2YGPXiBV2taeF13u/eqVy03XjL6vNRsTIvjOmORMqp8htcv83r/tABbReCzsm00lMcx1/DS
L8tumOZplEVFzqlkSETMz6QWb9oreGoCkq7i6+wvfWHPq97fTrzf7abKIhogtesnA13V5eNeZ1H0
nBYRSzMjKuAUh0/3TEN1webz6W+DLeA7Cv9txDPOFgydNql3GdyLMoomrUE3Xd7nRCGUmbGRNqZP
14IK0UmfctT8Vg/2/OIPrXzmq6qILSik11EhylVAU0RVNsaR1b1mqiXs3/WYGInguTM28xkmnblT
EUovIKqlah2ah7bkd3lMvqVmzY7lP/kmFfidKFVp6/Q2pnFn79ZKrnrbhsGFwEzht+kyOTeX0tZ8
tvHfbLxcAtrjm7HRLK5cghNDJTQEEDEVNh6GIoQplDbbtLPI3idgIpW2qTJueDhRXIeb1Alm+ZO/
YIZA/tH4H5RnUF+3Bjvx3/SN1qM3ncQ4XURo71y3qEgMkdu3k+yayMXIcPRNgfdIPsQKnNYcaFrE
zezKgDSgEJbWnslTypJsDcoK/onpDsodvJ9To8rTbD32HRdUF7FADvTG3DUtpDeCzfI5pTK88rxO
cmY328NmJIg9PbaV4kUBIgBVO7YZbmIo20+YLDOzWbEGqjVikSwI5/BDFR1YueJTfv5T+TozxZLD
5MZ90nRvHmncn2tHB5OGvFuF+70ClM4cQhTdTSUFFpWPandmQAsqMt37kZdAFqZRhZ2jsUlzB8WX
GGomDs5RxNllLpSw916ILcepCx6H3kTlBqmrnTqmorkFwriGSZ82Yrjp6LmZTWBdqmVVCKDKo8yF
2GKinsOlHzI17mGmEPHL7RjGHPA4ZK4TePJ5Erzkalotj6FXmHLbr4sPs8ss045u1pNhsKgLn+AS
ZLaQanptvCC9WbkPcJFZ2sOBCP97XCgVgJae+g8tWvRgpSKVyG7Ok8ybMoQbhTqScxORy4ofNHbv
ycqxNQnXZa6ReHXD8GcpMNVAVPhQ5M4NSKxpnv4Bm2VilHaRlhXg9JQDlXrC4Q30GaafjpFwMXpK
3oaNyiRPQahI104F3N7f0nREJd734xTUHJ/xELM6otJfO4SNgSCUPvXo6XAbPc0lfwH1+zTK8KOu
qkojD/jJ2HOymo418Y6tGiujW1buBLEtGC9T5mG8+nh9Z2uauutPHDRag4ts86Io0aetz/veIKQq
dc9IVD5pe3qaOcpavahorNH1g0M9wOFiNcW0DCs4I+KLYkcW5b7YqIGoGqZpFe931U3/qBTWekId
5Ej9VcUe3nhaAG9CcB0+qn/nKO1syx72CmUL7PAO+dShxhGAVhDMZ7I016gxXGyDJ6nJ04zKh/U6
6f3+BvAiFiwYJxYm/8GauMCZbZGuSJE9Cju0vbLiO//RJEXjloGLLr/u/jMv1Q63IKBWGRFUIpIh
F2yXBGwU/dFQs/kj6TBPS6PNlbiC+Ec1XzGp6gFNey0qkuw/sZTZfbTFAW/c2qiFkWuez3cNHxOa
RNPxcmj+LHnZ3+t+zeHUfemF0z+stAS79tohZ3d8YQrBRf02puJrmHyEY9xNN9K42BWgAh3ik6Kv
FFo4ieKTU6Ef/jjI6sCgvLvPLDi8xekR9opvX1cK76pA7+yt9DHQsbSXXE6YAZZ6uYsrig3s6Cru
dEgHIDMFnNItbaefKTGovMJki4Rbm4hun7zWYNv51DOkFhcJOiE3ZuzT9FqLGlywTukTL+cQT+Ar
FZmDbvrYygLHkL/oN0RTwqA8W7KTwxCkl/f/+K/SLwpkRisz1nWEUkckuINPxCUqXHuZ0fgerpPj
cyy1oLd9RSKmmcz6FwJebD5SGE0SnLlOxYYbpnp0A0mKYjeqV9U4eD//lTAZyKoJ7UH8vyMWBWRD
u4PVIxTqTgIOMqFZbtBy8tyFhEIOn98ff986Q8qSLJLwpW6+hshgPJuSSInScKKkb6YK6SjCpi9x
k7G1Do5AkYBYQpu7mJ5piX7P2XEajeECi6y+0VV9nXUm+f1jmqFID6/LDf3705r211awmN08graV
Tz1SLNMmQoDlC71dxDFyMs8JBcBH797oW+FsYv5nJtjCFwlEmYBuR+e34iPweNxjIjJL2maBPkdt
DYorzqkNoKV/ybWN34wGhK3JAoNiuwbgVJKlxElSXKbgAgbhrwJVw6I7vQ1eNczRW7BPFd1vGIxd
6dgE7MwpHps88j5Gjh4+3qyJ2NK/ZavZhjvu8aFItyGaonCtUG/Z8s9v/HU14CFJT591+WyK4J9G
OmBqny2oBjOMr/YtT19yfFsV8ZBHzNCaVpao5nTyb+J5zYNxnQJQvOdzcWU767zqqDrzYS6vDO6j
FzSQ+ilNLjnMUrOm6tbHXoyshncfVhljpZHm5SnTVFDLHgJ3Y/MWgDUYEURU/Ioh30SU02MCa9fX
zZrgetfnupxNPMMkq1f/dm9VMCygKKILLru1mQr1ywbyg7EXkON1JKH9we/XWDZtrlkwASNd50X+
nk63iazIJRXL0cfuwTgyt82IRndwPgWiUyqCiOwknqZZEbhMASSn/pk+uL7yllk9YfpuJytfLtoc
9OIVF5o/mI5ibJ3BeYGJgTK/5raUkdhGHLPYvPKkQ3lCdDKl64teiHGafax1MqlkSZw0XvZdF7ND
5P+kyj4tDN6OtEFF2VvYiJz/mGrs4FKXzoRiN+M5RV/OkRohC1Il6uWXPDh+H6zCyJohuZea7XyK
DqZQMzbjZNVct34oExYQ4e719ZJmC9I+wo9XDYJ5WKquXnmLLnMMmjEMd7j+Pw+hTX5o8/W/DIZj
XsOZNOGkA5cVOoMPXpUpOhP5d7t0aCY0RYagwLm13cTR85Ma1CzxXvd5icsCgrdktpxKj5U0MV43
AOav3X4shS2WN7/CVvuC/QRUhTxAqyxHOagrU7JVl6wH8kzRoaq91ErWtjMUaZWrMMDX1JYiCUK7
JVE9bOVwzFUDgY8YbCusBI97kM4Ao54ct+imgKqrsNLkkkoWNwszDGfHeKhe11NUKTqV2pe4ISy0
ymmTchDCKQk4eSsuUi4CQDJHUXSIBkXfQ6GOEXxnqso9yn7ioLfL5udbxuCD25oCanYWc0PENF0l
J1GbpQl25drWsyq/psW/MnBCTeIzC9kdR3tUeJIlXMjNxtsLpSekip29psdmP/GZzQWO1jFXIMTL
hRLUBRXLXHzkwY+ohRDvPXMOz1xSzKOJVhH7mjzGYqzivxvzGo0UOmjA9xTsTtX2Pm7qAcQMAIl2
aLx0FKMGpFxkQwSQmQzLqAKaNOByDY4D229V3yo/IHYEu8DTh4f54k7hJmDDJ3nfCkjPrc0cNyBS
t1BwOjEAZ5eRy0xw4qdhf3SrE3IvwZOPCUcV6Fx9+4zLcR3+dm/l1vB/FjoAsByPjqgDE7synoFE
NIcelOHwm0vpGSW13/QH28N72NMcx40781a10RWHenYd5KoGfJB+I97lxVLWQoZobq23sTu5fYRX
wuU7auSUWT+6QkwTw2iaZn8wWnmL2bjez/vwV4OBdMKA6eC7HcbiY3yFEK0HhXzqzVI9xrb8q4q1
LT0Jx9S5R079FDGFlWQZs6MzoQEnlWUuWDBUoI9qjDcLy5gTYqhgd8vplkQgyLB4FampAYMH/k/o
Vkpma4bD0nnEvU43G/J2qI6Td/YNXZEybulTakGg/ncKLrROqj0r0PjkwlcRN3XH7Nc8EpMXPSDv
Wh8TM593/Wwd+azFerbSmfhZKwdljGKl/o3WR11JYTW9o3fy8GrYl4F1D+eNLd8gDTH2KyrJIFVK
9IEU+67yGjPUlDYZaoZD69To7M8G7HNqbje3Ih37whTvBb3w9PIgxsNuR3l5TIqr1wHKjX7jqmbx
kwj5li5AzgdZHa3RoBBiAEl1BNrzxMJtBIA0WtcKmk8PxzrtyDRTNlnscor4MVN6hSGc5U9FD924
ZubxiCKN2uWq5rVSuAgdzRpwhrmanLUE0fzR0jcpLxCyGh7vQs0lDp8FKD2dQwk6N1MrvjsdHMGn
vghFp0RSgOJB0hHGnFVhGn1wrC99Szqw0ae9Pe1AnmmCtcl5KmYrnzkiY5526YHM0i00WIN8qada
UesS7hv3kQi8bu9DFHp+dbvsTvbXAtPvfFpR+OXbUEZh/RuJLr6LwWrjL8AKfva8mONunm2F7g3H
ZZxIKqZ1DlkrZWsYecOvmJmLFId2QOUUzqWn4LaoEom7I7N4Twryq7cXkQqc7V7ifOv/IQLSy6ut
DjGIqOMzi66YXFQKaoYe6u9QbT9XtbViXtAUxz1KfZXgfvsJHwXgkfgd4FY1C3fBh8/Weqtp06W9
av/7FZfVoUUnHHo+B57irkijb1wBTCV55n9pd3sBYPxlSd4cdf0e+hrvCHD4u6rXKJG4JNNvr4No
3o46GKtOad+oLEzJ2Tosay9hWdH1AViAf2xdBjRTuZ4G7b6LnBD5rgOm181ZQxBUECzxu79nVqw0
c9rJRSFL1EPjHS5ahLTkVNzitDEqOvLAfSCPRrsdt3NmixSLMPK3nqdUxqAYjlbc1BIubm7nelwb
hn+lcvEfvuMwHr36XwYii4UT+m1GFbM3OW2sVujgyAfP7w9cSH7CaeNXH4F8L6eTLf7R+InUUDnP
odJ9s8weAZiwj43HeTNJMh3shPkJS3/RkCR58wYjLsMQ3eBTPDtuwyVcOsvvLYuSPfBIPYFav3Wp
46J+bHqD1ZpGv/tiPz5uWH56pHu0TEzSM54Xj56LoknVtsfJJuJ1SfCXKK1oO4conbfEuPIYFHoS
023tS3so217HMy4QnUkRvf1obNgFWY1WluY/1yBtW6pMjtOyWXbyNpEbJTfZuGao3bFSB0YKSjGN
rC2+ssODQWxsgBS2WWu3Jabdj8+p2EXs0x2zH7R9/NO6ulYmCtQ+KY8vWquuJ2+iUfeKa93pQZ91
TMnvQEzQhLQ2sg3Y6HfCoOIwnLJLICZBSmMzKK0JnWIDheRevM4wQAfSUcIy5gkx+OxL8Cr+tUXn
W0dM+VQaJY9qh/yyPJXkZA7bF2gTOnRrmIVTSXme4EnEj1KPFHVAuT4guW58aRG4Sr+jF8EJUrB6
4pSerQAz67d+kJCrkIzmIDpyMJHIwiqGg1yBiZK1ZZTAQ+c9llbXNoqf4+V8tOBOtgmqnpaJfBgM
j6hMa1+46PkrKZHtfEuvvMx7200VEbBeZap2HffwbbFuQ5938vXUx1oTfl3nD065Anpq3S+SjxtH
gUbAanGe0LCbMv02o5eKImpOf9KelEIse8wdweNtbZ1CllHzegblURJ3if1qJgeICkS48gacoZNY
vDTYlxm+gNtrRIRAhc0fFzQILhQMbzLAfrCFBu1EZN/nUXyURMm6Ex4VIMLLKls4bAX9UXv8CGur
6rsKkhPZQkU4U08xCaEzl0v0ENFEwoypBRCgCq0BtqC/SWwTo1ChxNemHw/iFwnok9o57EXKAE/4
NTwxy08aqF104nOeyjr/hhrzb+BlcjT9GQhk9giv4vFWoBbMmKECdXO1wGQqOPC4Os7YzcNN3Qen
qsXYFXi009dlEsk8ycIu9weLFHjDjMnM3WrtG1vEewKuIOSQBzlcxgY4ntcBCl+xTcBbCOf7V9qB
FQDJSM5DsKuBiKiY6H6Nc9wbkcYJv8UkFJnD6xMT8kCr9wq5hOtqe18sWQgGW/vAXCbhYHNF5OLo
4eLwVGXGAMp3+D68pa7BcZJOy418+h6Fi6lYyQ8blLK9PliWQ7hokG+SnmYBXgN6ySc7LYDTT6GR
IprVjjMhTyf/dYeOUnJ+8AfVibWS1MIh8wuvx/DxC4MQGNf1x35o1Wb6uQHpA1AY8AKP3tCMfv66
HajmHq07Mjr2lSdfC4Um5cFJaLAWIAom4xvQFhLOO1S6DFRbn3s2eSiQcXlhNkZYuXKWiXsELwz5
Dluy4WWIFKDakwnfH49BQDLOC6aAoPbsIobDzXfEqTTH4Qof6jWSLXBH+W/0g0dcglKzT5aRS+Fm
Ti7pcNFBWY3iH6Ssb45eIwtD3rqIVC2nOGVXkaN1cy4b1ET+hf2PKt1O3dZFMWyb9O/WbBX2Z+ne
AwTrfTfOU7UMmPtvZejMc0ko0Czfx6duaJeli/+RaygyTHChoAgQ3G+8ZWuhSp26K6BY2Bvi70xu
bARm/Fl/5DsPzMyDajWJNiCvr+6ai6iPIBtSiBMjxAV5Bean43OaGbyM43nmijpdUFL5LDRFnki6
GOQX2s1LZaO6EH9ZQUUGgJqgMf6tul3UiLoFiUMGzpkam/DUXT36Jm/Vt4qiu07xnYETAIG00kE5
OFHPCXenZ7q0X51mRUJicEFhnpkvqQQ75X8jdk0KHNBe0oge4snXna3f7cO5chIC6gGeP93+6Y+W
+xlVd/JR/GexCYR8CFSZU6zamKUqUj6qmCzJyB+25ehMT07iOZdrZkrAYGsCLEhdwXCeJPDYybGq
f18U2n6dVgfZb9ui1uTYlp9UG4ip1jpqmS5wXasP1zcaPz12538fHN2CTyO3DeA7seu+pfXvmhYi
Y6Fo+JRdhKKr0Lp2u1YXcmcS6g7FSilPB7wXE/izxfvi8/TGBlCWirEqZEAT1HfAHjLJlDs/dd6/
+uN7JCGeCU8RppJY0JEwZrl8SZIGbGUoSgjns6n0tEiI6MPbkxC9UE6ssXu3aZ+AK/3d5lIALqaI
zzWC6kAObRb830MzeuF27h/bxyrrrMWmUuh8VxQY01sy76o6fidLZd0Q9MsB9r2qPXP7fORAb+GI
+Qg3rKBHQ1LrcCSQhybwKREKGHmnabD1/OSpIj09Ku1zSvoGbnShYW/33C8R0X5Mp5YH2hCvneex
4UxZAJfTQfQ8Drur37ajN+K5IKkwghPziAFcJZD1/nyiS5sjPWO6XLWvXc3+mBBsYR44ZRyxFaaZ
/Ntrm6zowt2rFYWSlONTJmJ/RphcQjsVWUMHyq3efOL0wILCuwkXiYyKLNlW6Ps9R16AcAOxtf/4
TjJyzhaOps8fCpthcaBwbNyvu1C7vc22hJu/8nJrQd/nuPNCsLTll0PcKqhwFcTkd6vLFhunnYB/
djP2Mnc1iJWUx/mBkULVLvxrguHqdHegmglHSm//pWx9DAkQNvYr5ZBG478Yq/NLUn65PUdPEqJl
JOOt9NNsUJtzj4nYJUCOvRKS0z0XK/ILhLRnD/mKlGbugw4ZK8VCcdDhoHylFCqeWAZqaSHPMYhN
/HJedz8AbjlaZxc96yeEY177M5lwbe+mrkdGY8SqX5tTP9k+34+5L4tQT/o9KkX1vufLXXIdVC39
igg0LogzmS9QkQew8N1/+u/lGazplPRAcAiczOdxTSYTkNoEVPwU6zjp/LdEw5Iuxu9UDEpGObYo
iRnw1Qe1pv/Gj7wyLkDX6EniYw5lsGsQ+ZcRLQNhINT0tlP3/SzuP+IlIE//aIxG7Vj7b7IKOnYr
Cnd6y2lXDG8HRdCz2HUwsHB4XKKrt/3UZOH/mt1Ltlq9836GTo59rEi9sZJruLQgZfnakdor4uiy
91pdVFz2mf0WIZYWgP6fVa3HKxuM66F4AaP2HE4Qt69Wv5Er4HXqeMaKxM6zPWis8o9xMfszeGc7
2Bfde9NWx0VxCsfNil6lRDu9d39khcddPyeDQ/XXAXJpnJQhnvUkbzLnnlyoR0a1ejpXVUjUQuy8
ZFINOjHAfvWg3UX9icsxwF2XKRZld5OCU9UNLqr53S3TZBaRQiIuThKzENfQo7Qq9RdUBRSPoZhR
z3hi+oNlUT4YWJRqGZ9+nATWumAUCkgcJlHhuY6TSgFkbGt5CG8veOdyPMGB+ueLBt2/YTMK1Mz6
UmPnxzq40h3Qn8lgmN+5duJyaunoGxZEZoxjE7bG7T6GwkfolGeauFNlyO7dsLfDkUc1/1Z/VkF9
Qh6Sk77Fd8pouXHzFnyozKavrR2+6uw4jXCfcNAwvxPGtxfEBTEx3M1t6CYErfk0DDrauBd5qf8E
+oq62vtMGjtiq0x5AEgRoVm5crBkMXIhK6s4WGYzDDMLjtjUYLe4Sgy1bAduLfU/jFJ4OZ0hXmRj
pPuqMM4f8Hnebb19Df95dHVjasGJuVb034wfNwMd948NunzM7fvsLFs+dswR92d++ot3u+GvyPWQ
AQy3MO11YwTSI0NUkXkQb7CHmdK0o5hbafL4h02ae0Ki8ryuR8lFOdz38CXWjZEXPfg4doF6HOQB
6w5+Cg8z84S8R0obgGEHOZHRL7bFl6mSmYaFNnepuNqJrvT/Pe3RMD5mK4OvD86ABP9R/dnol136
t4Gec3bOKd5E2rISyMw6YivvjExcm1p9ecpIIFT+l+lTHqhimUZ8EZYj6kK4OR0nkPgG7Lthxy1G
o7YADtsTY7HMxOAS3TfsZ+okeQK9jviShBnrQyzXnmb+D6uJ0VWsJcdHc0lT6btP5FL4Dhk3BYcO
9VTDzyRNReITi9rpqq+alP269Ahiv2e0oQFTB5qZ9nJse0BVDtdcNCcUj5L0UXBlV9Quy+ATKthf
2A6o86rcz9P3icC9Z60bfP3BEIaZABmPvea2s74PNcx3RMA5gdSTyHNx8Vt5PickIBhi+c5yb0AH
kYYEaR8Gin9jWFuTRmbobgsZ6lAIWAMswMIUV+5Og9TYJwwcmAZQt/4bL4tMiSbDTZ1adIqy6UK/
xJnhB15m7rZTGAe0aa7ZaXQcaIr37SLysDfRUjMW5LoRFcQzUXus9oqBDdZ5D0+G7OC2ekppdMmp
l5SNoRMjRYi5BmSsDtN4cLzdcaY5gH08hqrmft6xsKHw466BCu4vH6nMhKxsq26Z1wR0N9snerK0
SQkxHKCumD6MiLND2XyR2XHfzJ2ykgzYigVqgbDJBkzTGTHW8yWHFLfaS8yEZlYbov4yn7ywv3UD
sZsuRP4zUdG14qiAhb46XPge46TiqZvpHmoIlNBiqhlCDAdmqpAVh1Z7EUKANVd77qO7Wss28l0r
iL4uI8rgp86hLMdsdkiiMFNf
`protect end_protected
