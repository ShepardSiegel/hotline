`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UhG42VhKepIzN/FxXmX1WYSjnKfMexdKnDhWQiJYcNcdqCkXX8dv/DEJBMTSYHXzXUxkAU6Llmdk
HXyec2h27Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ogtL+2N1bjy75cc0I86YTiTvS2/6HKonwPm+L/vuPCD1rTFQfP2PsDhto/GAjGsPEsffV88XQkWV
GwEJqUCHpxuWf2MFqRu7nK85U/yf/Kr58trvZDyGCSCxHyDFfomxpD9YxwwJk1hz2A5iYbJ9XNa6
An1MWSIwsfmqX0BlkBw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qvGhWsDk4ZRNEsnOmNVT6bIByHTbMqTtganWvgou+6apsUT7OY/vrHXbEa8LUsr6U+KC5vwu07KV
+5mSYZxa3DW+AkROlKGdOdopv+hAb68WQ0c91zQPzXh3t60kQAkhzFSrkqfvXa0mYaLV8WtCV7LP
kntIn7z01i6c33TrhOz1aFR280T/mH2umtH/S3bZg0B++5ibxX71qndb/g+QvSlDVOva0ZBuV8e8
aQOxdKCRtqdzeKGLGYn65v6pw2iEO9VdXoHJYR8Fm+e0E3yHkry7XY3T4IsKGU/rir3DH7+w9Uzk
O4AJsfC10xPwwUo8et+ZD972YiaLje8YQt8ZqA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uZB0pf1VKcV0tQZtwunKjwhvmBLiYfL9JOSTEs/ZaWMNpY/XZHDQKcQe9acUm53UtKWXH9T2IhMY
Zq1oinAUlGspOlcZvqVXcmerOzrkCcouErrhMWYklDAo0muQpQbDY/vg8cxngwe5LzqpSnSIpP1D
KddU1BKX4xh8WB4Rm6g=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
R2fL6OA+Er/h1REzZ65WsnPfUFywqhUW2qbJBZ4ZB/dHpEEUMUBTUjVXOUePOZ9CThl0clsv60OI
6e3qzTQlbm7ZLXl7K6rUZCKg3gTz3hmi8XUZqRRL5Cl78RdbldUn+fdZ0Q21/KwiEOVAJtAYczyp
Nmw0o0S7d5oNKNrx5ilxaR3JzVwU1YNRaZ4wfeO0JOUiEviTIzidBJRu3YiXcfD4GL0Z+1RESVzZ
tDZqOphi5HzzFLwm966SAN2HjXGyMDAwj9OjNw35E53G5UnEb/emB9n414G98qkydIW/g2mV+YaK
9l4FF6p+oTvieOBPV/B4fSt02i0V8C2Ql/WnvQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 34944)
`protect data_block
jORvnvML9Al6HkSDf9ASlZByS756JOHnGw1c+MSWbaa+RiSqy3rfmHbBG8fTnoeP9S9oEzzx1RmN
83Pfmn0GVXtzArwzFgiwUkbD3bJO5Cg+LcCj11imR+IJwJt5N0Kuytl8bh66IM5QSQMyUhswSJJ3
KwXrawhCdilx9zJeeQ0jg/VhVsb9Yz8gCi4olBBkxbtcxPQXPeAkhH4yWRYuktKoUPD3sLQKjAtz
FGwj+xhdNVnpNNZD2fH7TO3u459IctAD5HI0C1qKA2mo0AZpUYqfTYW1SdEEoucvP8IP9+KO8N4u
gAfz6Enqze/AiDjixq2HoaUuBcAc9ocK9FPZXWxRtRSOOoK7HFiaybF5HyaM/eaBOTjdg6pZ/NrX
9GE6EDL9ncCiQqRqQao6TzYg5aSI9QHsaLfMEYUn6y20KcdvsDy6LIwHhKR9oVzk9sbIiVSU8kGp
OlOVvX7RbnHHn7S1elBvI+DK+P0I38O0xtkkOqgWKT6SBEvvV8xSnQnssbbX5sMTXuXq81MMmmPM
EtAI5mDVcjKLubuAZMtNKlbURm9ZATfhRhMVsk3rET/M4Gd/LZch3wvcY/1Phf/nBsFljSRReZWn
ziXqyInd993MUQ6p2L8d4ccUGUH7KII33XYGGfXQOPq+MADTQrItTjBzGVWNKj7T4Gcli1rAiklY
IYje2uS8+f5k88zrYZdAaCIp/Q7jTOtN60kLRmTJuFiV0ACl7vaDaHaucZXn68JJxD48lF5ie8/i
xeQ1ntW1pX2tcnxngk2wGTUoE4Om88ucMum26ZLZavl9UO1RYrc796biRprWACe5KW1ajnlECfFB
sD41B/BFMamw/9m0pp49ayb8c7btHVm8h3K6WnAv8JzCx5UYyavcdYqVT4/A0nJa5V0ZWxEJeQPg
iWDNWrDhpvPy2emBFXKLWJSn27cHN3wSLOWFfZCcnTx4wafbySAty524gWj+ed6yyab1XEp0Yh+f
tilN91hcfsFH4qAo4sfr2gCf5xy63UL9QVF5lj+vkUuLEtN0efdsu1lppSwCuQASk4RrzbTNn5dt
rxv3xNVOSlQJw023vFp+qrOcW8l7P0dd1M+w++dYuEoapYCZ2NPpIVKb/DzRpLEPtJrexSVSHWus
jRtt6ITKv9NCFRbFzTwp0gZmxiX+ExCNkHcPZ0BgrIDS+wlk/gHt0FhCmJCcz+/Fjef9HCXWM4W7
NyJ8iGNG7yNW8Ga3hLf+TN8TYA8/JYxkzduiI+ZBnqY1bLnbs9/sFah8jDAQU6pHv0rQ5EmjuMFG
t41bV+qN3rftp3zFHGmD+cOgZFjtS0u36rixPW3KfV4kSs3kJVq29ZXtoLpwavosbQ0pyd44EGxl
oPXMes14qQ6h1JfiY6BkoryaEQxrlHsDiOg8dTqpmCV7HotqiPP6hciwcSqXh1DfH1tah2aoFV4Q
jKb7gZ59lf2VD1AYivLMi3zVOJL4inacB9U5to6VtBejqrEaXkP8QqsFJFOQdgW41MrADLlCQH0L
BHSFkmTjzjkJgyZ54uC/Yt3xmpLwgew9Cf+hVUOW60WJTc/rgZaF67IV+4w9XxstMn4yDDHdHBSj
GZF8K3/qYjjqf8seRND7EvAGSWIFFnBEJuNow5rBMHIvtRbzkZbif81yDgRHu/pkkmLHt8PkMcSB
Opq7BoZxFhikMQqeffzxzeA9b1oyiouA/C3qEQNh0ZYvuARUA3PLnV6mAigl7/dGVuZ1xtfHFZEn
MKNSqqkZKTHBZgM8sk2FggrgYZIOaGqYvUuvh09M0NJJF4phU7HxEsAPLHn0USuoF1MhD9YBtTU5
1l67lNlM/gYX5u4ZKWXBA82tzhivnFqDMxSHTPta9JCr5cyP7bnQFkFb0VcORxhuGhWt/hLAZPyJ
A13Vgs1LyYE9F2yOSHX7VQ+N+Jy+Tzp0ANECaFTbpbwdCNHVZVgMNyKBZeajjGqOeb40skbAOC5e
MwXc0gDvmUS2T8rrw18kT/TUX8P0xUlM+Te2rSkH8Ch1JguRbpVuWQGECBS99/x1UVhM+u5RBz6F
WqC/NLl4qnU+VC5ENxVTU4zNP9/nS2Pt8eKAh54ZPhlF1C6daqZaRiE/+qvp3fO35VptIdyOW8J6
Hoc2jZvg43AlzJBooFZqXzUPVCvKubZjlFMuHrginXidzcO1MoHHWUc4/mhyaBqXqQ38QoS/W0C5
3xaNkXNDu9jb7EdEJpIEtqQtI2B9ydc8yB/fF3Rx7ySJpzn4/nbPhAp4FUF/XNxStvXcFLwWzdNY
dnGjBU6/AS4sSQKqPoElK45SQLN1j3nGZqtvx1pRR4yNUX4Hj0WnxXrWTYOaTkBPVyxotzMhD9Xz
IrWoXe/ePwUJCA/PCQcT8qJ1kVwgf4IJvWn+OSfj4woX2D3mxuG/k/nyV3AQJyyEEankNMDdee0x
QVCa3Shc1f8Xz2XlShKuKEMOVcOmHxNB/XdfaVOEkAdvmgNb+yj3pgzD9faXSHDUBRf/03kKiLzE
2+Gq8EVqxw+z+n8UWZYjS2AJ8ZUPyE3QodXeR3T9vOD+Vn+qrIbCvLqkEkWShjTDlH434Of+VVW6
XEMAuAaylegiDtSKFVLKKlIPFoFD/D5cuWLd+Edrx/HiQP++kSzGYesMf1UJq5HB42iT1cjHjumF
y3mkKNTmXaNSxxVENDekJiVDJpOqrrnMp9+w3qdD19mMZilnKto/dVrHRK5SZTEkL82bD/SzZ7wi
0FwMKExi6bX96DkxxwEURbb5+kWCwKUY5DviiIxEhFRlqUr2RlPwPb+O1tKPFtrND8G4WY15PuYO
WbFVFuRNOvSil+EVkSHBRTR9robotey8o1OqErAw9mkvijZeVzCAlGwA7nIh1hDa7yU9+CUHFZne
TsJrErJ4BS7wB0geXYWaMJTcieZHO2NWfWFjWV/QCMK0r8nc9zg3PlycUm+pM/M9od1G+R8yNSS7
Ld6dZd58F5eWEFQ+V+368DXt/iMNKMlLdppqWEXVWS4LKkMDt5fJKbDiwZH5VfMjEgTHB0PSK292
8T5+omkiowk3JOjR26TxKklLcKtshJq0DEpx7Wvk9IY4gemZvj/NIVUKYXHqq/gZEP6RTrIpO5vS
CekA3Qkc+x/6dAlB+PBKzRHI6Vo/5tEnJ3OLSu/INOAqRZaIg7wAbqetTYn8CiUvFZToYFktMTJ7
cc0IK10PLEdlo0Gvq12f3oXFUt1h650nPILxrC0BxcuoZuu7SuPEEb3I7HUne51Dd6p0yDog8Dxs
xuvY8duvb91ZFZQIh/ZLsMzNbEr7QhzDw1ZbcwSX+zBEhlk4D1NbmKFSMqnwvgrjkQLHAK7zUUUR
FyoTVMycKV7Nb9NaICLAirA1GRMO+tiLsnDviqTbNrRfYsQNgj0M36HKK12a+7Eirgpkbg+WLCow
iOHPCVKLIep6rD6RTxyd7N8lQia7B4DvTvin90gVRm0crApONNHfn9R/G8uWpWizv4e4kChHocmq
68xP7Veet86Ys5cU19n5sm4rtX+7+4YS2MFh9zvO/Nf56p81Ne1YSwcnn96PXPMqhHKacGN2zcKE
8FPrhTo8bNthmZaMDUYlPmHdchXQ1yjmaxDbtYYJr+B2GMs+S8V9OBQ2SVW1AsmGbw99TRE4dhrs
vcAZc3+F2ajJFgbIU8BKjYDpzziDSCuPKJsyM8a72VCVdj7ltzxXY/yMUstNO3ZPaNoWcCwmVmiT
JtxqOXbB2tVnl4t3vAooqUReFz5Fmz+fGS2jRQrix8fiwptYDdqES76o72hlz0iU/DerTJk2+9W0
dxrNAXYlgNR4mzGVhD+Oi35Eu+KDDUZniZJM+BqQCa0lu7kettpneJ6lhAUH5Q/W2twP2FiQvxPa
Nlkk0Wac4hJz/b+BqUtS8AADmlDuBXqKdvZkUdLhYBFdNdKMnwIW7bMXL3oqR8NNV8JV7xuaqDJR
a1zNtp/WcUmdLmyw2vShI2b2jyju8jCT2TJEdvQKMkln6g9t0/h08DYruRel1BtIZA8dxcre6jCo
Q3qatpVx4DtQbdu27a8AIfjiyox3ojzeBqgCWvELHkO7hHuq3WwA5HHyNAQ06D2MGJmpMOyAPYmT
U5eBfEE7Icd1V4NVjid7X1ik7T6ih1P06Pd9lon1VAhgd5LGgEcw2pauDpB2/93C2rKeFu1o8C7C
DyzXHOKoRO6NkbGxkD8AzoMnmcnnezx6ocmDEfbb6ghcLkvnxrDe33IPKsJ3qpl0m1JbgmHWB3hE
XfxhKHHIgMuVoDSBo6kTME5cP2Dxl2paQ+RJIGf1/RDRRW1iRE1W97rH9R+e9OxqaojtxKBIgCzL
pz5pBpQ6+3q27Qdy3vCdN9bhDZiwTWRaqRrPVyr9RD+Ax4A/lwAp6W9UdZ35cvmYRgntcGjhSurD
iGSdBUgspSmKqutBcwfBlwBnS0CAXfOLUZRxwZncGbFsUozBoGZkvNb4JInQiLg/da6xOnjgJLm+
Xackg8/F7tkAEjoMGv/gdDiOvzfxVlsdgIOxD5WONhKxmZ2sJ+Jc7F8JdNjRUl83yfFSXYqxHPVt
Gdi34iaWO+7Jy/nGKUs/kDW0o2iukPiiecTvwjw7MPZHnk22X/2Sd77ziPaCNSA15PYZGC79xQ7r
yXoF76Jp2NQ8ix0OKrIo6uHiZ8MKzUyTShquAVPtWlUnkuonOr3Gf4gUUshtskPDVHTYSipia2v8
2zmjFoiPXcfevDaJbfeFdSqAx5oz/e9MxPD28kLXuYuSyRFWZAq7N7f4Ivn8czRx4FC71gTbyk9D
Yxp2+KKa6dovQUGSVKTxOKCrNzCK0uOs4FsMIrOV/1WOk4CFlUWltCF2Ekf7lmKm5thhSDMZtStI
4lFPG0J7n/uI6r35J1e41OoUS5BgyfdGmEgChMeM1jytn/3CFXA0L4Tn2kTAFjc0US5VeX5XK0uz
/7Vy+Dboqlgl/3i4e+o86/2g8YrNUZV1CdSbLJGViGezFovwLVCir2cRce5jMSOasLKKfWA/3d74
hgvebVpHTqa+m1w2x/4g7NeYbe1FpAiOm6jVIId5MfPeX8yDvMxlal4yxFMPQIyRT4DlkODgL4nE
syYpapxZpW7b2fzSzUhiqkWZhcdmlGU+IQzQ5jAVI5cIbC2z2nz/DKqX4hfL5hwDjeMe+o7xoqTs
rQk/JJTU3e/ZXB6uelJnIqeOEElj0wuPE/otZ4CVUbrLqlPtbctAUASLw2IsCaHxYFZquh+5iA9z
DPs/hM+sN6PBHpneYSatuswuouyrR9ebR9KMhfzmA2eBCqewyZzPPTX1TIs2PjXUIFsu8jvus/n4
zI5EBgb+Z+pWze7pIxtNw+njwDSIGXKw1DD1J4qPlcUBOEg2/MoUk44ZJmMBg40wicZlSXie626p
xMT9tzuHYz52eNjflIhVP9+zx48lq0vWA/6fBinmkwy30gNklIFGYRXCGmpKr6EVxP+Z87Hz786m
J7pXfoBfwtEK8bX1MkYwAVtzS80wv7BbomzYZmUjOyui+KE3cEt9BFxdJOK9U3cSn+w//QHsFlfY
MvHtrdXvU+GZ5tPTPXPtXL9HghjS4eOKrw4r5v6ZXSZmW/Z1R/YnBZkNyn2MZn34ErYkye1vcpPm
BnQOmsnSGq65z1iFg0O0dsfTluXi5IqnkAHCw3sC7PDzW9kV4oEl5ABeRsTGpconEulveq0edTaU
kU+7dZbHJ2+Mvbv1pOwZXFEWNQa7Ut9evZi4rstXeVkXFDdxsHbCy8gw3bRiiMWT3z+EszGnPMd+
w6E50rjM0cAtfud0f65FEA9+036hFnWgIgVXrTPIgk+03kABr6l2yj7PYN0U6K0zFdRYnrJzg3U8
DuaJ7ajgrdZcjRhkXEJUku9lovYrCR2VTjeVjf9+kWS0nV549ubO9RtsLzFfO7UkD80qZPB+CMRf
R/fphtD0oo7BdgRFXRPQEJbGE147GhBzfo0zFsWaahFCeh6qCv9sjsLBWvyeCDwiUkkw4LkddUAA
c9/eqW2CGDdxp4rXe2JTLrHD0kESa46SJt8v1lLkJfwdrxKT/vIovEbC9kyfRkq3Xy+N/1YiJyE6
JcQhwq8OBkUQvmwLxoYyiWSWENaKSeEI+uEB9sk7uqU58Rvvt/awVEvncQ0aY8/8CcgJnO2aGck6
5GjGn5eWBnt8r/mYXbrtuOHHTM2omdYga4eJIG+JyaI8KeCdBHGunrMnsQ5Q9igEDrRM4kJTaJBH
P1AGrY9VoxLGkE1/vN7ewkslRaRCR+6j4s+a4phrF4PgQyhMttxnb6ybLM+kCMMh7ORg4b4UmsA9
NuT4n4NNh98/QjG48+9EYiqVq6epOd9l0zlvk6w4ALslVunvav/x/dd77KqL9KHMejpE5EX1/AZK
/uCYPMDiJmqQ8947w6XbWBQKUUTbvsj4QUxVIqu9YKHYXKt+9w6Avmp5CYlTjyjLGIp/qIrxvfqw
rNaHBo1jRQiAS+s73+wueBY6EbTG3QO2qeQ+ramN3BcRPYys8jxRkn1tnNDACKOMJjN+VcTE5IsR
Hl4zjxNlDgFZFZvF86v9k1l/8IwgGyueRtu21QhecMqba4uNOD/cZBhTrcBnWDkAtSf/SrNuKo0U
Yvc/EFaBGO9I5lt4A7dNfWjRnQoTSTspNrQ4R49WEiyNrbxRnjhOsRR4F+32sXMj5P7GsYUhg9S2
6LLwkts2SIiC3nXhmGx22+XkXLl4L4pCP4EsgTUfouUXDuNJOT/FfFAPaJri+hk8jlSkIPQ47JsL
fQRxo39vyWMjZYsxGMUTE0uCoDI8VLHDCBKT4PTuUGMJ12cQUTQKbG9+9g3x7jBnGoAjXC+cucam
biXqckgyRrP5If2eHWTiLYhXVN3YHQ/Qv/VyAdf5uxD1bJrA9s/ov+NnJsaes8Ge2YFprsEksfrL
eWEvZxevDklk44MkZZSbBgH2OBgpOLwPl3W1u8Yyt2dWp0ypFjdKABxmRScucrLJb2EfkdTVMYuT
8RGDzHwTgHVKW3K7Sn3TCH00jZcru7jSfhEFF/d5t56CwpUipJOU5h50ayHkg8l5xst9H07neev3
VDwqxKHFEIDm81DeWnyyCQXfS2eIXTSw92K0JwfsbMZUob610eYHoLMNXuCyKuDQPt5g7CUZ1HB5
tg/bGPBbNJxiBzsbxXgPLwgoXllBb2GJg6PAQ4AOWdP/6Fek1pIOWtw487VnD07oSFn2xbPUGTkZ
rsd8feE+A7FsfEXLYUOtbfI0MP4v6hpu3Z7ErXnO3o8g6GrSGHx3fAxr7u0fBr0+ulGDdD5NYSoT
3sE2DpFVHGO9AcQDVMzDazbD2f9XBCzSeBuq4VrDlYDljA/2r3Dog5OYM7P7/h3eqt/mNdxLy4aE
GF3baWj83gEMNNlgolcIXpfwsXFFQxxXYvtOpDEkuKgLPYJOuVWEhe+faRv4QECnDxK5XeOOPkXn
xa6d21M5xfe/Q3Lh2l5vUMEzW71mViduFrFtb4HAW/q4akrmWxKJWecWkbpPBNzkpuHiED/J2Vi+
R9xNBrMSMFLuu9xicKU8zAJoTWWw81ORGsjWOL1CpZEI/7fZiqoNIQZ4qu938OQKQqAgFVMayF5S
TTUjkWN2aiFyu0RWbUAKhNovkY/88mTzVvJfYPHBF6WNnHpEvFHZonSvFhzKkTBy5bOOpiA2a4+j
548AiW4sFK/dI4DZ4YuNEHOuwntaVjo9Mzq4AD9IaEXUmqL2OFXLAhYQQ3mmieWSNECQkYhxJNvY
ZlllZErXN2DyNJNsOlCF9sILT3+73KUxE25WM+ufJ3dWNWHAW3R2HscZqwZFIg2HIvWsZycD27v/
kz0JFbxkn94wVoq2BRr0nGKQjuhhpEYiAH/KHRvibJeLaCmp6bZLnV0lXQPkMBKVMiP6vm7QsBqp
PtFTkOougqJKGgAKaGXYM0bxdCnoE1lPa56RAu/oq6caxcdc2GzpQoUPv0lVZ7NS1jIFDGCoOjSP
wcVlur8PnfhTbtDqDxflQ1GpZlRqUvqpfFdu7itK88BwHUGhxmlrftQPfiMtQ33isZ8ndhLNJ17U
KS3PI/4uuXl6sLUNfCtZAk0TgkY9/19vS4aYfep4hMFEfLXDU2Bl0EqARCDlyaCrUICJE3ssAT64
9WERmN6zWEDNZKQZNYsEqRI0EqePWIhpy5Vtl9LIP5niXDMtKZov8vqIk4xDxODWmjUkd4lxW4aM
xwh4mGHhJYErIiv5yWbO6gZfsRpLLM8q/cVNwb+gKcmGuPCMudfESGvefFYgCMXdh3PNgC6cHIHY
UzLI9lkt6Nd/3lf+yqgmnnbMe+4kM7k22FnKzw7fRBYtf8b+PM3/x8NizkiklgHZSiDLHGs3G1EG
a4vYkZPKU1BGGe5nf/iTRyMVilkvW2uACf9bILtN+PCIYeUXGUdWzwxcRZuCW15hzxk0cPZTr7qk
jp7K0k0WxG7DIcseN+hooAu6D9dJBPBfGapkZp6frV7ngIOnl1LdmpJqfPfmkLUOUllKvUMF7Kcg
dJqNRnXdopbAYmMeVuYRbgXj/smfXvBayIM/nEIRMSorgWwZXIX9mTjR5Pt2qR3SaGvyxYrXs63h
7njH/yEclNkY6tjB2fRqh07rUTm+T6V2ueGz2jJMfXavFRWrNiO/Ym2Y2IjSe8/olP43OKndzVXY
NUe9YYWRGhzYmeX9MYSent6vLPocMP47xltfxDdzakXloFJemxnUcTp241bW4OeUCdSmE//pKEzE
xcRkBq7m11N6uUW+mxji9lSE4NXUjIC4OBVK+wK+OlzxmyFDG2zXapsgDKSFChvVdCixIpFFLalG
zuUWonSQHK6c1Rh25tlsMvhwYCApUycaTwT4sUon7DscERIJkbhEn9i16qIK7+3lzFrF8CC4y7gd
H2ccmTDs9dTPDreIWEbbbHKWsGJY+fL/CAoMu2LTtelQMHDLyLxP6zytp/frd+xHwDHi5LbCXYh3
l5AgBM/BoU9C40oyWAlv2IAEUigfoED8oa5UF3RY4z8MnuD1mOT+UMOC/vyiugJepD69S6M4crGK
skF0kbmwXnRWcZjgEybXD9E37HVh7ndmqife3J5lkiLGVmcyVttshSP7Fb1vkBvFAcwwEeEQDf61
gizl3Tejq4XWqurv3UJAZsd/Y0PN9Zwyk3yjh0rAKgtXyzHhU7AcUjHS2nErr7B1TY5UFbFrmFUG
UxW8rKaLboEDiWmhnB53pNRLiBydHhgNIvOXcD7wNXPBB/jheEiWTjyhGbSwF2SPGbrNRvBDqYlx
7e80r3KtkMLR6IPVV25TFz2IruMcwROCH1Q5yxiPDUBUOteld7CrVEEjDRkcLg9+BLRO0xa/iOGn
kW+/FL9XUKU7AmwzMQT5616CVexvQ6/6MXaK3/1EO7BpW4PP5MeGN3uibGQ0zSkKlTYZn7rzHqEU
jgh9fKjwJNZvEpv1igOwE27xRQNZYpYb3n4fiZ6QJvegz4KOgUFCFffCf9+3j9bZ92Rfz5vkSKf/
oRR68I9y9gEegNU/WXXQCSXywHPxP4uwhDmW/MlQWE3Xuy8W7K0wOdGziAUGbwEpmfQQjTOFMwSt
kwod0TR093IeVDhyee/Y6VxpC8f3OEWLYE6gYO54fU9Hyf42Mxn5mqPHZqWy3vcqXJrfNPcJ7foa
UzkR5oa7ujXLdkRvFUcW6jdkS4MBKdYTXA68mLk2obZ6/3Sy1pCiqTAjgrikB8yp8EHcX7wqut5N
7nXTnRzU+tNAWvtr5MzCLwzvNoA8mECCselHZzdWsquVDo5HODtyHjvxLLWckhKTDnWaMBmbzpJn
jDyoAbo9oOmKST9EYRHfTGG19ANBHRb5ofYmzIZh9KPn2Gs/ZZnwfpA/GIjUmgL0NPzGOWPtXhPe
i5f8F/ODKgX2MlIVY2apu2bD4z2E7qafk+h+Jz1BuvGihEZIxwQ0dGbaLB3VCRlKoxf9gQeRZorb
cZOtKgx7VHxWd3oYRr4toFDqyq0LLgeFUKqwnxZYaBORYeywmfU0mSh6Bz0hz0jCx4m9UTvxOUyz
8+JlVSoQanDXzGVMpDUBBwwQLXAsUDt9j+ca13TL0P3jYdR3JWgVb8bMXtb1v+a/EAFRjkIRL9Vb
0Zzg7VFmmPR29oCq2lhU7nxstrulLjVbpE0GqqR1lHkh/ebnPlyoJEa+tOkTM29NpvL0xv0yRFsP
s8a7g9oH0/Sk7x25LTa3Iy27jsgaXbU7Oi3uS85nkSjaDGBg81J9fUMmPY2fdEMQmWmR4J5lh1py
vtjLcBRbRC13JnxND4rC5tybreDBEs09lR8lzARV+W+FIUFaz9gWzrg6Qe9cNBEr+bUAkSD+CI60
G3F/LGb7PKTDKesPw0/cllmfzjtBMl5kL0zMJulXrCZXzLdj0iC1kq7l/rGR+3f5hZr1cIb7F5DO
q5MBiQG6+JrDwbMMYVQbWkv6OZy1SDlaw94Eip7KRs6q3LIW4azf1FZPac4wjRrW+MGrC+7eW867
ZMKhgQTPLGN5exYxoaHHZ/JtzUcRGyv8wkFxiNair8IiNWFm9SINcxfaKo2GoEkjMsnKTSYBbKau
XXx1pdp8EqjM2FjnMEGWQLbeRdVKvuWoqH7EsElg4E+btqmprtDssPALI8Dd6IKmC9HeN2XFhWoc
5ZD7d1S2nB2iEq5e+8UBoVV2XmuhQmtM2Bddl7zMa+moa3yYZmm6S8knkcJRTmhrCJ0oXiORg0px
sW+EJ/Me3V0QlcNyZf21ATw3YVd8M8cnRHx977dnUM/2gK+yJ+wpb8Wm+aZ7TjLV/hlgCJIbbnTA
Ai3bpQR/22R5uHnAqAdVKaVylDDfDWWvNVnGKBmCLmUA+6uScv7WrxTTfxtdlSGJEeIfx3RG4zr8
XINyRuW8KoB3DHLDc/Rg5FD2PGLcZDKPjlx9mrVziftyOBM0DiyEmKbChQw0pyG3+muF2gUb05ZS
IaDpHtb046BWWYI6CfTKARDqNIGHU4EBeXYdrgaFDUKFkdYMXuzMLZCEfU6zasdMD9x7TzvWcCul
qHbQIGmzrJwV4DJrfIkjJjFtNkkcYqTjSdenqUPU5Ua3gWzxbvUgnzv1Gvp04ALL5U+pH69x2dqn
17gcR9wCVJT+s7/2AxAkyO6FNo4EdA1xA/Vw8X8dbcXLXDfQN+pCpjlJaEDFDpklpIlFaSGbYnIk
ocl9QtHWwrYcXu+pk0yQS+RYSmiLeT+2KdcH22fH0RLXIx2N5Grb6kBE4QcGRBSIbY9CIt8rx/0q
m0gyZEocId6NFsv2nUG45gF+W1At1EwxRwzeK4AG9SVnz1tV0u1iwBuQ3BZc9vsgD1PJeZ7m4/2S
9hQPxW8+28qZtSEvtX0BemN6Fl9pEvXNHVObKNwj3AgNkDVJOty15CdukvLHww36cOP40KXnRzqz
UJW8bKv+PcXN10ZtG45g5dbYPGcVMfS7pEc50PG5q4461nzTKhVVTD9xaABv8NXVP4LcKj4g46V6
twcOqxUcC7XMe++UQODynsTVDcbUsxgyJh+TmVyaSxjLyxohCkYjIlcBv+YaBlHJrogPvmIU3pPd
rhcFemHYGPFQeN7DvCx5UDt6WxJQeRjpBP2NBRZDEhM21tI7wn9smMYuEdw3er3lB3gHqPTnyIv6
4wd2bJRfieol43csEesnUECOmTqAuSnBc2X4WakRkR+V6dCLI1emd3dTehPQzN+Clbz0UPU9y+Rg
NZry45q5hg2HfZ4MbsDweYDyWQWlmhrAQL+MEIf7onWxkfyLUN7vGyYssg68g+P4s82+9oQnx0yv
zUckN3ZZ4z/j1cmHKtMFc+LbsAvCw5EhSMfx2u03SBjnpo4lZM38z/Eh+CEO572ucCrQY9vfFavK
bQHJrOb0snxNv0ABxFAD5GGEwRF6qjosqIZoVwMogiroUg7LILe/lllL+CNzhaEZGwZld3J34zOj
W/NIE7pa4PD68YkKekNNNL7Rmjjy4yzlkZ7B61tSmWHQHNKS8LuxMjCqcMymTbINm4lpuuu1sL7B
xWV/ErJbBSPIo4c6fXdddTcSSI0jRM0s784ROdaxnO5O0xPwK63H430u1wurlgmg0Qfihktuf6m4
qXq1BydvvwZFYFyKwATVyz3pmLfSumm16SQD4cZ9MPcHffyV+6KZOeKOYsoTXquSqFvT0dU4Jr3U
9GoAQ3Lgd6ukDO9nSUj7zMeoyBhO2P7Dcn8leGX8SzW68xnEZpvdO4jWTaZLc5J6vLdF30Q8sXXG
tS0xfcFrcScFO1W5i8PTWDwDLsvZH1VBWtwcLc+UtAvf9Z+Ku+i5SSdT/9FwII5es1v593ZzGCVV
d78nY7n1ZVTEZBxjaxEzUy8i+aWI+nWuBkOuK71ixZfbQq8i4muhe8IL6HiYUaUAZvTOy1f/PeBm
b84O4/JYF9ujqcThgdydR75UMrb8Q4Txrka2RMiHBbvSZTl3VFdet8t+HGgF8ujChRQri42lZOTo
J7sAQ+8EJp5E+DyxzgBJdbnwdOqup7Y3w4Ty0l0Bue0ccHnkWoF7La6aNd6+cd5xedWRHlflr99z
e+X6OnIEJl8hQbhOHbDWa30A5DHPd/dO2MPAGn0CdPMjBOiL0sCa529sdowMRTjVdTJXa2ihXfER
8VqXiYXLB7xEz51hCPuo1iWoQaDlytciCZuBMArueFzFnd6g1eJ+L8BnShXDzbCNI2nknWpt5MKg
vFOg8ujvaUC9mpkGKE2vkAHLA/EgDJXgt5XMmbiQy+p0WmD2WyKWSzrkEwwWW0mtZXsuwYoSoXBE
nPzZP2HYdIE6/n/lLWQnVb9wLEbFcW9CSA6uaJKx0detigMk+XZeNcucMmCoCRr2v7/Fce4GmjEe
dVupASKin6QQ6BXw4OxyI+2giicXcHrKLSF/vI22AQIj2B3xl5bs8rhqSbt2TQ1ATcFiiT5emsrq
eou1vSQcROocV3G32O2VTZLOtwTz4NU8uyn48P4eVcElA3c0fQ7X4tggm7c4MmZ6VFPBJsATAM3x
izN3wrwUw7s5SeUe4ZC+9dDMeR5E8uUfFtqrKiMSnWI0Hgt01acTJa2NynQl9FLOWP1T8by0VUZ3
1hcE+kDdBvVGiM1yKRYHu3oPbv/jKZPPpeWk+dOGyrJ8ChbQOqNNhk+kczcArd26bn+p7J+dg/Ro
hOVhYCRmxT2G5sYtDffzXZPS2vJvaH55CDn0ZXqEo5TY6rkiBEjMtYJCgX1MDTEuOYr3A03Ij5Gy
N7KexddnMhGrrubE/C1Y+dZ9iwqvEIE8DYkulTofsEySV8X3U359Jgd5WSkWOwZtsMs+IZX9GJpZ
IX4vFpfX9Kxb6eAizCScM7TWj6O+dxUemiWE4fnBTbZ295zSB4qYIg8MLVmZC0IUbgoyV2yfmOmf
J28CUcl3pm0SdbY1Ken5wV3ZQfEDVbkwn3fbvDrQbVFX/Hq5Ozmakr7Yv4GJ7qm1DaBDNWX4nASH
qV2Fv3aIIQKS3dvZbMZvmCTAzBxjgMyjsho8Rrt5QECKl3eo97lKAhIATBUQMMr52Pw9PTUne+ip
jsnkq/EyjoDSzgIUH61eRv/ndaY7iMEtKOxJXmXNEA6yUmlPwDkUeLNAZcUzgsnRIRFVWeFBwbCA
L/os21BcA7Eiw+DWShOgqjNzUHoAtdPeI0W4m1L081F2EMNpmLbWaAHyj8Sa1gzAARMLjXbI1pS4
aq1KbAKUSa3O7KkaxXODDgDraOzmM3OsAlWYid2eyvsX8WG2BtcpUANBGYBbEBVacfZ7iyZRnQGT
AEenYJVQ3fhhacXd1wsbJVw5284ikAneSyvVllEMrq4SH/ot9fdb83AKZf2C3+IZs4RotsBE4w3E
4/n8k87bqi3FT4F255ZLbcHMdcnVQHxlJaizNLUb/ZKxXJL2op6PeI0+eYtfjHtUEzprvDoR0D1Z
sC8TRnhq9787oWnY2xMYGDZ0G8QUNdEYqpWD9aOVIlydYyvxxy0slxfCMlfxOu27dRGf22HXf5uy
28f+ilPG5gbEme3ImULan5AKy/is4nnsHWDOFBCCOztmjzkYeeXwhqtn5rg7BkHFHulu5ZI6QuZo
DV4O8pswVll2ERsoFHVi3UqO1P6UQUYlV2ullLBTRdmhZdNIBsISTn6+qwW2vQxgrfHhj8IDJYtb
lZKO+MODmIln9WU+IocFWugesWtz2fdKEoEIn1zYO4S9hI8LSeUCA0G9piREErbsJ8lbn1dFsNrA
j58GoE1yAPyBimwscfRZh5DVo91Sxkau5IjBT1n+kepe8hpkFTymiIqjlvX1tZan9H65ZXwHmY+y
TGgJOO6d477rfwTeh+h2Blj7sTp3Ol6J9PrOaG49mi3qTsEdmcA5hiBbN6pFERloa8JOm36HMOhz
ISvdheHThYTklTfCQbyt9eO9ipskeJkH0J+Y0fwMVgGiKnmINIxrosBrXGDlAlHoRbNTxPlriiAZ
kiJqxc6Ya82GvS0yIPARWqfgbufQ75l9rKNyBnIs3XriEUVy1WO6I2oYzDt5b32cRyfhOwkxo6hd
jHVBr2miu55fTYmx3OAoW6up0d8UsFuuemmgpckBE4yqlr1sS669ixhLfgI+gOGUI3B5/yB/8jOp
NKJPtPChiw5HGI0Avbg2F4d90O+3/Bk0DP8+EfJtlxXGes+RBVLFUbg+1m6EHjxh+lYJ46PWScQD
UTP5sWYQnDFkTOo1qpP8Ta/dHegGRV9PXMR5EAb/WuTjtfUiZRRg7gch2XB03P/AFHr1hcdXNko5
fNy6h2exexepo83LAXkrHboL2Q0Ej0lYvr3tPSp5fR/srIIidFtebL5fqSR0oi1We0OmhJoCHHlM
qA7zBA8V/0T1bv+WQl5CpiY5aQ9I4ci1gnd5Uh5LMrj/vla3im9pfYSzaXpt+FM4u+FZgDTLJgMi
2pd8gM/1jxJUtSBmxQgkJXjO6FRB0zBg9iAFJ5jl5c6JW6LQ+uwZ9ZShilsvVukFVgx6ds6Sl5yW
2BOsIqAVFEuXJGXzYktJEB1mlM6yd0XQTfAX4PHEhmf8vRRvJlbUmfEb+sT/Uf32xrolOTTJzTKY
kSUgPeoSI9AEzKzJW4s9dzDFNGo3kd3sfxTVFmE+irAZGkRhwrJEhUIFRN1uRKe+jXgpaNSgmz3x
yxhBPvzm9Zy7bIV+emFJ/SlmJruNzX3jl0Oi0uSqJGtFon2z+RRwESzaW2mbe/WdpXEM05ndIVcD
RZljETsq+inRPYLn1yS/3PIg+wSo1VY7muInC3D4PO4iOq0accQiqIobqMlLwGNL6qTXcpomIo4p
cHCc5iGvkiisJyvgLVVKWKWdRMKm7WgrwQL02MuZYOv+cucnN2G01AkYMfQVSVhCUDyHrCTSR6YP
WgYFKuq+gDU7cPyTYYC99VRDWhvQXDwtYhedlvyOxOsNz9Th7BUPVgmhVroGxAJM7vN6BncHZIKH
gRcHSMBJ4d71S2HA1bXkJ5xvw6wtEaVpDoKeG7QwS9+Bgx1coNIN6+ZpbMrbDhx4ntRaNJLXNWxB
YxQjSBi8OD9Lvxspv/eDmfeGAjN2ED3PaLZfqXUG9WEU8nW6rcL+cbVQcD1Uf8FnInuOoTVC41Mz
zZd+Eb4nTtgXJYSE4VYpeCdAUjEvukZN1P+OED1QqBrRuSy61mc8U4vH4/VarCx2ns2WtFWXrvc7
iJjgxmo3n9o99b9U0MU7CT4d4TY1gnx33L+GTmQ+QvdYiyxv6a576V0WD6VZGfagRpehik81B38Q
asidGipBQgvo+t720rKfay/cpgVWteJFdTuupkKTpYT8a422gMz3+b0vkKQwVk2PHvRhQbYBkhz2
tThV41hlsOli382w8abKR1avT5LUKszvA6ETGS0cgm+J5nrUfy/SaM2hV0aKKddcEpo9RE3mmTUG
m8v8lcERvXcX0aF+v/HvPQZAhBLue+CSUqBh+aAdtxNYSYeDw3slEnrZuvl5QDZyDVmj5Vb2jmGV
x497w9T/Snj6eRCOg+cchzPILJDMGuXujOp/b6xL0lDAgUZt5bptGdSl8BXR3rTdEotpNn+Lz6X+
oQIe2VWabTGDwl8z6t7l48SgDlofvFRXQraaR488RjVY288y9zNZJlzWO5opWIp2UqUL1H8ZoScd
HGvLJU7FnRZcOrCG7rns+1Fr35W4meE2x5gv720WClN6xSki0u0Up6kVnO14PFKvhSPDUlgBTgWy
ZQVpUJJUijWc5KCoN6KIbH0lngaHgGN4kj3+e+dhkZvr0ZLoInT+e7M4izhzpjAdq26Kk+yBpxgE
K2iGPqfjgygAh93CQYHWqO8caquged3G2J5mZqyGGDcaNwjEOofj+bBVTLlEMisM3zJNcemnx3jQ
jMbbDfeMqndTOcL+/B4+itsJz1a50mTyFiuBYLAk8aUaYrZWGsIhMS1L+VaCWQ11E/KmT7GagGY+
Y3NEXPT80X5cb5KiElmaXsUIXqn4O7ny3oAovC43Lab3KB/XWrJOu71kTiPhR/nyKCoElcsKfS5P
1GmDPaWCZIzsO+EWSFFAhGY/gxyxd0qCmoHJC/1nhond+L2puAOppnixrgkW9kHb50EvbVc7TzwC
Gq6ZKdxpb/JXYyO2hpTzMwHVu9KjeRPfopTpDRWh7rL/coRMQhxX8G1tVMwwU+9h4voBPmfEs556
zmEPd/ZdYMsW5JP7cMAdmj2Wt2GSeHc99JEcUfeX8C8f/+luhsHK263o0sEOsVdD2/dVfAGsARJH
fPuH4KgzkJVg6tQChCS4fd1dPGS2htPp8dTIaYJu12UyAeuGXQ+ZQIGPb5SXr+ncmkJs9gBB9PMm
/654f9EGdnRW6bQ7jM7/UfGCgIeRgHYwwT6N7ddcr3U6es18YdLR7z2d62YyvdCsBcLQ479MwCP7
hnWeZjiWBqog866VgJfMfYNE6Sf3Z2yR5dTb3G131QZ3ytFQ3mlttmOsO1xZumqo2vAbFe+XwEGF
QOjDv9BicVXkd+qL7eqmopU+i/HbZAkk+lATS66EGEWZKDSDL0zJvsILyiwVuKaLa0YOgh5HCaIO
0wmDIoq+nwC1ymYT2WZ/sQEOwblWkCuJGuccKFEMK6IKiABNWlHCW0TzL6dFXhQ/aFVryahKtAiR
n2rMFiImyliaeXpOmBnkRWbKvMG8zOuZsFmIfyrdbTg0MqyKwCH09TLABao0rxt0VJmAcJYiUxLw
xWLMawzMetZ4aG9EdiwFyOZ+VbeeOeMWMmOHNjsKh04rAwLLof12EdUJreQ+T6km4NAdCN+U5LKj
3J09/FO4cs16u2XMKx73fEj/FDIDcLPdWKfZV72eKO5hr6SGQL99MeDN+rnKbdcTv0+G4h1baKy7
WJgB78UtjBEWupM87tD96JFM7iU5FSfGl70yceBkb3qvk2i9S0GySUFN56VUnfFUMcd31JI9jCAf
ee8AUcQ0W+y1VQ+mlsJFjPa3AxJzGbjpG22WyMri+7s65OQLlD0alBKenm/NwHW4rxCguJ/5CtJ5
dEe/pshE5TAqMPskVoC5X8tUUTZwipXB4xEAkp2a/lMfltKTSyh5AXafGJzNZlbchvXynAQnccrV
IkKJHG8bGfJeBUY8vOFJtDjF8mwgf4JF6n781imRtwkXcVQrAbOkRTc7GcfggSZOGDXJ3v+UAKY7
ASF/15V/TrR8iaIDTgL/f7WOqA26EItCcIX/U79XtUK+JoqNmCWfJgRkaN8CXRVfcSrsJYpxOBcL
02629AgaNFOVHvwQ4tRDv5mMXg2geH7DS8WeCql7v6j+T27O1g8W8AvRdBaydVCIjIuKTuyJ6LF5
L6SizkX+ZRDsqIRBPREmimWdIHjZwot0Bjng/rhQaYOQ5clNn4SJdjZ+D2YKcfoVO/mLm9dXqqPU
VOda8MLtfGSqSMZyKco62XYEGVq7d6vvjl0I5rYNwfyCt3Aro7fFEIibUME6BzFx6f8fgNMzNtG/
CyoRVJiuvSlF0rj5RCTJwruyNyCeDVK3BQDxQhe2/PpyRhQGGqBn2L+ZIvYsSxfTrMCD32FU6QC9
GwfJVu+pvtlLsooPXQja38ajbKgwVUyPJ59A3LMNSLEYvruZbLpT6N8mMNBj8MIXHsj5aTwdcJhN
ey8tUd69OV0g4vBZP8RojddUOVGMM6CgQyVMkVYylBAdpje8ZKsSWMLkiIytru2lRmJBEzfTbK9b
mEQyxic0DEVTYIwdh4xSH0ocZ3XJcrYCUCIm/CLmR0Rs9eKPw1BTeu48UAFwe0oDd6obYX4NQgjC
gntIdPg2DgFR+i7gYGubNBJDxu1/JLIzjTBeZA4I4uWH7170zGOAb/lcmQ+PVnVaZTDhCzUl/myW
LyNcX7AL8lmlP1XUom5etuxF9EBv475eX9LF4VQufFboz3Sq0usg5iSs/jiJXsxAHuDIb6zM7mo7
UKGKkg6p85M7g4j5LKh8MKUdX6tORy5SDK0SKqTFW6zNbI2ytZ4LF1fTeGiuUXZq7y1Au2bcI83z
KrFVDIVgqmMxuKFCbbd3IWQerrRHoIh8hnUzPwPKRN0eE+ADjdAmSTAZicsxhvtrgnznaO/QBzbv
ZAWyShuLl6haUrITqXmFO+5cx0P387zJXg4X+lRcw3aNimu/jGq2vfcMxVISYc79WIiGPu4PRnRv
NyQaLb+FyQ6d5ODpu2gFgDTr1UQBCLIlijzbx4qZAEgupzjFisxP+iT6skpzwFotnBM/0Yn9qF3J
4UGfUEYqEgj57NhrvfEdsrrM8Kk+JSvyALYSkDuzN3OnqbnugX4gbBPUNO4SY1TBNdiez9LEumJo
HIq1+jekrXYfrdAzTFEnj74lsK5L1vrEi61NrF5I8v5ZsjEFeQYzpaXwT1CTD/yzdQsBETj1vlnG
j0Ox6sPcBnqquUzMhW+lnTcP2btCB354Utf5qy0cKtxnO5ixcwqnertDq30VL2LwAfZyN6Yczyx5
3CFqH9u9PvBXzn1vyNcmZ9/h3dFPde4hTFEmdpKNE32IFVIfRRvats9P7R4b8g51uTknBFrkn3H3
zV0BnfcmZrFDX833pHeIGMV3r3oD0hORFRg5QyPyy0ROILFDDmfFnPMqx0KuZd1gMTvmAlxOir74
GQM9GpknuHTc5IhVDgq1wXqb7PdCW+FzZ9fWCkUN/Ofgvf5pH2aObOZ+hQL+06+ndlcYSVVz/eBc
/ZB+sQPcVCxPASJLHMTPPziSWUhS38+iZkxWs3aCb/p525xkzKPBotia+V28Zx5jMNyw9OFzeD38
J+ChmE9Zi+VSYYEcLU5vrh0NqkqucnwIAZAwFWBJeZ6kYK84UgEC96AK7QCPBZ7lCdah5skedgFw
EkXPy6+225oA6tCZehSOYkXNKX3LVO1CNcOWUG570+p+FA8Sg0rHvsD9gOT0+8MKWytUPHB1wxM+
bZ2Rgv27Rr78p5p5KpencKAwFbtjV32Bbq7AlHWiY7mdDjyxBYH47QWbx2N0NXu3v7iq3azL8Psf
7INmm5Iw80HqVCLHNUYE3XUMVnFFL1Xdv7DczCCABhUMrd5kDIsc+CxCPfnKXZdqS2gOz+HDUd9q
5N0dczadSO2pvgGib1ZjWh0GIbzeBxIvtYZIIBtxb7V6BluxfRfOXJJ+V5GMCErOoECXMZgp807J
eVWfoH25YwqHKpjbjc8AxriCs1RKC5rUo9MoN5np7QhlY9pLWxiLAYNVuYFyAICR+LfzmfZp+Wtc
1FHXmXI1qd15jmCrRDQONE4CVr1znd9BKQu2tK4JKP16f+ZWN13H3rcaKKtHAxuPDWmZ68mNC1hy
5mUdJ4XXC/+OvFtWP0CMKfzx5WHE+i49qM5Nxe+TNoifgvMRcLBx2jSgQfulj+W4BE1QWLTu4Ju5
BK65RKb+gmbTk9wfSYIGRLc9byeAlVsQ+oLNl+pLwjkxDWYi4eYHwlgs5HozX1LLTDWMP99R393y
1tkINAgFo9l+jOIdx0DBNH6YHgkiss//1lZxLGNSsHAjpVzlPcUzSO2dHJ78ZxvT+B43nhe7aOpo
saUNkr3Z3xIPHtfwjPoaB1o8oiQESO/CZwJJlKcwY1zIbhe+ix5DFOumJFVnIG8EepyfhBlvmx1Z
U/Uz8/+vk22bxT3ObMqpB2A3QHu73Kdbzpyhk9d7TXU9qo5CvjoDSJR6S43qk2tWX8AaJ7GmHCec
wQOu5yM4bMeF+5EPVzpEVuVzTrJ9ntGHCo3tAtKBrlB2xW/ojHfZer03lD0pn8Yi7dSWXwqvA/me
Ikn1afszcZcU7N2R+DNwVt/NGSSljRBl0cTQVfO9leq1H13rAAmu4goSkvl2d+6LaR3jb6oukD7O
UlD189Y6sSUKh86qDooe3Fc5lCfY0g/RDb4aOtMtB/xfSLpuYlful5HOSjF0MDgDsB2mMud167br
6ekLFKM3lK+VUUZN6S3iRJLgkTrvVPw/IlI0jzF0r8zcOykZtpypawF0sOrZMLtoYr4uh21aGc1F
aJtMJ3iC68V05C9K87H+qalwlVGZkk2guGZhdLLMw7jmu9bMZHOXOMhuDICLA5ZP9fPmheMaeVif
9IWtt7EyNDmnTFEfqlBZbbeBcRoqk6WZXSVOWFL8VW3+iCuXTl4vs9wxUaNTzpFMxPtDGMRnha10
FKG5YQH+NosonuWkbApvXeA9tcFJOuuG8lU+yBsgJ5T+cwzGypwTjJXTsoj+L5v8O1ubjsnpHgJ9
0kMl7foBhOiuQSmy66vepsKsfZ+c5phSYiLCsnDfS88U7N+LeaIcPM+8sClOOYYrZ/1W7C8UOlg3
CzFEVLJB1qwiR1MfbmW+zaV5xdHNgE7moW7Pmye5zPyat1Gk604ZKamaKplX5ucS35JVqzbP00eT
H0wO0BdZOcUsB5XC5qadnbvp3kmZ4XPQw4+vSsIcWqwID5ea5+WhR0+P2+IiHXVWG6ZUMnGJlgEB
Or3Im3GNGOa4XU1je01+uB7WIKLiBdvds2783/z1pyTp740rUNKmLUBAcFc9UwV4qwg5WSpuEef5
jvmKAmOn2Y+6/TOl0QmlSQbi4QI418uWnXzKSTA6hqeA/kXiM6CTemJGemOyGfyUL5ESqQ8XC93n
xehs4xbZXCv8yZRa7RAbWhbBw7qeMS8+OLbueQyKWVmPCQuMC9+4F4fADQq1jRVz6JRq+qrXKLYC
rtfYqynguUuV3MhAfr007px7E0C0clitHBnA7mM5n+6awVXWbgCjB7KPfAZ33+hetObDxinb5gO3
WMS8Iqxs1ON5ZLWjhyQA/MmYUsjjdF0yhXSs28cmrrQwnfwM79O6UfV0V5YeEPBW+PIZW0oDhAMV
Kepey0q3QPi3saFjPnFFuHuUrvAPXUMyT+i7Hu7oHS5u9hnHrDxEFzfC6sw1n9fQpX2OWaGonB3e
yjt381cN56pifApL1PLR2lfkvd25HSIi2241IzUYuBsYPKm/yUuIxwRIetqGCqCyaWnYXZlvMWyL
xRZKfrFVz3N/GIvOjJYodVw8ADEZe7Q9MMuIxkrNHM7X5gpib8EY22+M3ZCMq7sxR85FE+S4ruuY
1T+Yc1xdssYTZXrrvSPvK1jH28sSAyaXSsF4O0PUDb0GKziooR2212qhdZAbfO3PHR7KPfo9I8nE
wPdjwRkyK4bomy6YOXFagrCJcy7AL419pPIs6V1Gp6p5xaoQzFBx049kyDU//XPhi+BlS9scpqqH
Wn3XcYGhb/wpElkqW1p1Zr7ecxJhlpBFmXBoQbuCeV9HtZILwhQMoJwdt2szwbR1An8iJ34ILf8Z
GmWOj7v+HR/srdp5752CfvqS84y0hJNumJBDQX59d47XNt/eNEYXptoAh73N3sA52R/HoH4E6pbO
KhGkyM9edLCJByx1dszaKjpe23PtS8+qxULCVENzgdld6Fd1jAlnoJ5wnVfJi8YmRs6lfpOi2mn4
JTxntCMo6vTeAQmsTij+MhbscRMXg0/OQKbgk75v61PHVrIwl3Kn0XLz8J1ksLhJitOoynb7b5KD
K3zQAk7kczZGGpwxehPonPmByDBwBnMLp+LdMuIZ1fMlwAnWy09ZYUaf/NGce0hWD/4fCW5eeGbI
aMlbXwS7qD/IXc0hY7hZ3VHVy3OllXxsUK+sRglwuc1r9eunI+MdaZbuP8SriZDcU3y5IAAVrDlT
JaybE0C7eoFz+nYBA9c1O7HcfHLfmUujBNLtOrmp6ThBdEiaqq2HuK8l2GM8UqmyCzjjXia2aqJi
UmvQalNddHG8S11HwO/9qI2VMr2+RgSW5D2IbJB5S6//o+R1BGZyjL1DKMtPp1BJRhKSxTBzsNvM
EZhSWiNJtFer969B+dpP92J1gy/EqGmg8bDjcI9q1+E67susvSX1Hth4GfOrhAwrAdejNyiUCOx7
TkL6BwMffUbssJSOILM5sF0cgdEB0f2xua52O8Lj7zfTCH1HUdhKarDf0hein5wyHcXs7y+3ULUz
QAowpZAO3PH//JD4/oFAA8SV2qaHRj7SpAsZ7bT0F0a0uhX4zL5tH587BRfR+nejrFlqvMpvZaI0
RgcKZesBR6Jneu37JHZqzWVyJcmdweZifIxYh8U43SiAOreAGJygwGF3LIdwaYd2PYaAryYDxiKn
Fshrepwi/KWCCznxmCFS52A0f63rFUkDnO1mA42W/3OkNVReT9j9Jb1bKwF4i2w8kX/FHUUCg5h+
4E2r/w2ncyvGFqwiQA7wgmXhWb1wtH0x7vMh2hwAc3r1nOgQem9diRCKoje+XBTta6Ru+cQYNi1b
65hdSI99Z/cPZ7A17HaBbOs0lGj3EJtzm4TVmGpFJ+QBsr6+K77J2jp3V0Iid2mHq5vgM1eGWY0i
fzEgW853qwZQeMarQpBNpAB7xJmjVR+Dt4sZr22bEqAXgm2jVQNpK2ppp7/SG2CJIz41hqs87Ox4
nhlHuDACliaTY5kQ3ArO7MbdDLj4jB6YvhL3gCJi3WoFEpC409ScMmiagEbvtll7hJTX4mwi735A
xhnYb4p2wpcLntG0P7MkizoZ2hbnceCKhkgsIpZzl8OXrDrAZx/C8BqzJ7qcvxYUidqKldx7+GOL
Frz/BsQ2ZW5qjIB2p85J3fJEFLeJKU5KIjs4G74T3q8N0n6rLTmcYETc4XesQiLhMyRpPE8aayDo
CoHfCth+XGhxkSa5RguZIoRkMVYwwjqwEzYRcfXJlo+wkT7wo4wUUU0pdyw7haRbNlIpisG/ncGu
yyC9P5eoqLjBbF9a0fiZnC3jsFRNvk3ElqP+GMsByjgYWa2nAT9NHn3u3/fZBcJIG/EMTF+BaXZU
5IFuu1K2xDwv5aK955izafk+uDDVmfSm9DRAry3PrrUwDh8FM9O1AZwIYm8lvjc1XbJinU3TeAUL
eEAAhMyNJoMv+bIPK2sTTu8bL3hqUc+DIs9uRS4LypcwP1bOIgHyGfqEBTVWVsZxaT5MoJnYwNxb
w4YQTP9TBcj2kUBt4TpU+8Lv3zuVKoZd2VYINhH0+oRjSbkecbL0BWq/aqGopaFnLQWjdhJhMK9B
qY4uK8fZTiD8BxKJjp5CJGTcd2hn82VuRPXfGdsdmr3eKNnjOA+QR76/ABxtIQpxd0ss1jY7Akfs
HPQkNfeBct+MwpcyYZ67UO8x1SQZ4i/t8fFZkxTKUY9kpqN9UunICnqzgbFkPWel01rI0v7/yvJK
ZqhfFGhbdpHIvGIKqDyOoFXJKm4HgTK71gyM1PwmDrhLeTXyNVxRyTp0kGhjD9jVyqeJ8z+dx4Lq
JF9Zraj5VJKp40/WqBJykJSZXAv2b6ZZdyqmyrFF0FGIPzP30ciV+ttyuVuXAr1djLrqs54dqfI8
l8wQ6gxCNaNSic0iq3ErpuMG/uIxzsQ8Li/98xQSN3Xa8TwjUkSP5h2B40LLZb1vAj1LQ/+pA2hj
T1U46HADnsnQp1pNORySIsukzdB2EdygaAbn8TcWfeyvElcLHdzdA5HSx4Wv+Wj1tLwzmZNyJ8Qm
cwTeSnv8y2551gG2Lkex+ClWJfd5MGwxGyGOguAHesn45at33iycpGC5B5mXDLnybkp9pDmxGUGY
MPm+NpZTH1CPLfd0g9XqSFSf1aPi/0STPMwC7xisjtulHaS3xHAC1modMM6T1ZRsEHeQhbUBYeFK
rEqUfa3qVPCBcY15XbgsQjD+61wiC0PkOMzhplYgd1kUvoinB5yNZf5lpdKzYxXmMN6wekILUAEH
mUoY5BxBxwyloK0E0h1/GzKUyb/Jm/z/vP88mNqLYvFChew6PbJoFG+Vx5WwiG4q/BG2ZkAw8Hkp
CQh+Cc5BWS+sa9Ivji6noIcX2GKwwrOd1NlIqx6GYcEgCGjjndEcvEobOflgBnMD3pukktn6cSKa
cBwj04ll09VbHx+XyAZfLwfC0rLcDZlgdqLn/SO/paw65y26Qe9od6VefMIxdsANK69ZJi9wIw3S
JYxYv0shpvkhhplibydIlcWEyiGcC3v1Dv0q8/ZsApi0Sb6iTLcPLplkNbFa5PDzNcdexXxahfz7
C4DpR/1KV3gWfLXJlxOtqJwjceXFPRVL4PUxqe8Q26mMZr4ObFrKiMnXmOr2NkGrrd88EBBXLBUf
cOv/2crWLDjnV2MIASKil3aFZ4F3tadqQh6tjisoyBGhDfVsiGWSXBsy/dvzx+wPRaI5Zpc5i6o7
i4jy91rpUguyzds/8faWhblODAUWvVY2P6iLxMTVBloIMLGNZwytIWwpz7IxjiTSxzaaI9k8eZAU
cve9NUK+z5JU9g4sUUBKtvAM3Z5NE9V62Zg+QtPtk1GYArnO5swnhLTBXRh+SQ2zlRNg3NcuG+5R
qD1e/mCew8A/16gSB3JlOsMIqFLqotSsm7pOTxDnwqZdtYuAmTHkSh7EUWYn/AZz+9XbRWy1mODi
0lFmH6ktG+8gR+mj1HnuL/6burInniP6AL5XEYTcVFxpEeGHnRorRQv2CmFyDA0p9WumfzzaLtOe
1rLO1qnC07De5chNO1YMV4+KXOJtEZB48CqpNEIZdnDQ5taFtDzluX3+AmM3Q874SAhq6kSUK+fX
TBp+yaap8Srndk1Opc5vXvezSPYwAt2qsASMHSmDfBgxj/PuRaYFJUpbTYTcgSdKvbSSwndei3NB
Z2EXXsGzF7tchNLrP5Dt61mSs+gNbqxPGuo7EuE3Krd3SKw1JjapPjJQ7dv6rT2Enssi/doxqF/J
hgd4inkq4A8xJTDWoo/rrlDojdM1g7Mg0FKEAO2Kg26uWx7UBZCggzh5vyk5wwphfg+RqyLveNts
gAXb7ZpBa+DXn/GRwehLAUgZs6kO5kkcudV7EXZJvErq3vTRaX+EYoDFulIB4RlvwyTwL8HTed1e
iuWeoDFYbSJoD8k1KTsMaIyvFD5ZjWUQTZmAaTCkOtttVJYQ936msjIIRNJnlh4Nnb2hV2647b3Q
muKpie3jwhf4EqEGlyovI4iNOCDrodHo2s53ByhfPiVhRn00Beja+NB1mrcGLdzIUBKoy3wyuO1Y
nMBtJBsXQXu87HUm89ISJdb3PcF0pPM4No7E4iHqo19M6whtP2v2Cy6co/2xPq1LkPB1ju60LPCa
S4klXEApl8pfVirOAGMiu38RAXRMFjp80YU/p4jJunk6AAWwHiQ8IROFMq+5bOr2IftH5PDIZmFU
J3cchxLZlKWak/ZHt29Pmt3DuWGXTXPyBaSaJjwrdyPHI/ZZPcfk1AOXRTtD68YS2oHTcoVKclM9
px5UOlcKEJo39Di+3glbMVGa1X81tbRinfk0oB/IFRqgzgHm0I09hmpjqFGZq6xtX8U9jxWiVgNE
ZMqmK+tJnYeZ0wiKOVtfMOJ6qajBLDzvOhYAZVuir38b4fWhyy/Zo/rZDKxAyInl24aOplRSXNdP
PpYd3LlGG9Ded2bLszQQGDqnZceW8Lip15xb02lIKBcEi5Ypfe5LeHhmF2A+uf7haEhmYe2yxAI9
cpen3kW5QqhwImDXyf8sl98gvf/A0we7YlV00iy0gNCW6HPJi+duMbb1RPA3CDAjEgeK6p+vbu9D
anGBxvaamxIM9Z7hM5+UbRPAkQHhUeFIyORS8NlvsOoQR1q+TtpF94ctwMnJA5G6skpi3lGPA+4u
PFM6X33E+PIN+77X08Kz4mSmqQS0bNPZIoJuAXeSLA2kpSWyus/hAL2zddsD0tAVNdaO992Z1ZPM
gAouEzIwiq7SXv6slipx0DSZcivJmQFuvTBZ89YqcuWY0n9PVtlSEp3dq0ppdgLNeHhh/TijmS42
vUUozJWE6heEJZbTaAb7VYfpzsN4aeGsHOJh5dKEzqww4HEBvNcW61vqzfgab9QsumArBI3o5S0R
tqkP7hXV5hz/u004QrwiM8fLOmL5rwpf2tSyI5nrOVcCnhciIABRx9jsuzBTXYTd7VlZoWTitksm
jJNg+o0rFVWJN4E8s/cb1E7sWJbesEKPEQkZIXxrxryHpRfmJT7A72WSJvcmxKA7aCJFl1+mVGHo
KYCxhxoz4lR5ed5YilHmheiBDgqw5Jgx8kkClR6twC/tqlDAJ6Un8ZnPs/zr5oCDnKN9bWpB2UhS
qtm3dL1uZBOMfj+ZuxA2/nE2wK+X98blALLpf1m3bmKYkX1VZPOL/LTAX4YPujn+lqdmhLVoyK8L
zx5CnDF9wtT+h1r/HnVdX3IXSgn40KEy7cl8glAijw780DHm2grS+IwreVzUvwbc4X9E1IFYIqjc
tdRnSnYPC5PLViVkzTTictSzT7EZegj67wOsvFWWRjcAP2TaXrIHjq9lApvnttY/Vp5/wGbchpUy
LbLaLqnGnj4qn7ocXoTe2+EyU9cZTfkv+/PrhZxVKblZIs22V9lCUn7fKVsRDCE8q4qGSe04iNnA
Rxiprmn2sOh+pTN7wGMtiCGa5gpDTCClpuYZTJNSoBdxFL+iHUUYo4ICeIty4uMGksRHWbHr1zUA
TbsBhGK4jZSstmOWoN+JSTPI3DNzZiHfnxaccUGxK8TNI+nCZZA/fkwjRuu1RigSStl6qc+91BZh
+PYPlvIVerOwmMgMK1tZGEXIJK6Id492/16RI6G2Il03NiWGRsJvTFYIWe1kptwj9DOjCbwBPqbo
2axpQ23z+qF7CsXL82kiHg2dT1dU/p6050wH9SxO/VU2Zfs8tx/bXw1ymQC4k2S+BcWCH9Sdzttd
tBXMgJzuhrctAcZJHn6/nckLEuWoryehIZh8vxcVO3rFnqBIcIV+Nlos93DUghxAl4alR6r5MLSt
Il0HHBrqhauV++TGltAh6wdn3MK+PxXeEnMuSyQE87BqgQsb1HhqmgVWmJSkJiQ5QIdAyLqiUzS+
epAhU6cJ4mOVp45akDx5nZxa+1qoXi/Jvhq2l3SFaMirWAjo77h7HCp/D1tH4e+J6z10mcyOzlmE
oQrb008BED2WZd2QiTJ1N9VvHHHwKb25ru9dsCfnyJXkmIWz13Hvy2hQgTWrkzrlF4klwRKEWGCa
BffL3+1aEVc87gHlkY2edqflDNXwRysYHFWr08fNTr7C9i5DGlx1jzNlSJVOQPQJ3L84V1v3Tf5w
46pCdAUf2sTDrDRWMRhmxi6De+KgLd2ix4eWabnru0W38i9gmEKffc8vuG5yIO3UTeB7bTnv84b4
KptjafJyWQBoOHTVHXNnJfA2ZUinLGIuw3JAOE1XCh2wyw+mVsHjjm3hetai97vxdzyG3Mn4iVf0
SDfdCDCajO5E+mqGvy55wXbMdDY0JXYd7Eh0TLsaFfAFIFt8WbwY5xkmU3111jSrKug9/T4v01ga
5uq7QqA9v4ZpdPZH4DBragDV53VkQMoLKXcGrgxmQSUPFTUPWmZLr4rV1dOXIJAWqIFtARCsPQ+s
/JuxfG7RG0xyBOheVztw64YlOCkYMbRqohyc5EH6eLCp4V9EA1TgFXwKQ4fIzl4/O6xRIGf8YcKn
Sc9mrVFRDm1ycRBdEUngex/MuGQzUuOO4fMMgI4Jkagln1f7C15crwrN6zV6SDMOL77F7dpxDMRg
vCs8ITQe6bB+bkdhUOYdpKwHHEzGHXDDDBZU0+qHLAgEOpsH4R1q2rJCL3bvbjjV52Ne3jz636bq
nzI4Ilu6IZGb/MF11O9MqDKZJzulPodVeX1pCtlnKgdj8q04/UaBPqn+o/rPU+4bOs7Mwf20Xtkh
9Y7E9R00ktv7/f3uwVZ9TWFLI4wZWSieGPq5TKUI2oEF/4n5vmU31DOQeCipN0xV5TPuHsc9ToNQ
pBojg1D/WmsiAAsdVmh3ehxNxMJJOBpEr0UOOr8dMB94BN5ZYOO5IMYdD7FtXb/C/nYMiDkB9ekz
Qu8fWYGC5RjSmnbs5Ut1I5iHzgljc9SRknmxoncdxVBe6bQJwfsRDlhHwz0W6QTYcP3IdBx8z6qY
6iLw2NdII8UX21UvJa7AovOQh9lNJb1D1ug65XjjYRHZXZQhnpTd/uzrPYl0TRw6u//XWLPavmq9
RnnY4T3r4a9QxPaT+nk4HdMHeN3+HAFovoDfdnlMGxub36FtIqdujFy/uMFzSa5UKhq7bu/s5wG1
P8V0cA9d4dYCy0mxDCxdimeng0e61NdH3qDojQOR+7soDH5MNeG/pZk4ZV/d0McBN+CMnkAEB1UL
rOR7jUN9jp/syHljj0JUGfvWegsOlxDJc6S6HnqFEsO3qDMNGRqcKXGaYxTFs7Wu5ILXgBc2kJ8d
sFiESIKkJpkmN4NZp+bM9LsAFeZKR7K5GWrKfQSFLDBEhIeOvMCJIJWn0KScqSKRbLTgSWOPrQkH
NgMTLuNfggN5clSbf1l5fl16w4f/2k1nNnHV6sXFeJAQ69+jQwAU3JAXfzPoY5gPShr9o5WL3V7k
iq3B5wPFCLOfGRIPHxAiTlde5tolG2egJymyVMz6LWCH7RQ9Mo8ZwDobTKIDMFyZ9ammeM8SgCMe
yxiAqRN2lNRGfyUOszx0B4R/LxngxapZdVDXeR8v9+c8V+SKXdVV3re9XBmN6jZ4bZwzxQaV2Ow+
7WIoCbkl0N0niW75oayj8oEvmGvlZJqlKl+GMgK2zezdEli1XCDNQk5ACCWSyWl1wJiimfuLrRju
LIgKXln4aNqGYZ1WE3yDy2TMIp5hRLEaMqhByiO3tLhQHN+bfWXkXq5dZ8epSI3ER3JGOQRJO5n0
kgwxUKbpG1F5iz5ysraHYXV2SVgS5M0oAOCDAIL+zhnjTX5QgKg7L0H7NWoToipSb/TLRVh+Om6T
VP5IBqEJWLdrwk4dEJ70c2GFZUwYbRl3+rnhTMBBWyWLoHyiSqHUN8HCenHxiVO03XIiBpbTN4eS
0iCFl9lq03jDXklxXcArRTHzXYG6jpvbUls+qLwxX8DQk1IVG4aM0jJd2zIMYn7oLhjqZUNOw2YF
LM9wxupOTDx6EoVpjknMAz7y8Z3mPrYxMvjZAb0HQEYfC4q2uiS4kH8UYXAyb3qp70Zfdb2LFSbp
gcZ9f/I8DSW7sd3ourBV8vpSNhRKTno+XFpDXF8miGMurDE9NL6fj+/6ee2BUKxXqBIsk6apiCnc
jXs4suotera/wbF09TX3JaqfrSH2oxGXXY7FubtzX2eUvUadmEWPdz8B/RSmXFSoIw+nEw1ZKpmx
TeyaT5wlbxom8oU/qFtmbOJ/hPduGHvWfiyRRLKU7Zd0KK9Y4bq50T9zFg33jFJdAofm90AjNOpb
zIjBCK+SnwtLg9UBOosIgGDAICBtYOs4AtHOp8Gw6x+y2ODJuJcfC2qP6RB6kvINNEhidPU66FEz
7dfJPEZmdZRY8ek7MAUg+ii+K7qtceMcAREbHSLT3KtjGhCqt5SFzDLyVAllb7dRZLwXYSXownWz
uk9FLDxWtLi2ajbCois8a1ZNDFGbQ15gcJgpflolOGJl/QxZWJ46f89cpDGQi6WxKoFJlqOb8O6I
S/kqvaCSPmfryarrA+OggNirZMZQIibSBu1INCOiTXAndM1X6CzjEblKPGrZ6GWU+gaUIx1NBOK2
kNABTLkCai4aOyrhCpei8RhFtDLfxwLLpeF/ep/SshvYsC68KCr1mwtfKXGxycHlJpMQi8QPlqu7
8KchltM5K71TYrIYlibpNqwsfPiU2ZxO6FK1PPZtq9akrBGm0WkcAcPCwJKuyLI8DxtVwLdFBtDQ
GtRcZqKNEW413VrAdC9LMNbpj9xj56juCC+5aoqEwPbZIphn4pHpbRv5Qae6P5NxQcHLDdZh3EYS
8WxgsYyGOMegFmBYUW6cPiu7UVY02zYVtr55ais695uQlhC7u7E1AIu+fDI6r+5d952J3JX4TKhW
4g5iOf3Euu+d+HJ8TlGQXrYoU52mQkYWHAhgVClgzOO25rNFzivGsUOVUp69qm+o2zm3f+VO/Kvw
WLoWVa743gklVekkmNJlgy6uclg35VjKJ1OddKudj+LVShAdD3qi1DBtyZzvSlNGhjvQFacTBmzm
6pCxv02UUdmsAERN5HjNcXRbExaxHVMLb9T0GjzWknLznZkO4Bkun7yNX2Ngezieo73Q1Kok/pUt
cx59kx1hWoI0j7pZVcViN4h81PfLGF54FobT4oldHhvLWJivhZGAGbyR/gdblpRHGe+gHoaDmyeL
dqUs6u0DBN9x0WhGgmiR/HmEjASKvhVFFiGPXo9qNPKXvTt4cBMFwOVlhgeCblclvnBxSgpFQdfZ
cRVGsE7RB59gdP2faFEGiFAppyTcnJakkG1mLAghifcL3hcRqCYWhcUrC6r4DYiL76huEumsmvs9
SaTebql1GlHYdCJtEw9lXvqF/TC/35ZN66WL90cE6iefZWZ06hAkVZgw/6uBBPgS+UPPBJXBQQRR
5nQlNSH4vMaR5UOZYY/Q8fsimPCRf40fcgtwWhc17ZqinTXvozt3ZOU8kbdXIxi97v3St5fkgC6a
YGYHEEfw84sQmrp0NkhzatMRsSAmvkmrNe9oNJPpwUnhl0aO7/fw5WHA+fVz8so7GFoDmOX4S/v5
emuGTZrHrf4L9yn0rQ3WazwJR5ecWDwfIclKeQAdQ+mZf6VVxAYea/Ri3vO986s0Rc+2q5Zc4ND8
XI9p3rgtD7E80Ns4nOcpfHxPC3g8JRAG+sZxdfHFsC2uq/OgFFMmiXN43QGL7QZX2ZZN5NoCZBvY
tYVyIPVvL4osRqOllEjZDL9TAxmwMYDDtk82zeyM3C2jMgFC/Vgpe8L+aapsHIJ2VEVnLkRbsOpt
0503D0AMMFeFXGkXKzY1/I4rRwSJAIKG8CQlceZVrH+toxGSCp5s/D4bgkkHE2RD/3/zstIvOip2
xofSdy+FXsl9rn4lEsdOnDQGlpT9lAQmkHomucg8nLNwP+YNQPkla5xeqVHjJH7etKbnLjjISdmi
TkOx94geG0fY7CsTco4OtasEtfjdIj3aEbofS/7OWepREav/clE+EXtpE041JjTZ59Ywm0zu6t9g
5EAVqRPGozzLBjzA7VNlmO3AbVpSxfJ1CS2gCAJ7xj2ym0OQYncu8iix77Ch8teqnH83enbAc3FN
Do/C8nngDnykX4tN1d40JDv2BieJapAhTzja2fUeb2jcQxGIgE++PxbVoblo5HdsAGX/284DM3Op
A5LlXxfXebGSc8r7xG6uASzWQKJyxRQiRwow5s7+KZa4UOQKapNgyhiauCtdvc9fQmSPhJjPUfw9
BWzRyyC2WEZbHgKIbaySxlJbCEx45SiKo1UjlfBcMh+1VTnAI7vDUEC4+kGQtnSedG8fI3XOFg5y
MTRazBIZNyTnXe7ddSXCx1CbYzUB2CJAuZhKEa5AzBnLwN9OKbCfhJuU7btvdtfGkrRbOyJCUZ85
DHJJUCPttbqw1aS/PtzZTxY0UqVOtog760xAidfdWIxlOd33DvjHWYCeegGkybPUObIbek0zwdKP
rfuAix84Jf+0WoiagyNWniGQ61JK5ZeA4vCblDQL6Gq4yDR8oxUbJ802O6lcxxN3xyWaABzapK+M
Hiq5DG1LK1H+1WWBk1X0fEJIlcFkICWBXXrqNOuoTcf0FG7Ua/7PaQSySoYVOmSG2kCPPjUV0UrQ
baRwyKct6n/BRSZITADKjToN0tZDBAc/IpZNxKB+CM/LxGILtA/O1HD812N+uDCZIYsznhSWshko
U7GYaHHal4ebDFlrlMapDpdHaYErre1rFgJ7Za/Us1AI2EMXCVIQ27AU98oR8Oi70jreoCb+GpRU
j1w1KtHwiqzSV6/iIMgkeZhLZ3Kdcq5Bx2p4Jk6EJXi4y3bMeDL7UxPYYIgKTmd/Ji8MAZFJ8Po2
3C3vdgEwQpm4AEx0Am58L9toY5rSflkR+EwKLssxmXt/9o3CxpvrMhhWIUD2ntxkzYPJhAXwKORK
gHHgGh21DSuhmFNmq9VYjZY4fq+NbxR9BYF5Mxe2AsdgW7eCkcAG7oPgfDbnkK1e5i4FyA4/Yig3
RXjVD3B+mNpXZd71ar78+j8M31GJ2ezh5Z7JMzzp8aRDmtgzhXFidOJ0QShga5X8k+eAVd7p22UR
czvebq5uk5NITp1t26M2dBw0O+CLIep/te1n9AP9KYftjVKQx1akYiNK8v1Y4Pm9WJQqg+Pkqzdk
SqzJWClbLVbYskME0C+nCntG7dBROw3eTJKC/LYxjuV79p6/p/uYv/fwD1OGwyQKaISiS3pfoPrh
XBi8PZ/OqgTjdfw7q+PWnFyZtcMfk6BNaL9yVpA5GShEqFlWEc1pN0jmg4mNstIsnLFC4ZPg4LUV
aJJU1M/O1/+9sQCgkcFXqx26Ne8m99LbZSOTKQ6jksvEgpB91/G10Wxhp0mWkVNB7LFvjN/aWlAh
xqeGlXdGrESUOkCfUqWm+ClucV6eFLSQq9aMODo4rAidoVsd0PAivzXzu4cPDgXUN4xBnd5/NNKA
dmPHDy0LpQnLPCm1xFByaFemlaHGoShY7i21SllNAV4XLRyYY+xxLAuVaK5zo8q0qVND+y6YUzGY
X2S6IxsDsvlzQUqQwUP4fUqpxbMg9O2qeJbLU/Q9rrr4yAlYQXxBbw6YFBeNgG4YqLHRqjFrq6wF
pdQHv1z+Usx9D1PSepdcs++Y6VE/5BjqbM1vQDUb5k0QueNBbEFWvoI3yJV4KKQNS/duV6FPcrE8
dKfsktkkHZL0EIVvzCDdZMZaj1pSpG+VsMrsAoTSRgm6sk+Zehi7VAwy/FpqovT/Ch55vZWJyeUk
i9hgCDMY750boABqL9zYdEdLK6p/bM3uolo1VnrJ+d8wHS9xPFkEkCuFfC2TY9pi6GFPpnliSvee
rLdcy+rw8lWeE4JQFzFXXBfcp37MrFKg2+2zwO4sUOhB5nlOZHVsyEaP1XMxH4OnhnxUIrKYaKPV
kt/qbgW0kX9kLUeusjBDNg2GRb5VOARcG5r7V7S20lWIFanFCq+KMEqYHAJuBsZbX3NRk57YhQr1
ddhyeRPdKhllYw/lp1BakT1hz7xl+cgA/AKGT5vwmzB2TKwThKhqZzwA71TEqx+X/UrYhLJK2Fxm
k17HQBAjJMOTQLJtQKreAxx4KwwBY4u4jwbQX+7zrkzR0WXxU8MhIRYcf5VKryc5IEwl6ygeNJqi
jkEiwG14lUVuBLkEymau44RwgOw54Y4UNpWSSsalwoBTHpm5IFyH7ksR5Kl6Z+NtmEFMO7VwQsoY
8FYLD0Q/ito7KA1CF7hEiaqdNhb7rL0ihy5x6ZaHOXti28qHfqCrbWeegtd435iw8wgHAOWysR/L
dRP5DbcOnQnZpCFbIz6ilLP5ifuvm9awl0ijrMh1ab+Uh3B/4K6lmeVd7AH7/it2n6ss/L3GzpUp
sCo0Kh/rmhtUc5SVTb9WlweeV0o1D4nLQOEPqROUaqxIFG3pHMrCsOUhlyFYMf4bQYiWQKR3QZf5
5XuD9mHA0QLGIjH2zMK357fpsxFlVbNkgoU7s5uBUENIRMR+uv8gL22HkO9mO2L9o3Ill1tRgYgB
cshMoNQoH6jXPe3Ju9OUhb77xozMvoPjoI13cdlGRp2EYeaRU1raLYWEZxIZYfZmuHo1p5x3vTTQ
z5tqW3Vd9fbE8elAT5J72Ngzv3g0v+omN8oASakDsepoA6w8MteeAK2VqJqmQ6ULW87hiqbHQ/2U
CddK1HNyNCUBTeFeRsqSt0IRV5VL9zy5u+Sh2H1LAT16/Q2T8djw2cLNZSWsv8GeJKBgFcXgtjrA
rjo89LgV/KDoxlEofIjAHJtSTeOH2qb+Q2xBIipQVF8NlEYQ9AfZa7rtsMSVQUpcdATTKvUzv+QT
9SSiX4Ri22r8vfqJSfZeviEnvkc/0lqHTWc5iZkz3+F+BIE06+l9TXKeOt61ZyX7pl/3KMQlvL5C
f0WbBj7kKvOX6uUebhMuEWj7dI1+RGxo9ax0+Z8L+O4c71RNKFzNaHl+EK6mf+AtJOl2Q0OYCAKT
B9movC+MEKuuGUsRnf8SA0u2IOa4h08DVSieCjMteMnPNNZwJQSJVD0PBWd9zQ3N2fsPC9Fa8mrx
Zk3A4lb/3pIXQlG4uniVRThP/ML5ehMQHG6Nzw4QStpaU8sdGlsvO/RcgZt4+SrDQfU7+cHskga1
FljRFPFw6YTi/a8lVrdSkfPjCdubFPBgW5sFQn/0sOIlkCJtMf/Lq+8KJmkgWysunJC5GcOEaQUT
pXll6l8caMIEGRH5338gqdGFee9ZuUqUGKQ95jbmrYVxiYk5VsJ1JZ88J881RgaFr5G69d6QfDp+
Q+cyEWPgrDCyQAHy7Vgb0kqHwxYTapdZJauct0wyPbEH3SgW2All9AbigqmXXu8c5fZG8CCmfbX2
MNam7m5SpstksStE6x0xxOrO5/c/Ck9BMKHafE2SOx/lrojZTM7VcYYv5/KqWFykY3yJSum29V5K
+g5PC97bLJXXYf3IXR5/iQfch8UswUUz4JYmqE0IJazCjpQSBjg4coE2tdtV8QGhmvS9B9IV1KHm
c8KNeb0oAQWJD5wGJv4ge47CrAZyo1NkQ4lI+nwdoQZwEr174wFtS79ph8MIT3A5jaVKUbXJGPj6
bgvj+epxEsg3IR1LteKAVJVIrmcV3p9rJer0A+7Ev9nsSJz86VKQAp0m0xSfqO3z+BfEW7mOKLu9
sUVYW27KX9izikaL/GYb+RlpZWOxnX48WcL9Q44pcdhDr5QjAILEacUKvbAyD2P/v11GKYMpYLeE
qBvtPodDfREFY3O7JNYxSwMmUI7EHvir5VogGFcICAF+boUo80+ojeNlXwHAaVM8Zq0KMP3ZaFlH
S6JIINoaRYYf9ELBXpdD1iuzsfMb5EQzcy75dctC6UF6XCyvMq9j0nFSQaDdR7LfBXBWEnhmoOfJ
H6r+vYcCjXS+aQkhosg/0Hj7ANJRWSqYTmCeIAoAmW7804eek8754pHvNAwnQ605gMZXAAc+Tvbg
SUSvptP4O8XYQm9+jiKC7bkhWaADVVNgdDQ+xeVkRwyXr2LyCout0BDP6sYFAnFzORv6Hugr0xUD
BKEo6idAk2o510qzzWrzG4UWTcDmeld/mgRjN76lnksmkjDevtcGOK1K4A+FDFHOUN3AM7pypqtw
CRBAzuTfFjNBQ/OphOJnVaAATF3ZkOhDHcsQ1rtszlCwTbmqRUFwHF3yD9HvDnY4onruGO/TCa1X
SMT5UlhnE7vkhwb1w+RHGfEIw6C/b8c1F0PLj5/yNzili4pIv2pz5lorpdXfSFY0NzmkMECN5nL9
TLPyX19vcjEARGO50n2xZiDJ85wdX+xt2EwEUsvOXic+yDM+9m+tBrSd+qHUjoDLSW6MZrpO+vqa
6dV1ZKbASVDSBpYtZNjDQpWd5J7qUd2kQNCR4nfpeNSsRFtTHhrHJumyBSfWj8QkdxRa9dkDSRsE
nPODt63pVZ3Es0+wInC9bhIY5Tm4cPiKIFmHRGZhaEV0KmZWRlShAvCx3ZEi1LZIl5ebfZ79FgtF
qGTklAZ8MqW9a1nFELnS23bLLpqWnGFVhQUn+umvdTDy63D6VL14p46/fsWclJMR37E/iWn9jcmc
vCO0RiGdLDp0DYHFa+nGmCH6tqz/geHSwCHQ59nBBbMaTn6nf0bx6SVVxq+odd1I8Hp0Ycs65CbN
wF8KB9gp0WBroAbFT4b/j/pEAiJPmVuj6bLfCVRuADPF4r8z1YqeYPDseKdzT7Ns0KplgAASwcIX
UQFX7rdJICk+jl1QCaH6t+CbY3+CkeViKrPqqZOE4fRzCYXONq77bwAQ4SMAVNhJ4Z+N22Vs7rDL
cbENKimWCBkYYSFg4Qy5oUz8/xDlrPBjKlL0AZeSZGOttYOB4tfnw74cjtEda/MfdtYwwKHH3QsT
MKgPiCNJ3gI/0C8+lIs6mDmyHLhEW9RrJeWvZ7qYd2wbIlMz7cTYmPrBu7ZCtVjBGEnkk4uCk2jN
smVfMOLoX7LReOoEL41e2LEvgV7dW3mn6a5y9Z0P6E2jjajbUbliftn8IafOJgBSKglT3Fx9Kx1m
HqjbQyfyIOv4VOhskWdtz76wdNz2qPUzTpV8tHzbf01SY0AkkjIywVTcTKsy92DIW2Q79YN58ynj
vDQBVwjZbVKypwMavgOCViVEEsOJMGqVUh4AfGB1xnytyOhcP0qBIhNEHsfryOS9Xz8YtbB52pZH
+01KVdl1ovy0E8Q/Y4lSII1rZBK+ku05BcnG+xLyO5S4KbEaF0dbkfJIFXIPL7NHTs0j87o1ZHjB
6NfntZLuxg5RLo1Igg/ffPEjt+3EOWMf6WIgMhTH3LFRMn8G9Vmz4bpZL/n2rQfX3AhPPDaEOhzk
I2C5ewvL7vPaW/rPZN0Y0XdNzSwT/7PXKUGap/H8SP8DjL85tselr+Iqvlq4KtIAcRyDsuSLtxFt
OeD3jDyjckIDlz2i0zKiywA0a7w8r9+C9tA5YKPdzDRZnazNE6Nzh18CHG6UfK/FKaqJMzg2wJzb
Nhlw0KFicHRR5HVVFS4K4ApVrBiVCgWVl5CGQwj+KUFF1uw7lgdWGtsFQXIljbaFfmkVfSLtVXNI
gYNMvqhbNTruuj4q6HI0jhC6sRMrRy51c0JY5chW7gQvB1gHmAgYGNQ4nda8SF2NXrQ9kLrlxVIp
8NLLN2SNYEglPs9lRsQuqSFR3wLH1z5nASFhXJ5Qh+YNzR+UJpla2jcfnQ6490zz9jga3V9VOtW8
tInO52X1JHFCT9T3y1lHpQojvvXQiYwhFeql0RY8A73Gd6jRO3ERwEk33lyQQNzuK2OInGT+ETaT
iF7ysmql0ZqhrybtfHpeHhcESpHELup7NYPB4MB5z0CMYG7K2oZV7WNcgQIzOqefhR4ZYWERjBt9
gT/0eppprYrcg8playyPxfL8YI7PCMUNJCkv+3EmFgaMA9NgmXKLO0fEf3GS0mY3g4w5z2A0R407
cOW01tIApOcaaIi1evkIxelXLlQlSWd9Ab1ThYiepz5stEkxugLxpR2DtUxarB8ThfeKiu+L8RLT
zdN3sACs0PQ3erGwf+fvZfR+6lrq9PY1gUOccmg3iNFWQnXqJk4/cRjxuXzHOfIaW1RlpsPykB8+
jXZ51dxJ7Qn0Ia8Bds3Qma6r2dwkQ7SmZ/7HZcCuVr0Utq8GZNHWLje58nDeJIs2VbEEQGYTRP0m
zIkSVHt84jUVgMRpX8TwN2ubmTowJp/fM1ebii+0aMlnSCcbcKuL8DFU2aZoeLcjJsEPntluGNOT
12hGtcfwNFnt8nih8yQy5F/16xJ7BDRtD1/Y5sYgw9uftgA2HIgJbtRinBd2XLM86oNgH2DSY7ap
ElTgHTPlpAnxlObidaM+Q2MJsrm2RHnhKOXgleey1WGvMiL6w7BFb5X8d33MH+L6wZk0wHhPQ9yU
/cV+Eca4FRnKZ9AursOL8OvsHd5JVHSjct7HapcwJ/3tZ5eu/xaLIcu6FAfVtgR4HPCsLH4BP+LM
O8bcLVJuXwTHNofRWrLvn6lHHSRPmdMPTeS9+2DQokP8HyviM4ixPE9DcHpLq4X0tbr+58pRrOwf
IJit5CLd0RZcVPR5mDDX75rWjElChQ8e/fE0RUbOn13PM3kvDu1AJHCRsP0SULR5/lOe8azDt3vN
ARbyY2Oic5yG7TZEC615UR1RHx4NXY23RATR7Kxk5lMc3aCLIEVeSmKjgIQyo9N2ooFzNE9g77PY
niJ9EokIOu414qlt9vGQUjWuG1Bj+rE80wT9YEJQ+/ty509HpaVXcq0QQ/mbro+MD17o9I1ppvP1
W82JLZQVYRpQShj+CAafxHiWaOsCm6a26qXh4UnIVg0TDqXSu2t/ueiHenBvh4Vvzjc4vRjfvNzA
JYWT8UGPYi9ogi7EnfNDElVqYeYarjGhLpLt7LrXK+aHHR67NbyTNptS2QD4jNHFcOdjtSJO6a1c
wiZ3ACJWKfUfaa9q4C1+TqMn6778R5c0KHtH3OgfoWlvHvxdmJ/TFYnQgTVbNd3AZYTORFKZQDg0
WIT3855gx2XfCJkE4ecHNO+EJpmispyAqm5Sf4tbzpj0mpr0ZVpYQTwo0FLdFBkkvhxYeJboLWcD
3UeZiLjndqg5UTPcO3OIto0ncDdvB6RqHMy0OXcVXgKLZR8mnRB9/0ire6GyXwIbduo1TQ0m7Du9
v9vbbvbsZHUOgVLJ6XUjlWJrSEbAmn+YwMBpj9FH8jZr55lptG3LoTXkwmVqJkpDnDMHBKi9BOMJ
3CGXesgX+61/CVb2yueMlRgIrb/+1kGLSYXl2UeD7esLNLUZzoSq1sUdE5dmgdaDYsKW9Uq2P8VT
zlmSfsW7sRyl7WlTiVnhrAo67lRLDdg/29C45efYtjKG0L/08zbbQbsM7pdSS+FI7mYEY8TyCGMS
JeV9sFdXi6VsS5lOcW19crgmbyXCynB/MXuTdL1NCr0SzCqTiM3DQ0WvKr0Ipaaee1Ybj4I4hEX2
75QsIj25ylGvYguFssnqBZcH+gW//NZVZt2YzXyk3rT6OhiwMysYdU++wY7crJHZeLC5IN+nFQWm
uehXBHBdS1qvYFEpvEwe1kIhyt1tg+NEUEdE2gaY9lSN3owF7g+L4Df0U+gyof86mIlIpnI+IIHM
3lUC+yd+eH+Rs0BN3ePoXD6TfKJQblRjwXEPPF9C30MvNp4uN5dU3QYWvQ503GM1OLI8YJZoGiSv
LAFnD/VGO2tz0U/3w+rQ7SN87Ywy9nDAyY1EvFK0RTTnhycupWQD93DsMql3mL8dEHnxE1C+0DOB
lbRW5+8bDQ+40c4SVTCrS1Nh0X8t994ForGDHpc3CWOXRXuCxxCBFQMKfWmmPctgRo3tbEGi4/ZD
6erxWjzpmsb0QZpWNBrgIwOhDJWWMuifuRl9yZ1uglFiQs3gdfObJcmwhPy1yHaOobmsBp/17sGY
8PF5e4uUkzbtzmzgfpjXBhHR7A0iFV5J4luiw3BjznTn2+CoGD675U9C3H0sLxDm9DeG3QyedqHJ
kbPI7OtCf9EGFfkDvHEZdmaN53wKQdB+9fOfRMGVwJTvOqPrILrWFS3cmGkPwDUBz/nyRlDmHCd4
lnE0KrlNZspl/NojybEKmTC2t1lRAUXL7TpzRHqwEHA8lTLeM4xQyE0OtPAvM6Pp5U13Huu8Bs9l
Yh7WXRq+ggd5DayB+druoyvA1LyZUtZ7n84x8354X7n3a7kEQHtmQB3WdBbTLa74IOY21eB1mux9
iyP6OOZRfeK+FcBaxWHS3LzKnp60ur+nymK7cyteBLS8JSZhwurirUlDWqI+L9YJ3la10XqjcjQ3
zkK84CyynbBeYg4WNYssPoL0FJWOgPnoNXDYeoplVwrOf3+7uXoY2w3HrxM7eoHNSh4mJBVyTjko
IwM/OokWKpZpmF8vwxRv/xSQqDuV02bYVCKCXL7AEvnHUVXks76aVXfobZy9J3h13xyWu3w+UysY
8+ub8JyKfHpmAP6WXZwYj+fLY1w7Ya6EoNK+K1wh2MrDmgaKg3lh1y36RdDFRAL8KeT8/Uv255hi
1rltIt5JAG190NxwUQv0CJv+zu1ym6GXodbaSLvcGKYnGFjfU1JtkhhwizoaRPF7nAvzlSTvW9nT
g1yXlQniruJTuJqxy7Glslb/9smga+RmuOeuhXZeemUgGPH1nrG5X+FQ6ZLXmk7PfeOklCdtYnC5
7dSByrCdk9P9QtfkGqG4jo3FlDWKE8lr3nHyoa70IZMWeAnTEGwbIRtoW3clfaExQvGeTQ5HaLag
uFKn8t1oTHSkCop2BaX/ZPDkR9SOn3S9dbI1N2RmPhfUHooyLhc83N8aVDe2zvQli0hT4KCcA7Pz
WMIMNoKgxe0Vem+15WSSPgkQmop5ueYWHC20eXRPiAhc/uAaGwUYnZbba0GTt0zrCoLor/A1s7OO
Q8JKGM2Puo8pwG+aZP0Cukft3rHQr3hkqmcBvdXRBAX0xlFakyHjA7JoiH+NPAZndSI8/ImHKW1Y
GsRI364sdYg3b+U5zHZVPL/iVck0fK+L2D309TzNKsNWoMdVfLekLnNc3c1OdqIBwL/k4lVwT/vj
Ji1aaZxuMUPJRXgetZtyYMyh+Vv216mYwqZgycUBR4DKqSyoLqpPsQDAMHgL3SQBpQd7v8pG/eFx
tE/4SuZ/xoICYsiVlsQBkBdQPf++ag6eccLwbWPw4xjuz/SbzWr4ZtC8/S6wYgOIH83nK1l3nMGF
+SPY63rsd6BKkjdIUksoiazfwthdXijLfOQVXo+yD6TF/7A86EjGsRCWlwk2iUFPHgrkMhBIF5Ku
qJ1mW6wB8rmrMAhm3igBFkdWYvhbjx4l5zMSLXMCGqWbPpAFth8ZkdMhs+OKoFju6XrPKPp7EZzT
ztQ3Pdt6MuQnWP0xCA8fb4Vp1RT5ttO/1myUp+aYxsHLIdPYr/hGr2M1UCBZe3vqhdvp22+oFkTQ
p9/avwubW+eVJ4NUCA8tdczdrndbTuxvKs2I0RlX6i1Y2aOQiC3ehmDXWf7R6Xqj/5jfEvd2QWJX
cHVAFFt1U4TU7hiUlOJWANOAvCEysTh56RWdGya7TBmc/xSPqVr5bg7mQHDUFIL7O7vVzzMfJr+P
tt+uYGZ50Tr/rC3I2Hyw7Se5uqCHRfyrAwOuoH6xUPGVJg+2KtGbyN7AVqYlivzUQXYU6+CqdCAg
aPhlnthKfNNFcPVKqsdOD+HOo5Y+O5J+XtBVXL8tg76BolMgzm7tVpku6Vzw7PgHJj3H4p0wf0z8
Djurst3B3YU9mUEu7547LXtiLPSIsUW7bAjF4x6uaN7U4DR6jcNW9oTEc0mqmWHZsjziiZNhbHQX
E5QUjTk2TJgtgJyHsvx9MlYLrv1d+A6yhdojyHwbJjEmKBvjLTWc/PqZ20EI0tcWhNMdwmvaDMCl
Z1f68lYPqipcM8ByiP8/KRiR/AXAI11w7xWBw3T6OXEwX5+2eHznTVQPoDTh+DxBSSMaLTrYMimV
wf4Uv3S1TLpcTLgI+vxi36a/+o9rVWTbjTGYgT0Yr5uVjQ3OXhSha26xCns7Dz0xfB7MzWtE/YPl
AmV4gkRv4dyJ/lLGFJ2c4q1Erkyzqqo+EWTwGPr16NB620SffdU56NsYtlSIWOKEaOq5kS2SrwFm
sYdi3uhMs9UpNaZa9vcqk9zi22kshYt4yHA6Bnd+VnT18dXGmGhPnGU8eOj8Wh8naio6/Da2e95u
ReM1dZcPRrwOcbbeF5hVWrabypMS1buuW44xxDDkdFwkNhZyfwHavV19Yhjs4NetSR91QADjmgJz
xSrJBGiRpuVC7NQAVdMUGrMLgEVT+U7l2+I/c4cfWrzPOmoLaVFBxtjOmJ7ELGBASlLfdDtXSyg9
gB6kpRVJbptUGlIVwWAP/EmozVCTW92qx29r2VPjIXkWc1z9Id3QO5F5TcG/qGVLxdvIokEsSUm7
LN37KSvpv+JrGhw/RRlsmAFRSO8XmWkPgC+7OXhv2zShxZ0xlYdWa6kZxr3HjaUlGj0Dg6asT8Bs
l/q37oCbt9O2I3YO1Yrz+muKuCU7JdAR5pv3dG/fOZwaf0HNtFJMeeEDh+ulXIrbL1Vhve269VI+
RwfYiPPNsMcG1G0/jd1aj3dn+9u4j9AhxDuWcETExBmDg5wjjq+wVaKROXShW4ExhKICrnwoIUyF
j3lRAg75Vwgq9OfsHdt0EWiC149nkbDtjCxKmBHbaPbOj2eJkZmPWHrwgrRgxuiqLHHVW2IGtI6o
31r3Emq+ub5BUpCA3zpzru/ruGdC6QeeuRkcbZ1KSDbF4H6B6zCeiujzNNZCXlsHN41ENkVd8ec7
gcrkefbiKzU9J9vNFEZnDdZkDLFv+BQzvhHNLfj40XJbkoWm4gIHZ+E/hZLuQ4f5y5M+xDKOCXnW
lEvCwY2VjHkLSuozrnDIIYFuKf1atm+hVjfg8IUVDT4r/Ng+l7oXkQt6FCm97ruXgvkHTrMPeX0/
UPP03JwGZaTIsTFtlxWejIau0vrX6kV+mptikOyMzEidLhwKDHhrEj/d33V6SEtt4hmiHKDTwLHI
g4iFQiQe2SDXDWfRK4ek75MdxuNjo6ZRxX3xtyq28xMk/22iozWPJ9CYtBC7m1cCxMy7OGyHlSzu
/VIKshDJCwTkSEH034O06ikH3iFHQi8ME2+C4xYLbb2kPHV6fD/8iHAJLSGHbo+6w4uruTJMJ2Gq
S8Flxw3KHP37UA3Jh8Euzs1b0pWsuNdPontlFGX1etGJufARzGHUBb+i+bQj1pTsD6ctNNh5hrtm
2k+XAEUcHrCFY1DGi5Vy3oczR96GupGakA1tZ5eCyaAPex89FqH2e50De/GBMlZ7x/cgECNK2vMj
cbHztTW1gDKpETRcqIrpAXcjV1ensCUiJXPbYMLh3Yj5aj22jdDnqmHspayL4OKARDFyQVJMtLWz
MnTo3skCklry2Fw5lzzAMe6vV5qLsLSoOgQXQmp0ffZjElLFv3nFEodssLTV8tYKYlPU6S9aJA5p
pB8m3wC76Obn4Pm4KEXwmR4NnIoiPMm3Qs1gyN4tAjnh/Om6Q47Cm7mohHArpuCw/ZDxdyuk7XY/
SJF+3WvvBNiUAFxwAo2k4+eZ/0urGHEqbjn0v3ECKpTFbTdU4dyjB4ENmBxB/RPbmInQWtdLp8KH
XssC8+b8B9VbXGM5B2QXQx4ROhqsuu31X1ZOpImSkxF8y3SJvcfxDHN/knjmoIWdTQjg3N+tXSnR
YRin7mf7Ww2FEgwqXjXc9LrwF5hNJOpbulG/vCkZCl9x6ZhVIXSRXROwTq59oBo0ZrDfzzJTg4TT
U4Qpm999hpMg8hBrLcx5VNRbpI/YBwbQzLb1ITl8tbGY2xgDFYRaXWdzd8kgaAIWcJXtWyTWVtsp
ssG3EtHRsGAGh6RMkp5rrmVqVRL1ohvxK0ZYiZ1hyteFXRlAtB8A7SfIkDjs7EuK2h2HfsS+CHYc
o5+XqeVd1y+r3vZmmYcfgsJYCkM9bEh2kx7XlbcGR4xEj2wsd1KmpG57QwgJ/vjWe8WcNNRN1tB+
6h71BZqA+iZOReMBDWtw3AJLgjDWge8YOrTFXu5tXh9uvvXECwjR9wDd3hoEIgPoJ1gUFFrQXfkF
LNxWYj4ZlrxHTSg9oJhoKIe7j9UDCFq+4kYnVyMpW476d1884/CBKSnJoAtusByGZ3ThBcwVxXtJ
FtqfCTBNBrLZQ4F+goLZTx1kCaOetGxPJYzw6hrhreObJ99RCw6QOmxLucayJSmX933yfZBMxpBT
ddKDNZeJoEAUgn/pAFkMzM6zYuyAPAieWRvFbSZ7kh0mmMMyrZdlq0SG5Yw6KEb9MkXduBbcXTIE
w7/Qv+40JWoc1B/BVdW1kUXUv0FSwk6Mx7RSOeWSz+oa2FrZWDvsr5PZiTjqqVu1Bz/G5U45+Oio
uHE2pR/ecoT4rnYnUGK20e4iBp5hYiGGy9yrY9q9W3O+8SGjMiVoT3k8vw2+7ihTjdakDyI/UBu0
xnw8O0WPhKWQuB6C5wxsHi0mjHBITr1YSVQ3WGXk5FCz+bdptNy1aN65Ue8MRYIBxgkbXuuO+5Om
O41c3TqR/3ITQQDpLQNnckluDT6J8e6TBmFfIqusmD1/3cvkB+4bEPea9apnuCOTUho/mbwUbbbC
iMXn01FRRQfwaWrNiFsUXM+CL4pkCAYoVDv4j5uGsOzp08ns5N3bP45X1RULRaWOM+ZJYUty3XOw
uftv+3ts2Mm/1uM4sFUjaeT+UDYbOuuKU4WNAS9OR88UNjXMH2IhPPLeklWT04XOh83TMiKyyf2N
U5WKismqzHmZD+aChBESN+ZLkFQruD728ugP8aLoK51Oc1b8NTs0oPErMuawqlkJ9W7+IuNJKz/3
OnR+CcnA2gTbVhCJScZSsheXgMc+zVpOHa94pbvhHRRSvl+O+5s+GUUwBOQK9wFld7Cq1JCBad7c
OS36okXitokhTGKTivJyQvCI02UD+8ef2buoHwwMJ5dAVg3ZIh8tev/P4MlpN82MwDXU4FivE0Lu
l0E6q+3Ak6yTusDQuR6/8DK/rKecnLYk9pQCS/4OZmyMUuB3f4CTLS2u7T6UjDP2xKagNGFYgP77
vbgmDbHC8lXsMwHs6nCRYaYHPuVNyUAySiequGW4ScLEtYgesYrjWTWILlAi755X3a3FrX0yqc1N
slcOlXYk8vpUwOHNAD7RI0ndfTjuYw9j4FeEmLYgy67XNPxy8OKMg8fFeXt2t+Z5Fql9pjyisg7G
exUlfn3TJNyfAV0y0Y/i0U20S7p7f7AywLqCaMp5z5FaoIz26UlmJTYMyv/9Ye8UfR/wfm2at5G4
k/RCWkTG7ib3YsG+PSE1r1P/D7OoulRJvT18CcXB6HcmGYjntfmDqMOtL/DqQ9KFo1t5vnuj7SvB
x/WN9Jjr4y95FEx3ZuJkSClUg+5chgC9wCngcNTLuTqgIoACbZ8Cesh+D8ErrCtXdDIgbhv8hQTA
vGwXEqFjrfyfwaMf23OhSxb/dNaNmFXITt6Sf4tSjMVcApYdWkaYyGj2sGxchqacIWj8/HW8iKFV
4e0QnwxUXuZ5MOeEoRjLoSYQWBTVn+1RuRVASdjk4SSDr5rD89eKGQSS9L7ffBJo18H5r80BHWtO
xeeT5qpBg4AJY+sY+vpVVyDnAP21MNREuaWEzbATeD+nIHFu3C+Wcw9vYsp6quILtXmFIUQR5xQH
dH+yzGmdkjJhTLqnIEJ+DMnUcevGsjw45leCk4cmgcvvvhwBBCYM9WlQR6rxH86lLHjkJu/4b9Tl
VUPFEtz3CNLhdmcNu8Qx/X3DJF4o9hAloveMOWWyMv9HBc5UbEV7kF7TEpCiJCXWdMqXrw3REwot
a8h5X2x9SGRYl40zMfHxFBgvRYFp3cFYlxzEgpOvLIt83FH4SqHqiAnYIr9rDefxsRRlE2Y1EucR
wj8UXNi0NfG1tQF+Cc3224BwPkmILUAVVtPBMgmC9E9X/FVFPi/j3AauOvyMKponA2QJ+XBn1vxa
oUAuEjR/Xc7Dq9xyZs6JVINK55D7uJiipCmtEwTQUg+M1ijuBKn/40M55vgdWf1jzK2StOzITHyr
KhUrkkfh/LyNP67fM2PjuTeobMwwBIaR63zVk6xSvrSbFsPdUZkVdhEfzKxdyAaSookJnxTjjFsy
2cXxMOxnTphFhNj+Tj5k0P/sNyaP7XKGdGlkgH/jyFB5VyU6MZTupSt00K98LSXX2603zT6de7FW
66xORYNFLRGLnUO92PQqai0xTcR/MPCXUa0cr5ok5XmXPINtH7JlWFaQ9LkElbzpTx9c0X4okqiF
LZ7ZmlvO5blwpwH7h7l1UT7hO6H/dNjiTliq6HjqrLOfWiVKg0v++cIoArRuQPWMvj36daSOTrI1
CvDIKSg6Vl1Q4QPrQ6/W2RQKqm8OxMCt0IPhM3WYfgMcAdNckIy+ZjZo+pIUy8LD347QZCc6Iue0
Qc3TuaFCuE/fQycWONMkN5PJLvnJYyWNO1QLvE2aXO/FFrchzEYouLhIOJDxtCqAARk7X1s9nzDt
EQJMCVVT+yy7x9aSs/13OCM9PYGyt/BbLFHxgvUJCrhomMdvbUz0cTHh1t0jg9fpkeaPiBCx4yTO
0CD/vefT1ZmLmnNRdHetPf2ZpkXLwMdRM1nC0Gz8FjjVt/30vJuzeq2V0BJjtrOMR5xkJGWzgQz4
Lf1sa2Ub2QXoxum0Mmg4RjfP0SBtS6FMG+A8prmOpfYHHIJPO48s7520YXzF0OlAMqDHauyKDLPW
h9fq9z7kiGil5C1TqhbsJE6RwRvhaZ8uDq31VaMuBKpdPFQrKbTDQeyi5r4eWQpnyF+MtleXIEsO
As4JzqrL7LLfhRpEFeBCHf6xiSO88e6imQwucqfBG37eNBXmgFL8XnXfeYf25EghbmOel2Sfbo1J
kXxVFUxtIEr+Hznz0kVRurnjL1sF31yPgu5AVAGmNDHvEnv9/jwROr0SPc8nhijgVO5XYqVfzL7h
95wpxq4qBLaIDX9l/f/2Vx0puI6Viy197nKZ58qwnk8UTY6MuevckvXdwj92/DsL4D1G2dZ1lt4i
bFpytRVeZm/vSTLVaaXKtECCJXmZXAE1SIHrX5E6ukXtDiYvbLcPeQT0dne/TkFdLjyNRGI4syEZ
iU2FfZ88EIUggw/QJ/jo2ylCMKCqsaTBv8zR6WHcXRw4Z0rs4lxWyviqSUgh2saEcaQtTDppKQDq
qRsu
`protect end_protected
