`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CcAMH4oQ9L9dkuCdix+j7SFW4CpnruvkJP5It3NlYG+eSSas5+bEKdWix8xLT/RLUlAfaUNkuuvx
UxUDFfYyxA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ET+/xWkqvQWHLsnBJkHC72RZR321bgQYThABwXQpdzM/8ftwsWY1TZ4xB4XYKEX9BBd8DcptDWZg
2ZGAL99y7UVjg2XNdl5/kMcVMOPnCFavB2dyDwkzqqqZNILgPWYHarFSZvUwf/z7Lo0Qr1AMt0am
/Oz1Nzr/19rGwPyjXm4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MH/3nBoBkra7x4a6gIq2yRpIV1mjTv0nSXt4rI1uO1pqiihI94Yuv9KPadoPMmrUhm+w41I+Eao3
gvjTmT7XVO1delv5OjxgA++lhHx/dCAxqIkDJ5E4vdfp6ToJ13xEpr7MCL0NKyex673tecYCLGKm
LOn5JJXVyluSdye06Oe2NJS3BLb+RUSDwyo3zLT4cbLOBnoqoRpzpZ8qFF2PXV1A2chAC8aEJjDs
jrM05EO5xDgSrZSZ/uonbhW+VLkydGud5kaOY1+PcDsXxc2VvLlday/OdLdUi44Ztfwu4iQGZD11
3+W0Y3abDuLLZRsJzdwl83nJMzDB6cxxTZt9hw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eYaadlELTritbuhf/x1FPmgBbZBW2AvUZC7YJCyrUTgsm1PmjgdK74S7cPyhBpFaJrFSKYbVQACA
fD/OOsP1OpvYPghcV6kOnYuBxPsUFoOIB3BmRoxajPWg5QMfJufrPvczN+6ddTximuRxkZnw4cbf
+a3QKUPBPNPFtAHamXM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tUNqVsW1K+T8k/TrWXD0CHJ4rozJ4YQbApBjqq7K5i0NeVBXmi9jDpYA7tJrqAGYlhSF9tuNXIGq
PI0AKeDh4DkIfTSEpFm5WE4bB1dRk8q3NNNT5BkwuuXk2cYUfC2NKB7bkF3ZfinzuAxkxjnx6Hm+
yjp7J11NUIqBz7FMOKwAT/zttWEpVvGrMrMWSTKOAI3YqXc5Mu+TYeh2CyCJ9pudPjlBcaF8vLX0
noIaJDFoEzjfZwEoj2EqDNRryRRlPQydTHpkR7XKkqGc9eNvCkUZoujKHDPnreRugzkEb7X1ORzd
GUxCmPz1qg/W2Q8iMjsscbvFHp+gkf1BznkCuQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25088)
`protect data_block
4pFAVQ1fHuss+y4DGnrUDhM14MF78WMLELy6WCmWEsjwBntOlMZd9NlBegoXXUBXZf+/5F1v9qXb
TrVFfLuQ6TqWrki7qPCFtwPXuEUREYkzITBa+H/T9eC9mhy3hOFpvnMcRuIXSvM4iGjUbiqRYi+r
TX1FJAvb6VqQf2XiRnsMBs7FFu/kzDDkoBIpo7+E9kqJDfGVujPXsxwFx4g6sWjavY/vQDKfJigl
txgeIHSoCJpy0dob8tBTMspKD1USMioGv9E8o+Pp3wxwWHuiySME6QmICkeUug2SpHWTu7epchti
zVVenZmMMeq/nuEMNWvyQuM7In0Ftyi1Vb7qJ1dO5IW6AAYD7/JrQYHx++KnoKzLOB10X7IDA+bn
8L8QNKY810/7A+4FQDkeDaTP2ah4Z4OZ0IPcsC7gyS+v7knjFv1RqCm3aMd7eIaVM62mw/FL+zGq
mci3RAtstG2ugKRP5DZCan6p2I0SoD3WQ8PlD0LMTVMpb8QM6eCDDlwAgZ3rd4DnPC/zrkRC6WIW
CQMnwPubewDXil46BFFLEEOOgvq0l/cNNqSeTImaJ5kSYsTgUWQ6nhStAZZZEMukDGmB51R1Mowb
1Rz5gENbJjlSTuY/QIhaSHV+4DxaXP2ea/bcnZtXN+IDN899qcuHKA4zvUGQ6s+gMyI1Tv+gY59k
1/u2ltVbv2FTUG/1KgUFFgVr3+aJbAGgxHOxnQgcNbvJbaMtBPPoxzVtBe1nMdiR6kPxR++5tw2J
OqSUZLqP7e0A1FyX+FiUo3jWI4bb3/YNTII+1Emp8dd5KgjR8CDAeuE/jLWWqqfaE81t8CBWD/OV
vEmtt50qeZNHAWT5FnirPo+i/PzDb4aQdCOpqoLKBGppdjTqcL/2HnUiCI90cyt+0CubysPmv71w
CkTuu+JdfqVtcqDcVQU0ZSaDpH6ykFQ1ufr6X7SHOFRbVuDn8X7oH6T3xDMqaFzI4Xp0aGPBYsgZ
bzHVBhH+6j9nwZG4C5RzEcjOx4c72mi5FddZux4Q6JWJhsEqcGYrfLYyR40w0t5ynXpt3lSImcR9
KdGyreUbyZYjUU/c8XvkMc7rPPfa6BKC5dVc0/E4PxHAlIlYkKG9IIbCPB6QPQX4QZkztXHN84OB
IYoxCtpHyyFO+WC+AOHHv0628no7Ffc/NOJuvFQQqUMprwaVDME/u4Pm120FHYU/0whn0vTSSyJy
pEhUSlOiaSi7l3obbJfdAesLlqfr8j+tAlWjH6KCzMJQdIs0cv1/5ZxA2o0TslWgrBbuJeJBvluT
9EFfs4gm3WSmeIP+5N8xp5/poPRAh8+CreQb0PKsJ3/nXFM25Uu9OT9Rv9f8LPvtjHeBBgq00fBS
zzuf6hiR6kbh0+uPG4uaO1yS87cYTvkKtnLKbcl7kItAjltIgBsoKcBk3thfX4efaRNzA04ZruOi
39A3+8y0CGQ3QI2o9BeoHWEL7hVBqdjEu+kyX09JAa/0k5q/pQ4RAFl05kVMAIfX5oNFBURq3ej7
zqum/qjqJNAwFmfJZkQMrOYD2hdjPkRfq/drMR6f2H1WeV1RHLg1C7OTtR+zcKtu6EoStbQl2lzG
1XcHrRqQ/RSe2xYM+YwkKph4FG3mUyXBZFuwVJ2EEdaJQzMFomzZABy2G2f+Lm7R0fy9vvoYsIsk
mU4vfiysrZV06AXnWf8mxoxhhYg33IAXie/Y62z4zBMczW1kUAiWd1tf7jsJgTh04e8kmxEjefVs
QK5YTDoduEylwPnmBuOrr8g9nmXUJ8wATeejlVFcFjoG5Vj2us5u/OTo8JOwALV4fz43FbsLdYr1
+9o1JxVKrSrwb9IO6/cpC2LAOwYnoWz7cMOQGruAHH9U8Kldeo7BVV4CKtjpK9adAn4ohU5rrFVP
YbTHFO3120Rr+LaPoNtYLSPlFC5th9vGiGRsn3yF6ZB7VbYfXEjVf/ZCtdlzkrwYcrhkc/HANsCD
d3kiN/C2om2vPbhWZiDQA/B6+7XDXbSZxFVh4wIdCUfTe5ESKYoRh6LLrgN7B9TwT1h1Kfqw8mCC
O+3m6eI79XXhbSdCLQbCTpz8zsQkNh7mfE2UsCnQZbjZeSVqfmU83d3rgtiV9+Lxpy0tAIuflp8J
Iyv/89h4IvXpyMOfWFJ5T+QYiG47Md1RzAm0TQl+pCsiSxUh9TWMC5V3aULU89HD+3r1sLkUzCJc
tUoZdhzuIpNxBchxyHZY+onfbokDu3BMXEzWRWCVgP0IHGVrwUcX0oL0plqUdS5Xwf2A+XMVVKES
Jdd4Jb3YbcJhchqyuITFA2set65oa6ekkOCxXjOdKLJwS21lpYzDelUnEdSHnl+YgD3vOIY4jxcU
2EibNAedH71yXQab9K7aztXVp7DHXeZ4twtPQjo358eeY6CEicDMkFtkSE0IdR/J6bLWIKaANvYQ
MySYp0xChRfyH8fR1L5oD9x67/QbvatWxSdZoYwE97/exA/Q7MJYvL9oDBT5izmiJdINmLSdKRiJ
OHl0wbC15yb58T6judDvYZ3niShpkCpq8McUUCTJxHsXBNV+gzIgOrCDIN+OZRDGy92j5ICehf9x
fEFGnIX6URCjoP506EyPEWzAVgWSXdMx1+nnqf4ifNcKO7XAtmBt4ZxCEZgvWxcCfiSMQCunWvLv
DjMz827OIjBfFNfJAEhgi2qbpVW6KqUjw9v70l52tHnCxLil6TrpuBXjg3ZaW93oqyMTJG/hZd8F
6SA+IKQOlSF85EHeOYz32pna0gko0ABoQ0K+bbfK2sYOZHkLARNHX04qFUmL48LlEdAT6xGchccu
VmJm+mmqMrmcGuxvocl2IqdNEGWkijChuN7MJUnGEa22jeUEwDuxZomvExSsFdoZvz9UCDJIapjl
eaa4jWe28eigdSAVFoGOsB4lXzYa0yI1AGKyicGg3Zpaj0tu4vtBoiGHDMI02rY2Xb/n1K/jUNZ+
QhrOsnsEvcvO3xmylCmggM36sax+9vfyyuCBal/3avVP/1FrPHGRSsQmkRk/7W/YY3dX2O4NguaO
dpR0aJe+JGZBdhXQH0K/yriHP7FTgK5cjtqnXlwTrp0xjl2R4/WoktWqqd55VycrO412e0CkHHlN
UINIhBRB90taKRlvt6Zzw6Q+uH8Y3Xw0XHLhFc9dhYJjUPlgQki/ZQWMp8x0E8zxWKVNkB9XxEbE
VSAQvVdrSl63ARE/Gh+xDtXvIJ4OJUgZo2+dB+ijxNVRIcY5TSgIaspYREU4iwmuUWixK8hteihq
zKKkWWxero6BfOXWTlTaGXDet0wPwyyP+gFoe+ivZHn36WSjg2Tm3JIFj92Al+Q00st4DMuOV8y1
1tPLMImfV1kszDgEnXJ+y/H6kEJV2oFnH3XZRD+bonAtPkpDwQ7q5XOhpIJQhfQwaN1W8SC+eQqK
0UdAq43mKpYfD25BlDMgGlkE1TA/tcwxf/4pAqyJP5VP1/rs33Whe8hsqmgWh3eQE9w8ph0bSSZw
+Qlbfa7Zj4kV6XYeV9kpG7xtY8VxviWWbePHI2Njemd9EZJIxddEdiLS1KgfjC9HtZ/hJSHK8iO0
FboeG2nPsNdTvhJ8DfwY3ttpYfk4FNlhA0D1ybbzPZQayTH7w+5WncYeHSzx5GOX5fdvEa1nF+aZ
n+SVNkajnTu7HMj/3ubNl1iS5nukCkPR3gquDdlPqxZy6I6Fkvv+gX87AL1RzLXuwU88Ap1ZcCIm
tKHngnf4ds/Zj3XfRY45L7QTy4/tJrW0Mr+TFg9LgummW/YPFT6cl/SkuxpFOzhgonRxzs7G3P8J
dNWqna9ntKNBTGi+cnGOsAbgCreAR2B8XiTY/zwqIdsjkJjoGWcz212Ysv0GPboYpDbSCAkcqNdi
EtIAnmuor45ynUbe8BOcBDHgxAZ/rONOZAR47YcdO+4i6MPwk/SmBOr9LX6shyPM7EEHwtzmAd92
Y4s+z5wEgCNYtTY4J6y00661ye+sgzrwe0oA0QeXpzC56Ftks9dSkMj84+9wMuEpJMDSH7KT5bjl
ZI5dun8NJ9fgpSzPaCrPNXCDyixrcYiINJykRpuL2djtGQ0NTRGSpTSoNIDGr/K6Tojc9aIfyoWD
Wdted9otUxl1Zt3Mi+2GsAE5rLIbCnm2+OKROdr82jW3sPsM6oyNM1x12vxf9AVP62oK5PwHSdOG
JlOQ4kZV6nIOzL2sOv+tMpUWOlzVbD6IBmfQfvrDnfa475jx4qkzBx9H7GKn6wLWsj63kzrUsU7Z
Lr6yOEZmwoBp2+1BRDX/bSUeWGj1E0Z0MPuZKVzHqtRAGyyAXXY9TYEocWd2W1uJqKei454ZX2GY
D4IUEylRdqBfiAJCTztvBD2DR9oA66cnvjMD2wocyGgW5hGgzl/yJcai5E72rxY1tJdnml12dEtA
lWbBNS7P5qpJqjDOjr32D9tCcUAfq70ltOtyt1OSdXizCEtVcbxOO8j8+Je0QqfiU+sGNaPb31ix
8ovXWZdcdt4xt5QPIlATemooHW1t1M1TqF4QxG4xUowhxFaZJgiAmkKT7snXYROGmRJrmgngwGTQ
SWztU2YcoacH6W3FmayDi0AsDxBVBcqJ3K/hJNLXu36cAR6CrIl4RK00t3yui5sSFnl6VvvZl4lI
saphQa486rTjSEndevK6aL73ZFJm/nGo5VeF2J/CXZFyFH/jORpN1R6i3ifGOwIkXFB16+OYmIE+
KDT0LF/7XQ/m0eboRDT71pU/NuvMumRp+iZdlkkZ52mzW5OQlc7YMUDOYrPUThZcPf7JSzJKFQsI
40C/yo8XWFXUTdXvjL7W0twrINFazWGaOuyvM6IeyjLBqP7eDSeYKUKWkfFt/9CqcIUVNyKqpMq5
nlRAaEPXnyAEzKRHDasfr5TmThQWEGC0sLp65vgEn0zlNkwnZKh/cTqFA3AupzJIaQJWZ0PeqKNk
O0HYLFOrueaDu0cEzEZZkQEOZJrSVevjAX77PmK2PKkyszS3JvvbUA+I3ikZjDSTTmaGOCxmue3X
zZlONh8J05e5pq9PrsiwCV4HNN2KOTEUqaQsgXuEbFJSBgstFuD04V++JWXcPvW6r7Z4750aEpYA
KXhMY4+l1fzEwXz43ucUBSYbWQ6OoCad3vbVscOaDwsYCnWccA5fRXYMWV2RwpqFlDiMSihZ4C2s
HBO14UUJNtTokDjEqGi3vO45Ead5VoNfsEL+5kOvIcVzcvcSXWolmjS3lqNGAVvtToWLQZ/1eMPg
3ME2K1ocswvnZtUSMUfn6gcdnb4Z6EMVu5M3eoQ+UzeSiafX5ivwhFElsxJWbLKEr1+nvk62jiOE
ufeGqCLQRf5cUfOwyeh696pNMQ/BVFberjJ/fRh1jil/9k5XYXaV8cWrWplD6oZ7CaWs+ifR6dHo
m0nRvQM1k8MekJdp5k9VaKdArPMskozFTToLTCPWp5linUeNlSFLttp2viW/kkN8NrYe5W7nF9ti
5y/yvK73LTjjmEauBuowrRR7ccBNziCqSfe+Ek6RX/51J23VAtKMFziJAr+Hp5NL8Ut6aISJnEKX
WJNfhr78wjdO15/SdCoFOFyXVp+OGQvnMFL709cIb+NeyCBWB+Ya1E4ryiwv9rvSgmgBadtAmO5e
GsO06JeowYo15wf+uV8J69VERwbA2/L8riHp68563PkjXFjxHHNsb63ZZt5WRDbnGXfQzyPfrcDy
Uly+IEpfjLUDHBBR2+b1h2WNA6u3H9EbXF8+6N5qQunTAnTfYUJaT6D+I6rfkRgVgq9AHkR0kV1t
GoFSbBIuq/K4WgS6lht1N3FsmHp1HHTs9NkYZoYXEDsbbjpm5RGA+nLWxbvAl0u1XYKcyaPju6FW
Fc086I63IJ9HPyMfRp5HBmvpgHhVlyiS2834wGxI+bUiksGPgFcAkLVuluSg+Pvy2/5c27Ewvwx5
lEA2Q/NcbzrVQf73Fg6IkLwBCxjIAv1cWovEOz76GPLmUZvSinYmfJ7CBGyPen9wnZkfORYeo7Ga
gVD+kdYh3p5u+oYiooZOwEEPfq7lv1JI3yVG57NE+lRCxDdC2UdwC00otNhuFclomh8bdeTBVrp8
EXk+A4LHE7TyIG9J3TB4L/QbN+IOLGJubbGVxV30xbMKdJvfadFATRsSeYmJr2NI9I/TcWTUZaa7
JRde5FxLTA5PzbIS8bto5gxLUGrkHF8s9uN9qfkbWcqiJteLkei1NBesO0yOV3k/pKxxRtXCK2nW
bWfpgvWGTVF/ypP8LLhpuZnapDN0M7Aa76/dyoaBJJbnbkVCFxxdDt0BF/IUHqXrRfTLLHKgBGJe
NavCa4w9DbAJHDSwPQlEi6v4cMHBSJoJ+46GFlaGoWoOadqmAcqdwKpocTIQ64QDOuWBRvBdWB8g
TN/63AaaJGbp7Pkho/LwYjS+sPOXucBtlaSPN0T02/5YQXYOW2hz0wH5wnRlG7YWlZI0NO5Vr4Gk
41QnFZtppmEz155dWzhNNN2YxNrKrmpoxEvcCc1K3f/wP6wlTYUFM12rT5HWwFQ48sqBA17/d8y0
B7Lf1n61n1MXuNJrDv+fVo/KUKyXNVYyVTKDHtXFIGZtYhEIpeW5CxWOXG3hUlBqNg+G1QIhkah5
Bbr378N/7K7BUpKM2n+mRdYh6d2tKqmoenRgRBFGKF/l/6ZGsfWLeXEWWteHxsEHiPVKus6RwEzv
zeSkseelxjeDTHYmQ2hAaq9kH8yLKkcKpeHUe2Hm4idqOdlRNaMJ57NDINT5O2phtnPswy3kIDb0
GUqPTOsraDWnro1qUL3pfubtJnCw1xb1SzEnrETPRcOyvBiW42SPydLJbEAw+UvoiebWG3yTRsz7
EMugq8d/NTJZaLwA796c5ucaqYhjeyBhksC9sYDubeSwo/HQyZwb7yWGlerae5VpBcpIc8yEfNLC
WpvmYJms5t1UtSU5bRh1fDzVk7ghxEVQur9o2pfYNI05zB4cKGdDUgxZvtEJI7OQtQnYAsziaggG
+DMJIM6e4irw1M1QONxhgbrgKMsHZ8O7+an9R6rmEOgV51NBYw+QyzL69m50cPSRaP/1fL1Tkgrc
1F5mLfxUNQbeoXPJHEQLoamckFTC9+JoXzBEUTjAJXgROegfVW2SuZx+wI26kQJisbt0G/3Hw1Ei
+Y6PfVs+iU7B5Q/WysNpMtftpIrHR+ezRxtrJUYQU2aGmw7ETdT7DoHhXSpQ6oRpVS4C+z5TEYma
A0F7OzRQb85TPjFIiNBBjTjeU3xrtdG007N74FnVQk98B9a5fCVUB8PTlO6yZckKiC+QGXZJld99
OfNnXvkd2WxIv6EhW+C00QPXLMcEQnDTCb6cnZed1L4QV1v81jTBAP2cppOi4E8AExH/rjvckqq6
j74VCrX9MxmQUL+vOqoT+H1d2UNuiLS3ZfSSWiZO/Y0h8Os23ONxj4S86qUOQPS2W1mhVefzfskR
V2EdiXHFyEOmccU09Jn216cJNuWrbdYgtlyzetIAmHwNUOzpNuvtO4WA8uAY1itFDKcv7V2IqYb4
nttJg3oi/h+3CWR6GMQqoowG9eBIiA+NNP4K3WtXVlUF5HTQG4drxgJ3zWAM+lofd007LKOEuQKC
WufzaVIEo0eb2l+dYyz6iW5msfiwTq4QkEBemmPDOmveGxcYHxPLVkPx4X5AZ3eh12dmUMDmX3n8
YW7R2o0jISmTTECLovZQxjKXVVwS3jiAopcPgLDgAoNutiM6IKxjkz5FcT23cRplmYxaEw01J4do
Lq8ANLGPUyH39paUagew5hY+oekPirnxxugxDs0HGwFcuCKChUPo8gUrAXcyY39ZK3NEXDqM0IFj
i1H8OZIcnixXe0PiIZV+YWtg2PHNo9nOUrOrsm1u8jsdL3hPPoKcv1lE1PO+nU0p2OVDp4j5o14t
HodHJynoqg5lC0iz3DOw3QfAyjVghr6GuDAoWrCH/FbpmPSxi0PIVTaCQ6pNO4Fuir+kYwDzYcYY
GFCZieszbsbGYtAM9NL3Wf7xCgJ1aF2qmT1PyuDYgLU6m+HCCC0lF//iItUJwpTiraN8kvq1aAkq
qZPRfkEoUgrkI3SBAtrInWS6NTD8MhQcb8ZYY1osSUOrddKSNXA0uTvYCeu4RlVtJa8Xu2cq53un
CVUv+bCi4FA0VBpROSbaR5HAosePIBydx0BEngjQ/uw7wjksM6WSOW7v1PkgW3jJ2Xwc2ItdLffU
V+m8/06uBzLchmgI2nH0E/hmTIuJd4JMnyBktL2+ZQwFRtQrSULN4g/9Jqg0QywHWxTfd+g6Y7b1
/K2feDRTFl4OVMdNYEYfHU5AHW9MaO7sdqjxyuipxsk7Bkm+zwlZMy4Z/dy8FBqclRgCmL4lePu7
NAGcQxgfZtXqwD9BAWdspRK4xVC45UjU3tnhiX0noMmF+Cr4rplMhe+/7P7oEBUa/BPkMG4S4XH1
0S34RItmdSl1OlIOQmkGi1EY17dgPQbkN5NEAZM4l1ds4CzKXUC3UYP7VELL2sl7cneztlE/Qjcv
5HHj4V/JDHKYuMWuG5Xgg7/VOZ/20P+JlYVjfIbSay/3z1b607yl0psqooJhLwoykZKzF0n/A9iS
SS0U50lhhS4rHd0bqWOLXd7uUjyb388Mg+1ygE4K4Ps0dCIUFaAoEQcVTZ0pBjh0M/p9yzmsemPW
Oym0VzGfY/5h6GbQje/lVgNWewG+mZX/OAOTg+RplXJHpsxCmteTXmekfl+iIzB+7in7PVQ1WvpH
j6IoTBem7Rg16VJ2mDUHlYCSE/4IX+Z1mZOLP+XIMMvXswPt3yJMYmGMkaghmL1bfJjgR8eIOZ+z
IMkpBwwsjx7rMz0PTVAnSVPItMKEsAXwbMOTr8BV7UdvHo4nDBYSRhCLHpzY4lw4lUvGnhKRtzoB
09/SlyEOoVlyKMP5HHq40cLgbPck3JU10nho2IIP08gx6EZfDCeC2riA8fCTJ676jQfuscjam5ei
zEfT6Li8TMtz9oQ4WUy5EuZKxXAE1CYLWY47JfUxw9AdDO6bo9Y5BJdOCchWqDkB7DkfCd6BsTre
b7RUkRHLpwC0PcoNDAKKaU1/hCtIPaiuvcn2TcyZQhlUe5WEzbUfedfkyGZEzeMfu+qsVgnF7eRu
1ZsdigmbE13ljTh0XL3iAG7shD6eYz2CfsW6Gr8du+8oWUPzbLtNokhYmOUbzNhZJDKTMwFc4ns4
QIFJJLg5R429Ugkd2mxu02imfijoEW2eOVmDxgd2CXGU8nqKGCbs5/VsKUqgMB9ZY4kWGx2Bptqf
KXYghmyHCgTclPRpfEcUxYtCqkncXk0Mw1VH54siPgmfFHX4bOrn/UJxJ+9LrbZdb3Pbf8wagkBa
Mm8o8JFtg44q7XquSsq5pVtto+kE1ocBwnDH7ae1egqPhdLRqtMI+m9KJoEBgXLWd4GIbzRdM+f/
CBFcAxDBvPD8MYo32ODVgpnmKRrgYfPqE69jtmIMUn3XEHo7CX3e5JZEjDn7nvWAzClJw7Kv1mUy
IqaX7qRHjh3cu4FsyWT9DB+v0jyr5EzpKGItrkj1veUCSCfqH6bE/k+NpJ2ljsZ0ylfy8u7GSmuG
d4kJ9C0NS/a3n5nbZAP2yQfUMc1aRDiQVD9KHEp2oWrjW+N4QvTgl0s0jzBH814+9essn7khQV8F
YUbtJEckObiXVaDsrrux7VwBCqwp2PosMsCQLYBNXEsJhwayD4jcS3126CwOQQQ8PxSvhpuDf71H
lDsaigsjziw6/GQOcVp2nBQ59/TJG72/Hrf6BKzeoHYcC183OiRmzDsIYsirpCMX1W2Qg7G1XPi2
kCVRUGonowytc57psNzClTzBQ1P3/zwzKRBqYtYTJ6dtKGOyKxVQZPGWRlPJQLU2tqaAqj/mYMMX
DGtGxAn4F0G/5rDoHdJJ/jCLUps7IluhZpiFgDPs54bjQ+ejucBmyHMGQ8NMKXu4SjXO7fbiq3Ml
5vN0eWOEOmBUNRsRij1SypIqnudk6UEOAC5Jd8RLFHuPb2gTUhKQG198vp9clbnliaa8CEn1TtCK
fkyVE02o4SrKfKra1dBl/YDchglSR4BeRiNEwUv1V6MtFywPsvY7fgm5yXwgUuo1nmi9fqIErtRX
PKmEknpG96DS7Yq3c2eaGV0adHzgRo/hgWxsUTNWn6bbjyo/FKt69Mo9AHLe+UB8QT2FL2qHTntD
JUX5ntpLr2Es2RERRDrvkmad4+ulop098SQQrEgQH4WNiBOsgTYkMZEXB8j6RSNiginDgCrCry9b
KwbgSc2TL98UaDyXju5ksNwYs37bSCoUcuSwgRWlEYyGyOKP+HQxx5r9AnNQg9b87FznWvTJHqlP
NuVzP0m1+zWDH+0uqsD/JDIav/066JxIcZbMkzvgwbhNSBdqprMtEs6cLom96SIwJmwUbHd80uGp
Jr2HAJOheBkIdlP1qcI77ov28mbVkIwWdpk7TICaPEjWPFyFKbIsN9DjLjUdwksPkcqoxMIUEbuy
jJW0SeCQo0caJPQ7xZC3uTnlTbfEuJgDGfgjiFY0f+BDpMFap5JRqeQE8l7Tt4RoHbtEHWw8ZQvh
dYNhtak9TXo4YmNGjlvvcv39MHw42z7qgC8QoGIi9DfGy5Nh52u+OiLRMHBpKyUZdQuJKUkJD3nr
D57a9eSkyCRrS1zP5QcjQ5Zj8E4Jrkxj02pv/3jzFeKbuYhlij1zQ1Bu5qly6M6ApQqSDdqXFjQb
TKSnA2ciIZa6gf0JUm5sSP8WAYg32mm8jWiBWhh7lhpOppd3sYYY4lUcVb2jP3cUY5UuXMzHkups
zIx/gnDo1sdf1e7vNGQR7MaDzOBGBduBP14IG5fcinpwnsvmZA8BXQExv7Dd8VhguLeRgerAXxtf
7kAe6od9jnIdwaeM7RwvR+aSaiWXk89Nlz50OElc6vqhS4FdrBfVCyNiSd4I8e6xdU2rmaKOgj0A
JE82AWbeKw2drqjFC6TGCXJr/LOrnpxgPSQLKE44iHbfTZVdEB2SzTl1Xc1j3RaXtwbNFN/T60Nq
7G/poVUX4MiugJ7DU01ttNL7rdvLidghn7MmAUKWf3VpUeswXC9BV8C/p9+ne1lAbCGqWL00HfIs
er0qn6sio7WKhB88a65pZ1et2r70+ZmV2vKjvBxsiRnxL/2rXvU3KeDRGRhkQyKyRTbfa7W8Ub3f
oFNqlm04OrFDhN64oevuwz/wc/rFm3sAgFFREVwLGF4d/XhKiuHsuCHr7Q+YtVAzTxE0v74Og9x1
5j5zVClt+QOCr4bXEMKlzDqjl9veqs+UhNK/Vzyl/17/hwPM8PAmsgO5OSUWG+eud6LdCmFFteXr
1BfuuXW5yB6mO8gSw9o0XqsPOUdqvDKGirhapAfBC7WZreQZiMjPZeM89nkri+rUulBmk7o1/1KQ
d2OuUmrNWiCgkrGldhkPWsOeDn9v9ru3tdxbxOmITskb5kzOi47Jpk61tKhMPoj5dWJT3f+8tnqT
zMWul1GkLnurWiMJZ7Ussch6+F05gta+06oCPsqvPq0SpSqJ2L+VlS0MMjvFEFZKX8Ce/1+q3X2k
K5Xs8Jotf9vJuSxrIrhvlHVk8plh32wyBhvcWQNa+ujK7zpD2+HBge1TUqZwmSs5eSPy7WUSQ1n8
r2t3rFTGfMFfv4nsZ/jHsXL01ykXobtsp+TMp2MSv+rbYqbZsPRFPc+vAhGHL6eQgIuOW1MwdZ/5
8pkc4sVUPVbSiGyGpia2+quiEypPX0nn3YA6AubZERQH7wB573oF1SWD745mlUEcTBxvCNbPuW75
D1QrNmlPIVLvgsJYGAMA45+IaWSXtwrVN4+v9jxqqwCC5nNXPprujtTKm6NP9s+KJM2iNA5qT1ZU
ztOfyG/TdZ4SxJJY5dlCnbJZLQSbTnZlvdf9zGl/hW3EqBHlhOtIv6RGWyRsmdWYifgZ3UGz5GQm
jtgHrphvfAmTDTIj7A+ks6em3KywL2697gmGUrQN8X/HdCVJxVHspXJ2wAIEBewSUUUF5Wiq6bqy
15EQ+1W4nKHh3dE+FR5YTbdKaUvDOkG9vm+5ugRZwmnAWcoDNX9OTbvfWaNZLqF8GtysArfjQ9R8
ohYmi20+VP0kVZM/2zMZif2OdC/Fbwn2no3qEjtONZmMSNq9loyf+TCdT8EP41htGEopR9dX/ADI
fmh9vgKe5CZgpg1zJ9WThi/xfFQyVXs2JVw2uvOopfNwuOZKgebTQ1QLzXmTMCZWMmW5u1qSZrdl
Wp+ubKk13Vf/m3pqp3jd5qMWqe0W+OFNcJxp6InH9ZmlpqVmZsz0Rgxb9nBoxxaEZRPRXPBmTUnk
Lw9m+waaYegqSbAvlLp9H2NAZOu3ObHSQYmVdbWS/Ka1HUX8b4O4cgfEwa77usnprPJz78WaIAzS
8Jn5eVNY6S/jyewfZ6QQmAiXykNrbM44xqQ0e+DuoRHeT5RVQ4jqDvy6XLqVcGp8Ta3tj0irw1kd
enSdFDOdlovUJdeAwO+eyYYUu9j+Cb3LbBXl8O0dZrdlj30FiaqrKMt90AK8E06M7dyw61BKUWlp
YMKUBFUdkcjG3MXoAsdktmkNsohoEIXCgIferB/AmHAqN0oafkqrPNVBuw2tTTf/mUpQw3VQ7UbO
QvcYZDKUp5oKMgjLVNTS4cfjURnBIwiwfJf6FkRfp5rU1B3Pu2wZ0E9NepkqqRW5N+8tJmyvP9mz
rkeImnqzFfHXvbMeETtR6p/PImJGJiuSPmTOkCUDdQG/99OR+GJ0p0x73eVdts3Dk1qiW4e4nP4t
tng0l7WICvxlcrSzAmUlWln+TikV1DM8Y6UjSnKhyLgw5aHDajL+r6HU5Aw8I6/TZryIXsyn1/LI
7lzj239sZQOyilWeqE7o0k0IjWXUa7P9EsOJXjylXuu01KZGg360Q3P7Grl2VP15dQC6OJIZ+5fE
lAJkaB0610iXCuWXl2+5T58J4kvXORACvzB7LkrKrWuyLEdtlItUqqqPPCyJoJT7ERX8gxIwCNuG
iLWCx+hAwAb+iY4YmVXgMXraLtKgDvibbSv5emYb4taym2WpYCJl2jhZCNqvw4S3iTTLoEwl2R1j
uC3Va2vWIN+bTg3sx/wdMU/cUFQyndoz0TszCc0hfkBkEniqDxL9xZBWhp4tvPy+siirpIg2wY46
y6iHlIv6BNDdgjXT1G47qvRxGpdVcbGXhOPqs3succYf/xTOdBwoe4TEfldrQ/FqzSYA7a89E5Jt
6ilrgEZv7pVGA85EQChGuniY2aENyNj/zklu4a3Wh15ED1OnQ7eKClRfO02iwgHYUj1SNd8tsxx5
4zeAoooDdNi89tqjqCQ4qyrk/Kn00B446zGex0qio8li81AZJG/oaicbz+7kcR0xe0DT3tUkODp8
wRs443Hy11c1yegtjQzWV3f7Yysw2K6/kDaxa9NzPr0XAwlh6RbsZuVCTxM/SqF8VehL8I0tQFO8
4HdQVRAxnFb5DtJZZMe8Io7cegNbxPwkzF7HnAX1Rwo178tGJ+fplYy4ALOpCrIr87GZnsgkTcqm
sWhh5j7KmUR4K/nrQQB23SVn9Kt6GRXZDveIQPxeRfSl/RgulNlF1yKyf7UzWcmsNZpojMfBoa+1
yXORzZp5ZOMRoU03WrkBYbNvezB9CZPem31DmKFsGFBejR7SoCzBc3BlSJ9SDiqVXNy0HxWM6Ly/
e0XKwsChc1kjEQ0+fD7TsXRUPQRb/yKJPY68dPp+sLcb1mDl6jMts8fsIoC7kneFrXmbRAaaB8S5
a5Nj/LYYPqBDk8/b5DXMDKtB9r0QICRwTmgTas0hIhnucCoHPfLz1LICt6Sg+YoxvSGu96XswcK6
lctUeUSAYFdpffNKM4rqd3TcKio9lXGjWtjX2D4NYcT95QnzHt95ukP2b9oA4FBJntKP6OOeRRkJ
3ynilFSSZ4zOhHBjqTV/OXGx7sS8s5yJUZFDp3RrQFoEE1pWYKHeqmktZA4uPdpwmcsn7Txdv8e3
KXzI5No1T0Xx9ZZK1J+Ik1wLHM64NOkVNZdPEKIEvCDwObL9HxTUr4AXQf6Zlod0e8HvpWvxk8KP
sMkco4VjHyVRzsPHlP2mJ1WenM/KzeyTRTNPrAsZQwNkEzXAOZQuZ62sw4vJUSSd/p4hWvVE09VD
K7qPMIN4k+wKDES2p7Fxh23Nlq+7daG0yeW3iLLzORpwMU0riZRxANy0NBzdEtgBRNvscOBKYVpf
o8TFWklnBJjJKdFVq1dWygdVViLZ4ZEFHL97PTT9hQCuTzkx3i3jNrFEPEzdrZRfbAHIoADgFOpw
1v3b4bHn23gbGSbqDJVDnd6IPPcl1IvdWOpCHOTH7qlaCmNI8+l4xdJRXLoUQbVvcnbgssawc2ZO
3CP5T0B30xXzrs3HClTKXfKaRyyHkh/nLmncaPIfoQ1+jK19a2TQCOBvonHNR0HIAZYZsblt4IjN
fmMTmREf8bU64yPqqxPekpgGMtUIPE0tnovbeZfL972HIuuVfqlD+xPQaGxIVr0KaTYhmA/Sx6dA
R+qZb5hPlGZ/IDV5wEnzAXNUhuFI+3ymlMI5sDz7hM3xSgAlgwGkxyoi5H5QP6hrjToiGoKgvxpr
7WuRRS3dmguHvxpqkZ/SJpY07WjljvUz8vTxrS7l1zb+feqJcXy8wqNHoF4qXojy0sCPC9fhcWrb
qzkgTbjsgunKSB601d/V/JWwxNX8GCTaa4/BZDo2JLQmDgBb/Xpi0lekTbJseUxB3/Y+ty83mYjh
rptjcW40Fykz1KOfJguiWJr0qtEMWK7qSB0A0fRXBDwAG/4ogJFFAo76nuGtcsuPxN8CMoOKjXeg
KOCdj0O2XJuHsQzm74oWW9bde+5rvCQ9rT4Sqs+/knmLZk60W4se/mS1UKDPYw2KD9+LrCgRjv8K
ErckjzV/NJo3z8sVrJGT2/1Lx21Uh38kZyKXmF2vbIhm6O1kTQ0VYGDvDoxgE7OIsgSJ806Z+mUj
TB25tXJegSU4LDwUYl0vdx+v0ZhvRyEKY5CFUv12D3ddZb/qpgyr0NGHQNvnJBWTUbIBu/ETpZoc
ZXfm8DH9jy3BfQ2k3c9F7QrvbX6NH29bmuSprs0AbwJM9Iouzqcx0ls8TLY+5zkp+90M0MMoE9SW
3vXeLdZPfd0tGq7GC7O2zOogkiOQEWwoPM6mapCET+1Lghws7nCGzde/38x+b+afNPaDHNeozawS
BpJdLR+qVky1nfPkPT4RosPjBaOEV9jshz7tPWXPU84pksIpOGkseC3EtiPk+7R6CMCQRZBxFsd/
VTg2q1fZL+Nnnp33FVRozl8pjLn1m5Z9xNaWJesJ34CIxzkssCRg0ir96e7OIzJNsvVnpdD051s2
JeT8oYephT6u3WBEuysHXcx4M0vE8jZcYobvsmGGQjsyttXrwuWU7IRw6rOjcTqRCl8XRD8UsRN6
t+QdBG7k209/3g82MjdEbwyd2yiy3JqPK2YURZvOiDcvrJvFyRIsDB1daqshnULev96XzMEBWu3z
Nq4dquq4cCnvZzwnFlcZqfkmjpOJUnDcQw2gcITtjCDeTrNYnaJlT4QV5T+/rnyECVKr2pAYqlMn
v32pLQIoTMAnznJPwjPArEOM34LTX7dE3GwQBVKG1qELu2uw6MtUN8WIVUN0j2vGV6w6iLY5O9DX
FOXVs6Rv4U7xyYCjRW07zABsuuA2a9kJosjVsE+9aMhM/4Xu3iCav2Kd15Aa288RcUevDvolt773
P0irkd+wUzGjasbXeSlKwJGcEu2cWn+G0RON9K+zpFXkXE9KVxwlQXn+bOwRHIhLGgrufH8/VAzr
ZSaz8mpU+iWRrTcXe8hREwVV7b2TWV4Zjk3kkb61mWZnzVXgzxNM+u1aGxabvRxmeTtyOU3TMZKK
GKJPCzUiYbvUTS2pjlgiZU79B0v8KYjds3Gt0f5IQmuTxaQfDN0IyfB+7V3gIGXmbQ94Xf+zd5Hu
D7OJSwQ5KQUoASJa4aX7ZMBWZvEZ7iEcAaTCXq5foO4u3bgfM1frwstU69xAueajJieRCIniUeLG
d81O/kbUoL8MMRn1Cich65frvljqzuTd7yXcUlcepYS0W8+y5h2+otVsy54QUkxmVrmxrnspsirb
M8eoBVH4m7AeMRpMindHiLM1L49GPEk5kOS4++y2cOvI6IB4ljrsbSyP8iPlaFu+kN+kEsPlOH57
zm8sV7C3PVVki4kGk880srKpS8rM2Kw9oaaDS3mIlxnDCr9EzD9WYO08R13buWkI5RygYWwsFrIa
NFtWG2+ThwOPTzxJxDFQHstt26zd773ew1nic594UwzS35AXIKjItdUdF26Sh6YMxmImws+1nUm+
Z6HVJn04b0gFckJ3hhieh5Ki6LemKOTqQ/Bpik8OsYxADE6PX5H32lV5zDoleyetKm3XXySkj5CE
MlnVODbMy8UZsJzCJJEYdVt5XBm+mWiR3w8h+QM7pSKNEOUV2PDWkGcy3UPOa38GnduXYIZSn/Kv
thersVxgPVWiTekc0jR9+WiGYZUlyDHqj+FwvO40ZpgK1WppULqnbwOjMzBagNYsp6JVArA0EuRP
qbH6J0KU3zKCvacyMREBfa7p+4GZafji7nEBDszczm16kTCGXHetCitwe0dylZUZFTy3K7K0CNlu
eOywTD1hDC07xFmppO6kaH+HEa2RwkchVGonsWhLxoRXJvZDXuZkiUhNvabrIp+ZVAQuflp52foS
md1lpvPXxlIptLUKtEnUFUDyq7KwXRTGXZxVUq5fm/V85VyuSw3BqEUUr4UNZhTbJLkWHd3eou7z
jmWZ49TvupgWthGj3U/frYj9QM2ZeJC5cvSzqQ3AE66A2Qvho6TtJp+6YfvCMFk+Tu2Vgirh3KyH
DCqwWtpggzSQoHaxDYxgKghA0jSIX3PYrZJwbO6auOPzBGie8ZetLbTU9p07L54x1kjD6B9IcZLz
CriruaPyiTPWntThzKDo+9zcWkcZTx3D0xLnmplt1j2FpA7jFcvUrV4RxuYyDRSC17yKdubvNG96
FJOejbEXSnAToIxAjUtEpTIRGTJDyAfEYgY3yGxPdKo5gBJQLUtvr7KljCIkBspgp28GeE5rxJKo
73oC3W0AEvv4TSsVQZBXI634GGuuoBM8x4ad6Vi4ek34HbE/jmv939tHMLFjknjNKcJpO7649d/T
tNCFtpiIp1EWI6xmPU5xWQmrmPYUtNAfX5XLXQq8heQd5qUCfvgVr+eneCO1LGEuCFgpOROqduI2
5LVsMSd9XzYBzyOz3rWhkyiswwNiGDv9ao+4Pgt+B6XG27HHhQv5jlDZB71f5uTDKRt4D2cJOYrp
WTnOp1uca+Mc/Y//REMWSzV5ttaTZemKqp1NtrKhZ6gilgK1/d36eD7c0zSCGuAaYg/NawPItnv2
llMgemWHf6yafNwFlMQmvT6uV7Kfbn7qcUBoCYu43cAvv6VbhsH7YfKiaX8fJ1jJUZT+wQJsX363
/x1JnS4tX6e5ignj1Sg0edIOmk4N4vwhihKh52nP7aMtfvSUpoz0KJQ6G0YPmA8G+nH6iCAshBJP
aZNxKxUSy5zGuPoQ/IobFwbx2OyvhO9Z8meYApQwgjMUGJIgGZTtO9p89l5oS2FLvKTZRMCPRroB
G03aB8t933dUhoYmSNfBsHn4Pw/2T9u5vbTu5+XdwHKmVJ2RcXDKd1GkLmO/VkhnSHlpsk8diCoY
JBQuuWMHtBFg6vUFD7x8Nv7eUGlpYxhc5Uhb3J2eoCPk2lgtohYDvNqqs/WZYJ/IAgaTy8Y60Y+d
D0K/He9u/eXrTnYa6DO5wgHvscPBpcymZ2VIh57MlythosblDnIdeR7ztxIYHqKw5qMxK4NzH4+L
nxqGk6J/PlXp8gWyAitwraY0kWNiFREsWr5DiyTHgRljDOtx2y3P8bGh5Su9vfdnrUVPJy4Px6qy
+BU7wNAibDqdDWk3OPd4wyOmGmJ4pW5CcLCNqM7B3pe9Da/GVq3QSZIZjwiwsU7CjB88EE4aSjUf
FzVWn3W3BcY9PntmNjcXr3VuKYCoTyTDPPCObsgqpXejnDCL+k2qpG+3Jh0SPHFzHioQFTUtSrVo
yGYeQ5xk3WpK5+QX56Cu3x457D42CqGwsmuCDlvLkAt3fpZyVokIkapKd1xOyP+uG3BUh3vmboKm
rFfwe7quBCbL4j/cMq7aiWfA8yI+RMtft2ZGJLUDiBYK9GdUxE074xlhr3i9wy+PBcsx2qpgoTg8
vqZ3ApayTuseoxPgD538HJAdu7+sKrX9MVQ6fL9S0vKYYyd9Ki7TyjkDRHFj3s3gm4o16JMYWimD
vddKQPqtMqW4aXRBRpKIEtvWawWVoD0HiLVdYUwW2KyKf/WpEne9WmuRMKYmJRNFJfYn9FIHojJN
Lp71r5FMUB1+rto+sYEDiUD/8AiICsJZn8FtLLL39LVm2Fx+t9ZnqapS74da0gc8aYc7iCesabgO
QNKgLwI4Zn5cOdF+cn9z5iTVQ+hBq8pUB6P2TXNHbUW/6XCUbJBE7vcwb8SURrO5D1Ks7SaKPGVG
o+0+XwaPOYJIY8wfqV2MgFjBI29BoVRjD6/hQipgWWFbpJmFEK0YSgyWbbUaYBjdzZrhKaeJbKmy
4SIbtGRPFSRWNtUqr5scMTVFiSFdg5WDFIWEZ7v2PFHu8NIn7le41fGA/4kHKRSWs/BMHo6FXq8T
FqKZGELW9TpZhgsyBUDZWE0Zin9lKgWMF7d/UVYV7/oc9fa4Un0fJHN86UAaH6Z8hLzgDkxyYsAU
qpFrz4RyWYi4nw4GWZJnoGLutpCdNV3KD8pGReSZaCuUeKwrzNfS4LIjuM1gqR7P6GzDn+5TY/BW
CPOfRq+QlHPFzuRueFSXLT3aE+sNQ1JQ/5PEc3g9ztxBy/Pe+acThqfsZOHKjeKsFHQtDsG/dVTl
vGjHDg/XUzLoE6qJ4EPcuPIVq6dxaY4+d7ogDgabkTLn74ZSWas/gW7uSr0NHivQkHCG+hUnGlsF
R7vPsiK5B1SH3QcCwHOxsLyOYdqMAF4WXTQbsJarihlW/VE+6Lr6e5al62dl/Fwnx7PH0+IEBZL/
9nVwv7vfjSxdUrGEFIB2y2UkwKZ5nBRDtV8GFO4voFH7Mexcl7dv5maq/IBBYotPqer/y3GyueiS
C2OaQrfCOxxIcEsJuzoGxjPaFcV8/+AEnOXlrOSNShVHzN2Mv2j3Q4KnZATLkjEFJ4zJVSwuXWgR
WxwM1rZQCw6luFuXvlDQKVWh48IRD9CTtnJPIpEuccR7PW/N3JLDqiaowt2Bp02OPG+HtDIFe9oi
DQi+cMDMZQ2ciA6s7o4GhFLaRxi5ZQbrrm47PLjtHHNSVWbnsrQYITvcBQnqV59D9dLetDBEGPIv
khmtiVMKIcVGVVpyX8DxMISFCHOnzUmije7azS96agsMx9QmCwU4ZtDfRUllFyPbSuJci8E47O9X
dhkUN2AqghS8Oy1M/+r03DDAMhBEHq+fIvDF4PXsanA37sYf8Tq0cUxhSp/Sz+bux2h4bnnMc0Pp
jxprpLJZUI4LDB5O6am7+GfgJYMuBc2LXpsvCj5arJEJJHb+69Y8TQbNIJdoV0zTr3X/KS4kaRXF
b7PP5MCvmvTptVANaDhMk9dZ/Y9HoK2f35/e2kBSi4BVM8fN+d9Qc05HZEB4RpqvVNzek0pIp/wL
ZBio1NXkpO7EvL8qGUYo358cpcefPhYUdoePapqpvdpH27ca824LZstImOeeVJxNuILOmCC7CHVp
xSEvke842h48FbYl9plZHYXyxTWtrtbKrgiA/5TSjIss7YTdYw18Tv04Dij7eb1lFo9BJvdiEFoG
/mvBibJfQsY9Lt7dHGLhDHTUJdUutG0UYS5jUdTvIrRGBGBOb+NtihGfzbCzbwjesmGgX23XqKDI
VCf5RulG0RIZtEUCk2G9g3NbQIdjj1CP/TKgjxt3c7z8P+IwbPghC5P1ViW+ShFIo8ZZWhdwwtyn
lGYYuBM745qr1Ul5Y+y1vxHOSSQBSj/aN239WBiDZ8pjTipSMkkjrKJTfZo1iSYrTNpRPxubP2a1
gnnMR1WkZdKpdLFPvS35/Nxk425Ve6/jhIpwVPX3oXi1p827uoWWW/suaKUD+ILlIoZpo/Zurs9t
6VXgG7SAfUtVRVwLqRcQWVwzqj1mv2s2BGdcZjXjGJLd8h7c2qq5SGIh1e+BT4UjGUCDwjBQ7/ET
QIg0n79SP6YlWp3810tl30+9hzcKlbyXzx1D7E/dG5Gp91aMHCp1YFCLp2h40WcokFihriv+tyVt
Dw7vft0drxbpljdp2m1U0/MNkNfohFLmCIfcD3ZEwwGy5o+frFksDUPHBIws1fT39Rpi0Yux6wRL
Fz01qZiMGUgz1jvfZFdSLc6aDtE2m26gAR9AVmkz5pfo/hlsngO09oy1ssntH+yCL0Td23AtfXdh
ebGIY/F8vW8uMZc26E1gYhW8gy2t8G6PlqEMgQcvldgs5txeBWEzwYJR+KHDdKsHQRCJiQNxPMZt
oIdZjsmJCWKmNskp0dLhPJUZAV6sFVbbucgSsReT+/ZGCebU+l/Yc3flBq8nTXfcgpLRloWa2HvL
2M2l+3GqI0sIWog+tVIPN5pp/Vo22Tk8GzLQahVjjRziGLD8dhgJVrzmn2rMHHnOwQRnp0DfXFJc
SQHmkRiM99Hd+BpBuZcsMRLIJ/Qny1xoKwQ0uKOBz13LBvqFKuBmAuT8kktmKQv9oaTZ2vqs5tP3
cORlFU6eUDdRzTHogJhseLFDeluNlJVA16V8zK0WchvL2oxDie5+3S2hWyp83JKOq6WHqZ+ggmGK
oR/iyuYg3t36yM1oqvTbXquFpfLWPG6+jHjIpLtJIlYw0fL6uZtC+UfA1lOppQbvCM2cvJVafFRR
yacIK/anBkEsUqVPDmSrpRGggSj2A1kxf2fxg1Qgy/jgxKciQjQ9Z24a/e8LZnSihPch/+WbvXL1
n7hdgko+T/V5UpKMXeyj/bZIXy7o8yMSxY6DyUf1jde6yr6Yal7sdTSMWmVbtiCi6rUpNJAAGvmD
lPQa9McDVljA1bURLE4722G5SS64PTepFCLxahY1LOtK0Meyx88bvlfd+L7IbXViQAy5j2FYduJN
pmB/vZ5ClEL/T4KlzfGTuPu6uZP9DtS7UOPN9ArSAsvdpbPrsQVmXhX6rr8FFqzU3mPsjm2xLV5a
YZKsVAZg0/Ih5/0QcZryx80DgrPO9GfzV4Cu4OhCdVCixR4fCTi4k5DtX5u4AuQfA5FFWcxb82WI
fCXpK8Toq+XxKFcFvSZF2jd57KE4fyFT+KhaqhcomeyBWmjnVVdrXix83TNckIZ1LiSjntgzWy5h
c3Fh0DlPT9OkgsdkNr2spe2eDSK8WpGrIfa10djaZDixQRYZCvoAF9zDjG80+f7Oc2b8WFLTz9re
nZni8oRQayNzJkBQYWHqsHeiQg/xCBa92MvEhxU4DdxulKbARV6bu+1dpLbonsNmMzF8dRxBaZ5B
vN487n8v2O7pMXm/0d6W4uw6Y8aM1gLFVGSBFHPLWqmVCrPep7h/OKxTcUQp/6j12CugmMSVewxD
TGW/Dtrpn9v7CktjOv91H+23+8Z3SxDAudvctpyEyALDYfg+1vjFLr6hc1NW0eYx4bQpucA0OFBh
lZ4iewlLzco49MYGfYVy8xHpHjJl4dqtEKIXYo6JDgwZtwOJdZHZA6tRei0+GwCeTqLof1NSNFxX
PY2eZGp1sEImw7Tr8tHlwWUeQifGNUfFHsGReCvxFysIajP/NXLqYfvtuaQ8UheLMNfrzqDXh+tk
AGucp9szAnjXbb0fuqcDr/bvX92EvbOYiLfxdNtbAAFKs6SQ4Or5Uj89a0b7zgOMwFE1R9Hk45Lb
aIDY5M6XythPNWLuGVCFvOs9iZqg+zBs+GpKA2h88KFtJPlQfoRAMmCkm7F7Ya+WnCeT/AhA/6YO
/PXqs334x9Mfa2sIIDbiXAmJ0GyZFtjrfRe1tCwwm7ky6nLUDnIlLOTrwXT/XX7WJPv1ZA+WvLtg
pn77CKv/3Vxwg3TYmVoF/qraPQHtVuTBAzUYKyW7ZBKaY7WL6sx33p2xGU84qdb2jBL5OVH89uBK
oPp9qjC4grZYaP7LIRZH+3qhacNfd8vXuI0TAx479qvPVaFyBQo1Kap/GW9+nXpzXinSpSAyMi21
jf9VwWEKXhyp6MMJbCKfH+8XUjjggI96u74PHcfaUO6OdjRk+2tpaNm/J5ROdKKh3e40GeCcNDDK
Kbg11w+LXQnGOn8bndQB3xuTgh32z969YwgLjXmQrKgOpNfVdeBSSoUE9caKUGCUkEuao+cZFu0C
5kcdu4enX5kbhTkkCSMykUwpqTusuWZYF6lkwHoFcB+SUohwgomVLogIRWXY9LtPCS9bRL/idVGV
NnYz/iaN4JRNGrK0lcEfxcRAXoIZSiv1+zonaH3b+RxvAd2KUjO6clg9YVX4YxkUXNWwfB8TkFUF
w9sABLesl9aGr17IwRhD1O+hkYZccjXsjrja9Ii3mW57mj8Mk3WQLo69lI8Iehi2NMzRrT1IJl1Y
wGI8e7DGXfWfREkMQKLrYPYteydExnXI5nNehhFJGgfqZyUHgW77JIQIOgXTTPg6Nw2e4xYDqCd9
ilRcKthbPm2rSFSHJc/XfKh+OQi+qxZglC6lcaKUg3uefqKutuXh2BJ65uDZn+jCCOlpQD9g60qy
RHQDIYNWrGWAqXEIDKJj0schW2YB0OxYYcuBcgH8XLEZC0EC60TSWprwoaP8h9qu5KGsrms4Hfcq
hQi8EI/19mGoKGR0pGV/9eQoGKX6c2183G0HDdZZzaRFXHb3zfRJaYvQo6pqbKhXydWTLad6S2lm
J3pCRUURHi5e/SZUVaRRBn/RlXIndYfV6uuMZRgQ5JmTbhoEk3UjNyPXM5CvxGRPkko3lSm498b1
0yz1kkSTI8IoDSIwe9rjhb7VGz/x83x4s6qnZXRFB0avG+vjBL/NmjyJ2u8q6+ttIZHyeC2nodxm
Vtd7vCsZze1Bo1gdIh8jg7p2Loz01A8AZB+nExGqAHhEaZDcZ7Y0oCECWFcw7RKN0f3248lEt49H
h+COi7/w4OwE4mxATnJqaerrDE28xSX37ZRFnfCxkOxRZVqnd02NBQpLN7CGW5tS3n3ByiEqyXUj
YVqhymxGyk1vwcsodayQY9cMRuV+o0AXYdXek079ry4Wv37VFoaPY0578F3PrAizBMsC4E3429EB
KHjeugwA21r6J5S2O81kiGmGNe3CKUYxGXDQMyApsXKfJ7iR3P0mQLTVuFss1iHZDYSsi6clGUer
44UfS8UFf/zPAUwL+7q8CZgsLua/+Cv0h5wmXVfh1LG+xZD45iFjqEOph8QdXDxwwCmr3qGHTp70
ZOjA3fS/v1+VWHPJ45r/KPx+vSnJ1cHnDd7EGdGajSrloBxwAAYhEzBg7GY8453pxQWHZy88mWe3
vyGOmSEK0sWISSqSN7JSeFJVDoEZdu7L1s21lZXSxJya1QsU4/4ntnxrKWfWkMdR0UONS8O1sXMV
8lZBbCc+b97UQzJRhasGbe+1K42N53TDx9/B+njZ2QhqeZkWTFAe034IRzF7l+5ccHts6yDeOpcF
CxEXVSJyao7ldh8YdKui5YqMTZkCj0Gk+4IsxFB5PWm7GdGaZhM4d0Q5rAjtbxNOck/Da9NUatBq
W0PZJ7epjgTD8aWs+RCc/YyWGZjG5Sv4CF7OpgP+ckI1iXhn/2eXimAeL8w9utS3NLiKE1P4B2D6
EC6+2bPgCCfUH98isz6lgYJpv9GlDyeFI1Xh93wFOUNMjXRH+3eaBrJrE6l1uBGuEFsP70yxrIen
6Qg6k3g9IDfADKCBj2GCvxZvyeD5jpkTvs93NGR45VGJ2lpykWIHKCoWvLVFCJCqrgBO++sdGRvW
SAqgOKI184QSqRxS9A7dmOQE3b/1A6uhgbfJl4YgzrAKyt/UGpq6fmrXwAMBwuYHqZ6DlgsYyzi8
IgxJYQv6DyUzGz8SHq2u2ZWv/359ogyu1JWleE5Z8hcUKY5eKJFcNRgtXjGdwHf/yRnqAResNwaH
rVg2u8R9NwJQH58HrLW9ia5YI41MK060HSdhcm5m4mK3b9sJmciBMuserqnywZ9qQbHmJQEhUx07
NqAqjNzc+iIR9nNXvESXlkBk84YC73gqYKCg2qIQ9JKHOmPnKfSDLtZdkaqXrvGYNbmr60emPaiH
7Iudtx1I8fWiwcG6iBoMkaJeNAkyaMFIUruvytDeUGbrlPU3XUxpJtBjhTOoFIuqAwpwcpLklIQ9
8BexeBlzvR8IGE96vsFEf4L/Kbz9IRxj19CqwpSGYqp7zDzsB74ZyRQaDjlvI822UnlXAB8Yyhqt
IA8OPW9M0nKOs7MJsc9ApHk4v9V86gaRLoV5KC+BPRz5/djNAHx+Zn630+S4y+Z1xGedtnrhNGoK
JBHVM1Nlmlbf4VHBJMwB1ipd2Jr5ZD/ygKZKblJ+DyJuMKvL5N5ewQXJKmBL/fUXDrBrBPfcyVhR
/rAeZzrAFA6sjf+bvUjX9yE1fBRGjP5ons/nJp51lpcBNRbD2RUBjIDFS0hox8xnB/nPgmgO5gv4
X71y+k1dUThnkfmksXV0YOv9hgqTTotXJX4HdcfUnamauygXsgdxjFkUWT2CNfCMM4EYHcCIsOWC
9Xwj9/jWTlqj4hJQwCauOIZSnA+rP7knY5n26uGj+0RKz0rAsjm952md3g2Ln2SWKFRqfCoh05q2
d2qXO8+4cDZbf8QFhSRGuEQDTZW6tBl6GhJ7WWETDWxByOSuVXlmsdoPnJdfgIM5sQFdDuWPmlXa
8z0JeJ+gbTTD9c88G/pgFde30fXfJAKHRbKelZIDe3vgXtmVUXItSPqPHr8yrtXqG6WJSVlJR/nA
6bCEyQz9+sWQ3PBlUCNjnTTX3CvujpQ6gfHabenm1NPwGfxVSC2dT4fP2uODyhwfdE7QASWOO89e
OSMwJ10o9E8MqSayWttMPchGFJWX62tQ7Qd5h3dDDdOt6BwR9l9aV7gaUB8s6/tY7Lf2A/ORAcYL
hJshHsOq/SQe2Xml+rFyGNL/Cto5+ljbNdSWdmqRLhrjPHphhfwW8LxmheL80qPsChoEO1/VQEhV
hmN0SrJkovaQNJ5X5yBMFsZ2UBHCY5qbj4PaeLc6jhO0x1/PWRFcVjWEb7OoNw2TAhNsvtHOrtP9
3XqOPyJ3l6EQf+tGdnhfj0dzNeqaVd3c4czxd9woT3+1D/myGjnCtMCI3Kv9KLVgX+yv0VpU8En6
69eXTdi+v2IbNDNxKLUcX1ZoBLjcmUrcKTejXUccCE7As/z+Z5pF2LKfpcoBduv8qyidm3qxrLhC
XitEDIzFrWXBPOwa5lcqCZqZC6BnUmzdFzYI1IeA9E6D+PUl4wN6c3AGo4Xm5jjmQpkXIq3xGUY+
x8X0Cep2xghY3MOUKxQOLuAhwNP9EewpWeYgUQGIrHnCSTKqa6dosIp9expyW9YSoahIeG3p3rCC
5vCTylKwB1o7mPFAXlfBiYp6IMivEI2ScLOB8IcFIngwf6xknKc2N1JDeqePf8YIhvTASDfA87pS
oSHnUrwtUfkSvehA2f10TfXc8eHw0zQ8gwy3osTnW7YA/vZ0rQmA/bb17hUl2AlKW9Fj87SO5roX
kMPhhP3O5ZmoLRI7FlKDwWQNM8rIXrks/wL8bIxNpM3AMF2Usfuhhj3DrdPSACctLJ7lIbQGLQRv
hdGNSxAWSKZ7umyALaOp+trPpcyNgAotbqXiIWiVjfESe9Q0MIijOAwa++abI0vwooiWhyGHn/Hx
m+uIj9zjcrNpWqhQycyRMbVqgnuT12aMr7V1Z5mOX66VsDTqpg89dGt8QAb84xygAVbw+9VTrL3i
HOYEYL6FL+IUNiW7Xg5r/gd4ilweHTMbiuipXMnXUzcNceooSUMTpO4XapcGuSMKeQf3y7EIq8HP
2VmNp+R8M8yCXpkZB50nT12Z389UfQJM5SfvRx1wtY3/8bRF1xIXFQA+jve2wtQD6XH5iYxupCGW
cjWxWyyujDAtW65RmXLvXKwPcseNjnK1P2nV4uHEYx5JksxkiLV3i1JcQcekAw/IGZIf05hyt1ez
6M2tuAnv/E2gqFufJwEx0kkoru3G7Ts8DLjHN+G1w6mggv/6/7o3CYgje/Lp6yyE77m723jP4HKl
DcPQpaYMBNfxVwf+UrDXnAg/1KIDDK59bgHorih86gApvcaOGXd3BV71rMWiVnkZJHtb0dlpRIau
53kj6DI5SI6gPhczWmERE0/V/JrK7cMECUn23HTFs3wTCVYBbTfaXXZ26K88fH2NCwOYiA43oVB2
Hb0g5ey868NJ562jQ+PrZNyoXPjWqcnA7Sy0wNVa11aHB1xEDK7IYv0x3Em2593pgwpZ1udGYKZW
bD6ucuba800hg4WWYbStcUKSfX5Rvk9GN3928kxvoccRloJ/koTOZjFfl+p19j7Cdkf7vW6LrGJ+
n7u3okvbzYlLTUVPYScWeTeOq253na2uOZuNf80ubS5cAqkzo49dBBGX1ZEmrI5uyaxh9VVwxfdf
efNE6rifpZ54/Bvx9AeUh2rZD2osFouHL0alguxxN1eRIdeqQ2rLqOsWtAh04U1h677GOzAbhNLQ
qibUb73g+h1Tv+XQ1DJnhzU52GWUlNWlLz6GqmiH0bpu8phnc+wzZwdg4LFp+Z80Pbk+9t7ji8td
FQhFn5BcRSDwppDKGUhpoXHKaIga8nyciPK3tgUx1NUXUiMQro3YOo/7T5K3paIULtgymmb+uyui
cPScHpPz/vonHaMYsiTJqdiHlWniYB3cZ+IPsefk8cO7tS2dYpoNOWi28i2AskkPEAvmeH9TTdXc
tmKMC2WAbZblGTqiSYeoib1i5I/PhbTqTbjP1bUqs9UZKKZySzjHXFpUxrZidvGLH4tpV+lyedy9
ftMo5IYPYnVDetw91mzf5JMTjaHuSZHwXPvPaV/x9rfx6kIQYTnzDzEyiEruCdQMZ3RXCNN1uDKe
eSvgHgUcUVwXmc1RfMijDnOJfdDotXtMs/CkbfUr75m+tYn24NxMHREVz42om23nCOAPL8nBG7OZ
b03RumwX6+dNQ5VEGvZpeljNT076fjgPGr0PNUcOYEIAm8/A+pDhH/hWQwAji9k0+J/dVYK95FLZ
3nEXIr3Rc4yCMNJnYsXKfLI/ItjXhMaek+Ekm09ZV+IZhcb/ZQlmi+t4tf/6zV0KUTRezY03H1V2
DLDxxfiCbURUlq09l9NCglVWi54h5zvKFYd039tvWb16PGi5vydwH7tpLcNP1deW/34uNPwMx5kH
dSQuUKOv98RMN4IP0InVJNOtcEAr399P0VaOk/rAZkb8NzLQJAQf3a8IoPL8dWnm4njw6FSGfMXY
Yyx8iT54Y6MTU0Xqb0o5BeVVGBLUHiMxpTQ8a1WCVKvkrTLThswMf0oGG6XC7aD2s6wT+ARjkgIc
sJ4kRbHyEmYpbhtN2tuJ/rhyYhymCYxxPEAZiI1ZOEZY5NRu0muJi0KNrKCP7LtSE0XJSxLS1dkd
5Zw5eERKNBg0t2j/HR13zCY7rwcO+oCBcSIQ6vR/HeqSufdPqNTYkP5gYOohq7UpJ5nc7Jim5GRX
2OKYTHA3QjnOuQjc6ra1tmSsrBY5kHcjypIiHlG4Hw7gGjDJeddjEtesJw1stulyD+8IsHeTI/gv
6bGMJDS1yFA+xhSYUnZzO6NxkW229CVjVucLpUs86PbXkbJPCVTI/oHNbxH+vteDgSDRW0sY+T39
ESqcQk9WjhvHaDR9mrWm60PKJArG4+wu/bdMTElEeIzSFrOraD85pk363qusYQ9FcR0TsDmC+FCn
KgTE0XP0LYd1oyxSHk8E8ypSbr1HVF+fhUmTduHSr4CXntS42k1zxRmiWKGRQvQ/jTfHsamyr2No
anYY+Fs+gQ4BG0ND8ZBikCQwiokBo1I7IWwOBZ1/uQBIeA9Cos27HZ1b7AUBTnW7XRjScBDQtupu
iTyCmbilFFDsA1kzmh7tcTr76G9Xv6TNSxju+oskN1ZSlhCuvtNBYLW/RldDJ800R9sAPBlfEbk4
YTvVHS6sQPHPawy7kaNKTsyhGcb2WzSE5gTlUxmMvU6vfBNicolVO9Hw8VLjeGiehVabtlsnEIrE
VwsJmgzNxCPep0kWnM0iophWYBGGn/IMJGYKom5IRrzRtGNgsrRZOrJXMBnI3kiNl2w100l0gUKF
f4fkfHrJ0ragOAMkPQxPexrdWpeUXXsYOhnfE40T3hxiswEU1nkAsoig1NTiqoLTLjXQUoMfXgYr
O64BBG7p952uvMRGlDL3/Yqxz9W2Zoj043KdhhA4B0ZgbjzVFXa7dwRtl7GdM8+iVTh8OlD+NQdE
pn1pT/5WB7yHr71MQJ+6Habv9Sx1GwRVDqR9V9y0RMC8kJ+pPN2o4gECUWCALgx/nHrTRSOAghRG
6z1Yv+4NK6/ZGQYLRawKD4UCM/1sxmeWQkyy15+wRSPkeTKFiMIW1R9L5+1wVb/cjbUs156ThOHM
VTAj3GRGdDwjXlnpFz9Lre/ZtlAbG1O0sovJg2HCZUlJ/nbKzVy9SCWEbZBw6slNO+khBIS8qHuK
S/i4PJkLhh9oi5EWoIZ6uAHx5UZ3xD0gPafGMn4Aaq6rAXIV55+HJJWSo3fMb9FT/BI60lDIBzPS
d2lS6+itMA+n+dWldwVPr9NbaPLIgarsZWK/US2UDy5Uu53bKBm1mod6S2vgko9bvP6HGNVwqtzh
45IMVqIGrlAQne5G2ZdOmmuDl8IGRzF9OOANK9BXPI8G7JpB+TarF1wdt6KvHpGWPq2qyZ7/jHML
e+JKwx4WrmRFzVwde4tFm2gD8wnmu5rL6D6LAgNct0otKk7+tzU7/yOi5bKvyvQrNWvG0nYnCd0+
gpBFa7VhofbrY/sKYzRC1omClJlmPJM21oM2iMThISXZ2DZoOJPBzn/Ek/Bl3TAIdE69ss0omVO9
9va12N0RhGRPXR+swMMKEzjf8MCnjuUf3OBUVSqYY7tIhxXb27AttK+7Pnb54YY1xxBjDSDDX2EM
zApS78x8G8kAdbd8kNpQzOELe2/5RILqpOx3BF0RlM9KqPUk+fXpOwv/4TKiLdQl46PdQrF7dcsh
6wgoZKJpcEWEgg0fS1ly6XcpX41bIbvrbt/KxIob7lLg/xi3rVKGYxo0WHyIgPlLL5CHukXdJ5fn
QqWH94N6PAnQfvJX7RAooheFK5lLABulWI2LqmdbzbGhL9o5SpR9Iwg+PCrCuiNRg+KGfibo88/M
iDSTOCTxRfSYakTwBPy243wEXoS7yY0ABM3imNNftYIEnkbjXtm5rVzXugVtm+Oux1CbaeIhia4f
2a2TK6KVlYgXeFlHVIbDAbmskuZp3/dON8sENKU4+O6GTdQKGllLdG5ze5f1yOyVTHmA5/Cxg/L0
rNtQYCWhZRZz3qS+AjC6XJjgwOv+0JINMZF8b8mLIanXhBi+uHKOYzS5GgNCb41EPVzsqexv22cP
jYKxaHFHB8ZbjZRq6odBA32ZQ4ihFrsUXzoQRr8V4KpE0vEnhxrgGxbZq9GKAXUjmF/EUVZqEbBT
FOGz4x75N4qz0G4vPCCczWLyQigLryuSb3ok7TNEv5Svsq7+Ox5ob+iwsF2F3wa3MK1BI90IA/oy
0SiJUdhhW9YJPk0yAfZUTnn2DC3zhEcFmArAFdRXnv3C5Dlrsug+rzyYmTH9MnZ84Y6BnjlqVbyw
vZTAJ1dN58mhk0eL9YNzl2y+UvujkJw0X5/9/3uIXvqz62HppVxNKbcyUJKQHTNgXOMSuAQfQrbB
jCHhVzxTXynVqzb337dakYk5j4F35u6JMNZOhQtsTrTzNOMwNVJq8KiGkIrwDxKOBNVBKjOP2Rrv
Cdl0PMXQxxga9H+TjcRsY+9Vovd3zHoM1tdWAE157Jm62LtaPOVx9MoIOOD9BZ5lHHGoA9IglM+W
U5svSoB+1jjpSthwrf1zwzL6Ec6Ij/rN/kw2YS9QGRCsST75bEIndX85jpckOUtdTzsCXdmytktv
x8/qoux1TJnNG38WYcE+aG2XaSUQ/o1PzOHaRk+lgRG204ST5u7Rj+exRNYzheE7epXQrVslliMq
e0HGuO4x+5eo7ZmRCTp/BjIVwnG854EhUFrGJz3H898liUTrvVunZL+wCCYzYFu0EIxDAv3qQAlc
A11RVSL4fnLd5f1aFE4wcesH1tiQsoFrxq15rUc9CY7gRG/u6PfPNSBbbpqiVev/OVCeQ8YNIHC7
oYAYtXAEw87ooMACljBsMBIPJCMk4zYifLMvyAApCv2Zq2MYL99G5GxuwfTmTTyXgz6NATM8GZmL
OAHkHpxjKWmKkNbFuouxamEg16C93ecHVKNms2/m+hTkbfmxK6Hk/NZ76w+oTVArlbsRsBWix5dN
B/tloMEfiaMEzR7x59eYdXlCg49mOuZHM8hv8FY//JwjckNKhQu8S6kvLp19IcRhmpxe9RIs6T4R
aRr5/Pw2n9LcVkiVNVaejPFKMvFa3acGHVoROe0fwpHVnWDUg1eSEQtPiobdiZz2ISJfPEFc589R
kcClrHNZmdyhUtDeBLVeXffNfie2hB26ut22Iewb+u9bE4IgcYxP2svvRaSzfjAYTkw3kWBN5pjy
SyVwzBpjHUxcnWk+1bHYXNzzLO53G+gTe5D3iErl64EkF/nwFraLms9hXxT+DNzJDgRFnaZLL12a
sYUVhFiBv05PszHeNAFbXzaGH4zFKpXhOe2Jd3Mqwh8Unmflty7fKn5hpeBNte5FMqH3XFy2JiNh
wpppgX2NF6Ae5SeVvT+xpi/hTtZ0hAvScpzD6E8Yub/TF4/iZKsq9QQ7v9LmgCCGGPrRlI76c9pa
nKBl9coP2mkbFqWJuGhuFyY0/nQZwMoq1+SDz6SoJ6lJiJaMJ6ZfpZ54dRS3+TzbDTHksl9PxCk3
IxsLpk1ye3cXNpSS3k3sRnaAGuljd2du79L5lTyK9fjsj5d5wip0Z2F+WLCklOb339Uy6mD20zsX
9uKvHSLbqZJjDHNpqKY8L6PRNPcd9IKcTgD7o2FeRyttS1GaKb2ChzvhrkEbtYOjU09hJJQvcOZ/
W9FOEq9PiJrgpHa22d1x5peEhFWW8dT3Dn1D4s4jD4z73gSH2KqVTYtHzsLvDVWCG0bmDvM0S64J
YrpiEd1K1bvT0p1vGBew+RCvk8CcziWAy+L0RCzHNbGSZa1OzqGp2WwlwGiXvuVSoxro6PlY7RWb
Egz0r75nWuklKriuxBMwMca9SGFaVI+VUr42rAYT6GHrwtO7nnij01gezrJpeYLaCaYvvG6vHfaK
tFmyqAwC2DzO7mzssA/MDVZqy3mjHlNK4i8ZjuYNp3h5AwvdjRNxtK75Ex4cm4LUxenKthCWyePK
EGS7/h533tDUfW9lBkBy1Lvy81bmD2/Zw6dkj5ZYFXhjYW7rqy+IUfxA8aO6UVNhn5E1zN9tJyCH
UJ/eTOagY772k1+ajboPol23ZBwYcpQHyVdlf6yjFlPCa/mUGKFzS5Z1ua51kPMzFV2Q195qf9db
sJB8cn6MQbbRIpYAIQRkMJY5eEjn49bDPjqH55YwVuv5aNGL4KSa7jq94JU9iM8hfD/ST204GHsT
Yg9d5NEU5hsQLLA7nfFUxz1JSX2GM5+JAO07negyTCEw5B1FaGb8lAYtZSFG/2IeKid69l+458UE
IMjCn3AgghM6T2DTQC17dmp+NWR1aOKamqWFTGLhXnEGQuA96IXKu/380xTZnVbc4js3Qik0aJ2a
nPe6pBBcVsms+GqhObaw7j1iwuww1peRM8gO24RHlqf89LBs45sW43qqAejM+IzhK9UlqiLW+/74
k3XuW3wHLmPYFJxU8uxvGnayQGvAqItMCoKWsYXe/Cj4hbVZymkUailFjvYHHG3J5Br6wNQdjIVH
BW7mhCiD7RSraexytjzaVQhizZI0b7PvF0EvyMvXa9ekbSkJSwclzPBn2JZjk+fJZHXCbtz42TWY
qyKPgB5UQuOCo2hceFGy9PdTusdq5rHGpKio6qkz9dJ3TY0mzfu54zT185zPkBkzuB+0cAln35Ty
gHe2Fvh8nZPO5vkDrO/oXvfI2EruJ+/p4tTY5QK2iz+WN7EN3aUocLEbBItg0x8+E3uCUIYQLfBJ
oWU3QwGF84Bade5Q0ytxIcIbaJAKeioIiSCslCMv4BadjcxuoQDgm5MGKHBXzvytC6onNUMIBcDa
JQ4iDpptoRM710obVr2RbXKW984IFs+NPUKZkgecYXZ6csmkfdmSdfr9H2EDgGscOgO7MiGOdjPQ
xUOo94H+v/qogLgEt5q66eWQaKSCMPVYpMAqmkQUA2++fv5hlAt/dHLctbOdz50SNK2AxGC3cKv6
ZsCq0sV0Kc3tez77MFwi8Yh2HimzUj7e7w+SEJ5EhhEBslp3WtNeITX7WuvjIgLmGHiQOE4yQ8r1
wj3yEb2Whd5ewUZ2LsAGP9MaBj9yMOYPVfku9zH032S9QJ1Areb72eB9syVYioAP3C9Hd9QSOhhJ
+9Oh/v14rdZCXLUax9/5Ofrah4UtI8W7OrNaLbQn2KEIe4Hd86xZXsI9UbH/83xiKQRdb3brPPkz
DuTo9QbbtIBVamipT8Ftp01m9z8KxLVulb5EzKOsJG3asej5jMyHgAMQL2Owlem5/SY4Jra5m0fa
Hm6ZehO+3q97bJmCWuAbw3qsAfGcLsypNC2uQk+NJLNVjaxxdL6eeDjg2EBct/s+oQBFBideLFqd
QOM7FRaojoSyXdAHqK6lcwop4U3cDwyoMTPluc4mBpgQDMVVPgUUE5AeafjrG423cWdWn+Lhsut/
0BVxXtzA+D09ETd12MnbBxfu0SQhnY/gm4NIC4i4R3h6/zHWaXCg/919xtveC6TZHvZZy7Kw7OIV
amh4tu0feqSFSPUatasdL5nCL160t8EA4lYuvQieQzCmwOzH8fE1Krazawyqpkd8Nh1ASzHf6twL
/tme4n41kqPBteUsMDltHlz7TRHiZzEbr+gr+MNYy/YEoBiWFJLgiyMtawBydwKWSvd/5rvZ6GhN
hGqEdQGxNr8VMcWb6chTjAcpKAfo8VFGz+j4T88OFD4FlsSe1acO6qo/mJikJ+mFW01gsTs08cLy
x6B7RXdByZ/fF6UUx/KjDlQdI0AdATI6l0FakB2iPkrJ1ZsnBexgWWAvA4DnHUnyHRxKvhhRhMPP
PqMtW4JyQFe2Ih4bTueTidYb6LDSNQ84f6gvHfjTYduAqci4rNbbtb1H3buUg8yu2aedboJGJRKw
gManRfKFivhKMqEwhKBhZ9KqRMH5T/fdSgeD6+ca8crSRfL6nY/UwbzYfXNbTd5e+HTGnC4E5G9r
7gRsGglKNck=
`protect end_protected
