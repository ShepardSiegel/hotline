`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
he3D2OSbxrE+4ttnux1o4tUZygr2QXNxR5YV25pvCuE4tFagOcmBSPHocGW3kieZ32cnpSE4UPdC
LU+TldnJnw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oASYliujHRqKb3JRwyKr8IibLaR8tbrMNNlrUaMLKL6dY8d8CSgJgvfeAyNFhpcIaTd2qLyE/7kK
OspM4SD0TfGa6leAMiBZmOOePfCy3ISEbqGsiWHP78WGLoPZiDgUJCOCniycY8vKBuDPUyA9jQBV
er61hV5vW3QD9DZ2Kx8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aNO/diRAN8g06wKzRRaTP2HG1p78XlJzsq60sqHxEZN/D34silgNTiqzcqpubM5bPGmafLX3gFXs
kK9L91DRMfJICmXF+Mdil70s7LPy7hQOqNviqHyJPfU5FZTQfL1okTscJMfGhcTS5UxsTUqwcBVi
xFrfYL3qlRfFAJuIF84TnsTANrsBLU9GN9UII7EQ4VxaQVYzg622DdMcw0mivSAeIOKp7CtMru/T
EWby9i23VsTO7Kq5+pUcxEE1ISm7PZPtCRhmX5BCkRiCF9499hxgh4wK5RS2zd36KDJxlM1xCm9l
atBvYUU/C5JEArWBM+BC/1Nx4mnhE3QF5RX9iw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
V4JtVMaVdmGeWzj9BCj7xucSNwIzWxaEViEr94NksRPaXYjUepw0oYZXhavcfR0SiSS731QE88jt
tjXyge3zqOKw9Vg4wOy4WD62bk9kkahf+ZdxXaDLBgO5ykFGD/BWhzeczW1tphQJp5CWR64owL/q
2w4qHiF3Lv/l5V5H6ko=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rMnJnjnru4G6s1+QlFbV0JnvN3gNajZEHo4e0WpGEqcENBw9uuheSCZvWeO/pptPb+SwGYJJYX1g
UG075hhWJygVF7Sbf9H4rYKSbmj5rs6o2xuoYgCI8YOxUkDX/a7AXBAu2lA4NOY8uepdwjHoEiJs
BJGO39qBNOyVpvCayquRWbWrpQ1WLe153XCuy++PZcAAIaaNBsw5kSdBe5HVal9Wef0vqn6pm3ge
vC6aqtszEs92aSxEjBeeUP/7iftrA12z6npQyRhMN+rd5DwahBFF0RvJA4/UslPQ2wMdeopmfL0Q
k31FiJIZDWNas4d8Iv0kAZQctP6VF2Qy2Iym9g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5248)
`protect data_block
rALRDoVNCu7LdFyUXcWMjElf2k1765txDoIGBG2rNmYiPXeFENJcusx03WwIPdqGJ0SgQva/uPBs
hqVC8UfzFDz15tkrKa4Vq8zHMKrW/z48Gy7x+WtKDNk3Jf1Lli0CG9zh4wyFEkbbFObP9qXlpfbY
lJCa0N9ctEkXsh99aBEHlsw04xz8kOvChfMStlXFxkcciOX2e27S6EUprXi0MKNwaru2D6kKUD90
oLpBaUlaAOV1Q0LQXujAElvk4z4O6YXTDW1vLEdukoqtgDFTE1ykkTFZfJ3rypknp+jCzlID6R+2
KPYxTXbp4H0hBBfLIrrvEzRiwlvRIxgefFvkbh6yx0DgiRS5L1PTun1TGiABJUplAl8/v+PZ9Q1Q
X+AO0Z/UFU0Uc6VXFGFEwwK5OpBO+GQ0CeoVpRcnxwPKdZiizBBYh3SxRr+AhDwPV7uWD9k/P8YN
fibI1h/USeBzFQSoxfR0L/VXaVOtxo0+EHKzkgDdKPGj5BB/DGDmO5ZbQn7ulIvEDqP8hhU6soXS
tXWO9cmWawI0KoD2iT9rHCZDxwE36EPyDbnwioTdWpyeIWbpr8xlm9b9JD8xHgv2kgjNwGcdD+uO
oOfrzBTeAeRM1qgFxX0AaL5b7lA6NwFX7UTV9QmsisPfxwOtxIcMcG69+Eh9DPqa04aoj848cZH9
kcP/vl0T9ODZhY3o/KVUHBWJk6NCuOmZwfhzsf6F3/nfB9r8gztB/6kaM9vuO6Glc+ju2gFYd+jI
aHDxPz/baIMoqMcdpzyUwGvb82F8B7mrjCLBVYVCNTCQZ40FQmqMC4TIZpuE7il/JFgEdwLSW/in
Lpr1u9MZuRUzzUxucQuSQiPmJH4CD13lg61OiO4E47LEtaAn0VqQVt/AYb4bsVUX2heEcPMmyJkF
FdSGVj8vnP12DqTr6kKLWO73J1T6+IsOa++yIXJfjpK0Qh7APyZklsdeXQnGZYTP+mQ/lySU9Q1C
qHHJROUp18zEeS5WjLjoRlQTvqbHZ9hl+zvM+FCWfDvDX+roWC7c9cJhBFe81bwZi0kP5mdhXg0W
gCSoPAKz2syzsv+tMXacRqCgQypAbNObGUttZb2nTF5ssudpghiQtnWcpt2EQmyRe/KL9sRpAi/1
0CkN/dpL0xBCy2tuijpqO62+7c15degB9u84rFoyieAKnodk2prLXNpIa64sOWVNunw1fI6fNQC8
zAY1vbSTgwJGmddBrlEA5ztQCZI3D/I+L0O3rRnCFlui2k+g/IVPao3XNAqi0qUnVkQ7m/SEm11q
Qodp3g2/ihQaF7DHvv82UhIselyn88SG6v0W/u38M2Z+12x67L3vV7FLWWXD4Qdaq8TMltQusDWN
Aq7vQss6V3qlS0KMWn72IPTQcsCupXGRYuvNak3qvO3GpvT4v8AA3qu8PoS6B0LmhCB4Xs5D4Egc
EJIhgOsAv1i3u3Vqds7N9OXxv66YrA64CHJIWp1aAg488nmHUh1XpjQPpWQeYwEdK2erViZbrYN3
1nuTFZZ33cW21SPsldK/Vppp2ylsk+B1S5v/RkDW01xEHMqzf15nLuWS3+yN5rIK0NF7mRcDS2jO
15/ktXthEm0oklAcf3qaUzHX/JXfqkzK+JKJlklTt+RHEW2k43O7f9AuNU8PlajhK8bkbaBJ4rnf
wF/TtKSNrgFbP15y5kvF5t8DRF+FDg2p8GnsxYwR0+0eCJT5bnRZpm0N98GVBA1t2FSXHWoRe7SN
swClYWqa/PL4y77vLyyvriYm/9/2Gr1N97WNQd8lIHNxyuBWGtwN8uot/rzLAZ8vahHZv3epWr7V
Hx9G9oHmBKTR5XbjqfZ0UEhBAKnyfmEG2zPJpsWk3AhFxH3tDTxTMFRXh/tmd8acNhV5HJcWZPS7
eXtN//jxgDEMfQ6yX40nLk9iaHSJIPJG1WFsU9Ywpl+apgCy/xybW5dSvdtHh+9ciI/gSv3u+jjE
hSGhuUrjpR9YG1+jpPgH1UN6ocCcVZI84QbAVkvJpgGGS5b8pDgNRLvtPrQgnzEu6e+9vrE4A0a0
xGp8EEpxRRRu5onAm6jaRky2EdyY4hAVR3GlrPeYpeiuCiCGzDKQiTuBYvkLSWqvvFfcciWNDBJS
wUR/pwaAMkxqqdleV5vkdL/fa7xOGEibgTGWpb6cp+oiEy2KuNyRq0mhxHoLxhH2pEMq2bcnvGIF
wv4YwKdDPGVuknAbgXbbvtb0fhcfPjfbeV8J8X1sMfXzE5TgoaPrPwjtFFIinEK7/3jmI34OgzA+
p4ue1zk1j76cg7wD3HU6IH2+4Bq/rsQu+s1LDkTfGVXbhpjqBjPn70wQTYpmYeZEpEEOC8UevZd7
0CQUDSDGkoLH/bWv/VvDLTizlA6YVyKPyJDku69JKI+IWVuakeG9MPa5482sB4PBlgRYUEM0wY+3
5jR0JvzpfuKjORrgciUk4OQ+EY56ICV7HO/bKaw9EyXUG2jgo3lZaPSz2Uo6/f/HqL58omLS8pDf
1BeMNpWP4baenJTKTy4yalGF08tDlFG1J3CQdFDJMQeKZM4gI31e3VX+Z2mQoN7wH2M0z5ofDV4y
iv81iZCuvLCDfT6KLX4kRGe+4/cZ36ymmGgbZImdethIiOMFAHAVPc375oSQop9PAk8rPrESZS+h
MDW5HwCE6jH1gZQpe/RxSxgihtNus7sAsctpfWJyneOHbSSANU81MU8S9m+YdzamoMama5FH7khm
vMOeb08tyffsr0ba5ZP2NEwqU1b1rs7XKB4ETE/6bh5BySlnXOm5EAqIXBmDiKfsf+thtGcGMuHT
w4iYuginljsWGn/mRHeRELB46JBxO9UCvunOzly+OwVG6/PgQs6Ku5VtniK/kdBoMCOe4B215ccX
91wjJ3LoujHb7vGHQYs/dtic34WaGxpfwIYBsu7Tjxcx3H0ZXEnI3Qfajd/i+r9IEq+d9oERKnNh
2uc/ujOKqefimV81eE+mCm1EOBzy6bfi73mcaWdxWXJMQI7UuQJq0LLFOWqHUDip+lu6sHpnMtzv
DGRmCFQZy1sbKA4UIpXJY5VDNt+IOZ7HfH/p48/faBf2MoD4MIvROIGBZrVmDhSDgHzavACy27lY
SI7MHt7zGyO/p+btv5o+6GbuYOMhmnHOPg1apYJwAc3lo0TRmNR1CiKCVeDU+z7HpGr8G4q0siPm
jyzjeZeuj8bDoGFWFoEWO6Ld9Q6liJlYrFA6foJG+xEYAdB7t7QFUdYdPAmhXFANuGbYG6Puicjh
kndJ+UivZqBjRV3VR7QLkdnfaQ5U4wn2k4+puKD/aUNWgbSx2Yk54x4dgXmNPByvTQ/hBDh+QViU
BLCi2Yc+h1ER1d3MnhnkRYGDovVE77vVb0uNeHz5GcZxJJK/KJHhurWWMVUhOTHe4H6F7z6gvfwk
kh+jajD7PZRiPdE1Nfskzys4lcnVk2o9eArCp8RsEuNvMG3SjLDNrqcX1dqlP9eyWust1aULYLbZ
thp5eQKcMsyTbD1ZK29YwkreOYJxoB6u07oI8Bix0Ai3c12ymyQ0PKmb28CzJFrXScEVwQHVyyPd
p7R/A2oJRk0oPCsal/08yXB+xWx5xWyIv7NIDsi9tPQpCfNrprpNXSO31z7R0jb7Ze1Rg35BkKvM
drlUjDn/l/fESTN5VRa0u9fDKr592boVOcfck4bilOJQ/uREE0RgHI+3ZmVTQAYHzZPLxxgnNvhw
t754GvPOBHJe3KNlIneKfMo3wckLgVOqsGhZjfrL/7cqle++MKL4aJOveJTIMV8n5Ze0/LRkfLeW
vqcqauPpogDNH04w8Dn29q8aOlcax4wKO2NSUEQQNaT6L60vtm/hexAN+osoN1yASds8EqaKT1jn
FDiM4WllyOTSUFYYDFnDaQD3i/VN1Q8R9xtzP5xPDYWlTjX4f+AupaTWfymAivEL8p5Sm+i0u4PU
jx25YFRbK4Qoon/r385hUaTlnKQUS5ald7jNKmMMLoaA5fikHIJ1Db7w6hJEnfuR0gZmj//H8pjq
dGnocUiNCVvVoYYIYMgtXu9Ikh6BsOxb76Jr2bzMXfF9OrcViLzLTqU1pzRd6Cwfj3i6ug7rN1EG
MLfB5WyuKxSe7C/0MWpn4E3Yu9E/ma3jyDesvoDvI/u9+pQ9rN7X2Qf31gyA6m+FndQcHquuiytK
gVK7yIT9N7dxnEExX3zNn2ooZFYRLWSIRCUmu2o3hmdUOUKCpH7efM7loRafAKQgUZV/f7c3K673
kvzQy37ZhtpwBq+HFOHE/3AqzMTN7byBVdvcDSaLKtkWX1Y8j7msMsxw2uCY+rzpoIiD2U9m64ts
6LJcIbyKxwwgXyG7w8bb5PRu0/nAx9kE3kBQcJG6t9XBEfcfEwdw6bYGCrETWNC8OQ6BeRM9OIlL
aN9mDgSVFewQQLDqE/waA4nQEotTfRvi+pNB9AR7QHdlbW2xvrAgrUTG/wyOyABvv3oK906/8Tn/
rFE4kmlmh3gqlX6vL4uDmACSyKjOCMsf5VGCzsTRs4dgArTBn65prvbghtO2EV2qDk3K7+GAJDwd
4O76uzRL+dqUIrnuJElwnZ9n0PY+giAQmYjgPi67pRn1a8qunmJECGWFYm1xB3B3/Wx2vPNdjsmG
hfJQX66eDvRInfzxqCK+VSjFIRa8PQ/LOTmmaZjJYq3EO+6ExeRywiHi2pjliPuH6ZdEToHmMl3F
uZeb67KrYiPLuDCBCUYP+ID7HBJEcEKb2ybXGXnIxRpkcN6aCvcAn5nLYtwD95CTIEa7KBsaQ6fx
5QurJ+ov7LmgJ87JeZFSoSrBA7EXOCNS53uP6fcg9qJfn6f49LBUbYNxDxgEN3uF6RlfUZNOcaWA
tqKW4uNXSw9GrK+0N97con+Ou32FEkLD+OKaKd7yelW+3BouLkRB4b7/ktoiuriHGC1PzQmlPFlQ
eQkLSMPbPT12E2lM9HxIdgStDqQ6jRYDmANHRFBfCRWarL5dv5sLF8RM+9ynTm1odfey9sNJoRkZ
Q3K+SuVYIMCopxLQGpdKmZ/N3rDsrV3lKrTWJsPRw/0xXM8y+VWsfTUUbKHam+UUoVKyDZN3T8C5
i0bGNIcPS0Zmdb57p6DQfthDmEjbNHj1XytZ0hhRezLf/TShKwUupysyXua0VS0hc7xFR1ruCzRI
HFVbaLJvFN3oZa+XF7XPNIesDUV7a04fNI1S7MqwBNRTdxJnr0O7QFQqGPmw8Ydfp9KRWNdCq/GH
CFgFL3l3GRglCkn/JDkPbxNomQgEkIl6Hba0OkfJnjxB8Pn2HW31zswsQv4aCqk1qpf1Z3n9FCQ4
r2k3Dwm3v2sz1FWMbjiJulqC9BLyEQOqAw7Vcz7u6maL5QKMAqrYDWcgfj3bf5HTQO1+QKWxnpwI
VNQb/WUIsrKQILzoh/uo1NJs5E1TOfIi9xpqE+wEFKfrk9GJGPIljsIzMmxKftzTAIl6AD6QjEhY
89Nok5ra/EQpQY/tGhO+NE8p/CNfduTW2Fhq/1Cm7UhhHo1AoTURgcmQJW3VP6GK6J4Afx6gHhlJ
sbv8dCcExAQ8jqaiN5yuKTZMCxNH59RGFvxwAYfOT+ZbJZeHv83vZq2/B9xxRykya+TCUr8PgBAi
7SuQHPsh9/dWnieAKH9FO86dE55BHc4OjS7qsT8GZpnjAOPPdyWF69pcuGBlETSrFj9Wwg8to0MD
v2+Y2vzqaYgvxElf5rk101YyiDVgZDr3Hqch4MVPLx3hWV8Pp1nS60F5Z5YxLF+YiiyPX3F3U2Bq
4H42soer2UsaK9f859wvKMFFdPi0oV/slmkwDYM8YoBUTGdXzAMrLH30sLBqaGVPNrhZzVzd1abv
qDFizSPoygJxS4/iTOAc7myb7tkZJmvn4AheCInl+Mbz9melD6uYK7k+AYPmzPj2PoPtQDQkxGQL
F16kahibjs689ohxIhyj1+us6JxRblqkCKPUIjf64PjylkY+daojn3vp3jIy1mKBTEzv2e3vYK+O
cisrJumLeTsPyCBL9JXXFujYgYq3ezSe4N1dLDXDdPoV+F9ttIg2QBnSztrcLTOGPObNQt4jC1Y5
YRAhgg67mEMAdQsWYvVxCQI+393ovm+9f5RJfZgIKD4Un9pn6F9rJbAAXW/v4ojAKr6ZMjQ5Tmwk
S3ShV6qzmnkpDHLjucRUAQ0HacsStE56i3zpe8ih+P/IiEAACTGIp9oT7BQAT22Txk1Z3eLMojvX
gsLGyhmomWyup1z5S2Nk4okEkyw/yZ78zuBrQGxpPH0pmmKzO/Sj7JsHpa947o640taGDN2mEJEI
8ERxyFlphAS9KPMCq0XzkNCpNrnUIHEaipbFe54twe/4BJ5RpmYL++rG2qGd7reUiVw3swC8Sw4d
jk4MiYOgKeaJTFINZcVkfAtHmcEXVdTqGPD+VHpsIGY5aBywJ4b+xf0lQa6LHwbcfD2XwyGawzpL
Hcibdf/g8iGBZjhexhFbpbx7v8C92NfhIzW1dQPUTQXs7WqvrjPU8cvbHrZ++cqSnjxpWUKsuEDr
VtBXkiXE4YF/r/+tt6ncfqvfzt56p9YSQJFWsQaa9h/X2JV1ABgdGNFqeFBE17O8sRPGbWMgcvAO
tma4FvQwovMRgQ2CxQwrSXAGZeDxy+ZnaOgE8rYSeE3Vkgg/cPbbKOzP8czsHDN/0iR8Nt0LvBxY
/8hLN2MGfDdr8USp4AT4/ultxE6bWeIW3iJY/wq0fLto1qQvCFn/+M/Mr+RFqVUle2Tjc3LJzykk
xkd2opM4+FkPWEywhoofPeCpfsh3ASNtZ6r9OTS8yjxwwpj5LFkJakmXVz7lUGdCYFrQG9neozIy
0XMTnPXVIJ51IToYvTn94r+lDr+Z//fKXHk/wWOKYpPBUiPYk98hZSCvyU5JRBvX6k9RrAwH7oyQ
rOJoq+unloMfdZmRUQhIGQ0xTldmGmXuoSHU7zZc1mXmvU+m7mMc63qvL+gXJ1MnZWnmbmJcMUUD
TeQebQ==
`protect end_protected
