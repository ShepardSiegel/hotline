`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cpvtMwUGXfKspP+STpobBkjqInqQ+UVW7diR0+HZzGdtoSlJE6+s0qRLOe9RloLnXj0xxcIkvuVq
+lFg/WoEaw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VqvzYSZmEj+6lXbWJuzM+VXgbWVbvtDDZ+JvR192N41W2vxxfDYfhCLF8uu+OiVlm2c+HkY0hCSE
KLpHlmVr2cid5Lb7nA4KpHb+n7jrPrvw+XspMPSjD0HUnGFCzVa8D+G9huiDSiioIbyA+Qakqp29
bi/ITeGVHwU62o1PvhM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Rpzlj+yAGuUzzPWNY/gBJyxWK3BWwmv5tY1j4osAxUSYHPPzM4Cq6GdYTzkjikDA4Z0MvRHwnknD
tNKV360SIh+4KIUSil2UwXSSABsO8qUYXd/xmSFXqTrohHHJ0pE2LBfhxNnNkL1poEN9NyxpaCjg
3C1DaVhsyJA51lvHY//vT11EMrvWlSve0//T4oJ6l+UAkrbQOZAoOocCDvmkpgsUTSz72cWo8VZM
MwS0v6JjQ2DqQ7xPuF9CrzvYPM9TS3mcoJ1Qx9nkD1HqrOuuHx7XjwzAPk0qlIlgN2wD1f5jSAgW
mIFdNVlkI/6DKCnozluk8dDe8/eE/I8HxlE/ag==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
V2q1pQl+d9TkSrYm8GX/YMEptRWE8e2ZWDQQJZVbTCLcF7re6MkBFjVjAhAXpEPM37bOjMo9Hiki
HTjh+fkUvO9m+fHMyuJX3Q+fOZafyrFoEc/+rM43uSt/FCSbLC8ip3sxBfbEorXqFD3j2m/KzKlM
+2xcFpxNAqnXtv2j56c=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XMNz0xTQ1UW3hjU895eBY+GjB5+QmrflOnmn0DuhP96Js6u9UFLEHMrGmpFBTZH9dGtDjv4jMC2i
+KoaJV+Bmlh68PBx4B4gE1wEu9rsNi8rwWmWiZ6Gt+29mWoYs0LDaW9obnGQbZrrrxbrKBwqiRJe
Hj+hl4wE2/DrdzKo1vpDvPpsIDgvXkEjfswGe8a7hrTX0ncxsYrmyOZ2nLy5PhOt+7Y1QlhTKcO0
Pcth6cAs6J55wSQk4plqM/4S2qekKXKyJk1Ry7e7pHSITHu+2W1iSLHeedooZgnRkCl3lEzafiZq
rDM3wGa2HT/rjbvn9YivaKBlPGweLMSnOUXNYQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 42640)
`protect data_block
R2uelMkeYySsYhrLb0ryYsHIPp9W0nV4F+8nAsJeKgcoPcPVTpR/yErBs/hyOewN1knf1jmTFI/x
OrUNH3aSOuonrsqJe2RpYizdd0Zxh/jzPDTVdUKcbpyO6MAdaydmlCc2CzUTZzAxO//d9paLOgqi
qe3+HdDT7Y5eVUVGYv3lxplTU3GxHSgNvUTs9kjpWmhawMWiJZ5/3XnNFFvWWm3CvRK0HqbMNxOR
iNsLWCtdVwzP2gAR43E2iOYnFA5EH6AmiwzKIe1Kh6IvaPjUuToSSIofD9DzJXhHxSO+6MO3OHia
F1V7Z/HyKD6SDFTOuvI1q6IlIfAJ5DDY2AgfJtZnWZGcil47hWCIKogbkH6eKwiqy84C6qxcKtGD
0wHLICGP5ODcTyyHnDCk8oaAHlz9sd2DGvWsMwMas45y5NqBLonuzztXlRigSkDNkgLrb/eKDR1W
W73mkKZfoQ9VdBYk4u6nhsESVAeTykelZguHCytJsmT9ryRjFpLh6ECzbljvunikR3a75iOVSzAA
c+plV5oO2mEe8HY09ZGcy8lwc9rIOaynwos2i9Bau7HUsTkcA1LpvOLpI5VYx6e4kPudHHNaz1PR
guQCSo/Ew3ojg+YLZYbAjChx4ViL9ItSab9ZXD+H0T0DEwZt2J/il4CeDDhJXyGDWN3yAi4s8FRO
7jmmlVx5JCPD2FaA9q0MbE6/hjcKAhkecLaz2XLRBKdTGPlKv8b29u5KzbQmAstuxuSBSaRkBG2Z
I0IGJdtEVVboTj+LAL2cCfonev4sa6JSp6pkxLvf/oj2rrge1zu/T4n0GRlK4N58JOYm/bzRMeRg
BSuIn1HlvqaefPdldy+cRNScWp/Gl18iuKFz5gp4IK52Qrvrnx1t8jt5KBfGBRQZ8PaszORqB0MN
YkqQvijEPqK46tkMh0vRJfxpBrt9SKpFARA6S1ZkRpDqtUOyfLz085OPILxTok3L5Iy56eZebTkp
HPs5B1BJhGf6BDe3ajwv9tenB+FNkKksxBGK5gSnh5hTwXmB7WmrnS1ejlsIbhItpL1QBcKyWgOM
A0twPChMWAYyAYHZLRs5oTGmz1rxjZtBBi4ES90rH1aXl5McRzrc2CnskMg0Wa3c1wU4413fZC4y
fYApbENWvgSlAWpu2Nlnvz/k39Afsis9Mdjlr0bE5T7Hk9qqV4vsgr8xcIahEqGtw4gDRtKCMJg6
adgTLMIfXYAxgc5Lu/MF+Dq+0ItZ0Vfb8gTPDIl2VvZlH9LnLUlSkIwOdC/RaE0x1Eb5CFvyTfIT
1Rh3ZIfmxn2lUZgQcVs+Tt0JelTkhJx2hfpDcN4nJT5h5yCUQtAsBBM8sIcJWiiy05Ink0u10t6Z
n/a8zfPN46RhtDzMZrXClGZohOQSirol7B77yauJzTsk1iAuvKS/Gd3VV5cNi8Ra479V2lULXHg6
Pm0F5hBeq4aM4rFpNPoVAbTnVeR/fXCqdrKCDM3to6nU9HW4rvcGzIUS0WuEvRd5eoe3NF8Oijv6
byhNFB/flIOW1Ha+wzMP2JKMp4KOm8z2IJ8NdBXqZWm6riFy3aEm1GQ4N3ndK8Kak0V0fuIdw+PN
3uViFlEJsno624V8hsskYYClduwKBUwN9v+4CwjcMsoyouueosqE9AOtNYHt3iNC/6SAc9CqPp83
pnpEMM6sNw782eCWS1NCcjD5Vq3lNvIU4gfnEhgg9N1B+0dpj5Dl+KuLO0YlFfnKnVgk+HaqHwzy
MxQgrxZ/aI+ky3uvT/LA8Yb1ftjXrux6e3WtsErhtqOUqIO3Ly9U4vGEocRGCXac1TseRoHNE7i0
mh4Mvg8Hke4ATPV1qAu+Eigpv50RrqMBcROq/0r5XnlHlCzdDpjUVjeK/0aJWz1WKBKL2/MgyXmc
WGxdyY9rwK/Uom3JCuXpB8A3H+XbyYyTHIP8l9ALTY5wlMh+9BIVeAWRp/SaqFnddPhkT1ID2V5o
1aLQwvncUCa0z1NCm9SNsWxIx1QznQFpbqctpaD3oJ1PZRvlv7SwRdloHinrJhs4yGAd0E/EcHOi
Wy0t2B0+k/buZzTG2FQBl+TfBHgg/cCVXEfMve61MtfB9OV1DO4YI2EfGAW2dRcd11kQ28WxkgG+
Q+ZzzZXWDQOvo0pTWnHHdS6D056gEgNIxhGzjSdskObCwr6IwbHcbfHmRP5MmUa7tVieHuXas9Ht
7u4MYDix0LetqaEd7BGw1jvMmAfjROf7cteRoSOa5IwyrT4nMvHguLl2bD04Z8f92nQAaphegkjZ
S7/dyQPn4mejxt/xFGswhv996hN+/rLpkOSenfbfzuw6UCTImG9gNaTdD3tp4MlRzBgBmqwnGkuK
RwAfP0ciz8y4ANndfkB5ge48VnC8i21iU7KSAb0MiYpFvrk9cAkSyHrQD/gKC/NMJjfgiidT46FH
qOQnG1uOSjrTuPTdjxln7N7hKvQgREXfmveZia5RmacUtd6UEnrL6WNR2ZzLsA9zS9aDYK2cWaig
cdEhISYlanwrJ7KzX85y/dIIrPn53YRAIuJmAiqR72r3jGP9CJwtTl9DVTyhSyXhXU9uEoz3FtuG
tRmWLstl0MX1a4F/Y9eoASgCO34nCEF+zPqlsgHafpQo7qw9ovAQTbhxeIS/ncH9w0zZQMLCkhEc
riY0SaGbsAq8WslcoQICwOMMRiqfukVkZik+0kQpiwdyJJ5XksZqkXd7Wtgqt66p235JoGcPq0hs
VBa8BnwcrXVYE7TRYHOUlQSLWPoazgg727UsSdOZwVxci9AaSvs1HkkMtV/kJ97yCia/W3ZMuKxA
dh6hAf+MyDcPDezPkXBW+v4uGXPRMWixm+t78npKtqhMXtOZzjLios6+HCn9k/4Qe3Ienf5t6I88
GCXpa1gGdHRpVNSed4MVQeiJTeZpoyRbfVLS0pIfgPFvOCScNXaCP4yKtT1Edp+P3MHAuGghvI7Z
5wrOuGET44/t1KGAkKegW92oXS750emc5+P+KSLih9RtYGReg4hl6tT55+saTD9HxWVFEIXrl97Y
4R7YGzHzF3+tNfhtkP4DbyqmuRtl5l5NwF3sNpohbb5wNccCUrydrMkB3W6KLVqk0vt60EsLTe+j
p8eh6FAnUz4zT7CR3+S7mTQcpQP1ct1Vm2GFybKrT9L1Q17DeOsvKvIxHWkxAIOO8taA2b0JcCrS
CVGPSRZrlsKLxQR/EV5y5seSixK6RL+V4aP0TEw400cZucUUTNVdb8Tq5GG46TJ7DR6HfVJMOgPr
/uGRfFiShZYCn3869qSK8oyjv5EEHJebZ1x1LMWHD+EKcOLW5KYTrRJ8QVG30cnunoAh9vafJEy3
ilA6SBqP8KknmojCptFx15HNC4rq6hDyLfeRQ0KbWCOSxXmr4mLYdUPZxNeVZOXF2lRwmeXuNmXS
ed9HPtcVLZxPhfruGNvfnbchhx4QU/E6hCRSVWyl6687UveNALA1sch99J2+rQx+cEFgS8n6K77U
Q1j3tKgvOjtYjP+UFVZjIQ+Ksw2x2e8r9xSWipn9Q4GpgOYYZ69IVjXbxHjapWC3A09Siz4RNCXg
5XVaW2jrMvEkQf2ADF8MdpFkgEunZjsMF+SYn+ophRrWEUv9BRcwPtXT/fbrRPsY8giN4Ixt/G9F
vqyHqGK3gsrGRPsqSt5vpNFaxUmpuzaZRP26WMXKkPCBcrFtxNK30KlXPyHXC8YCCzmsjT9sCsYk
RcIvcXk7hAUvZC4oe+7Lo/EGInCst/AffiIPBrU+/SGoF/yrl9F/KKXnMePff63Vy4Nb1sMKzr89
jgspVqEmhaX/rpM37aKt07ivCJE3bjv0+/tOGnmzPaJebVhe1FdEg+2dvx8PtQSGZM6cBhdt/bbQ
MWomG1MB9+N6f1U1cHv2HpWDSf9FDUI7JxfmcIm7BlQtFcmmU0yUuXPKnTgGz4rl9Fgl+SCe3lzX
jFlIkMfFzDcrHDLJ39Slw6JdN7Qt8pDQS7DMZpwy+zIX9Vtdz5ewQEf27Y157WJinm+Fw6YplnU/
qhpgGPWj6jk39BEPxYtvx6lmo+MRatQ8M4Av/4ETVcEZt/lnHvCM0b2tnhec96fxdIXTH0eXWgTL
itivsrchlDrL1TPvac39ipQN1HCvMie9B1xqdo4YBTi5TQ3mukVs4+LDJrm9c0GB3hxJv0L/oX83
ZfAI7QRp6WzaJcvhwliZmVYhitnqv9I8vxrNIMbhmXcYH18BudUF4yVMCm65p+cYxV47te0K6cD0
lxXKlVWUp9TuLdGW6bWM+7zticWgPzFA6zyinw5veg3ZudzVHXrzlAAnGYk2Oant9PSct0gtdulB
1UejuIuAVt6cyLQ9d96S0FSx2H4PbyZ0/jk5yh7zAv9RQsuhx/fjyWwBrumHqksgHVUarBYbF30f
0uQXCNWjEMcmEn7giaiak6BC4jsjBsPV6ESYDkBjiH70r5Dn6u77DyksUk8L3cYorPv0eNLK+eMA
D/hnGRG6omWJFL3uEZVVtP/iZ8hpJEF40mZREsUTKtp0lHPd6TRU95evIXcK0JONNuHPQLwkbPsy
lPMsN6DGkPn0XJPAbqQfaC3KoGP25Hz47Rjp9EKEuwiLDzrUGyDmt6pnkS/vNLtFc/HXwPgWeD4j
amhPsPMG+MjtVo9ynZeB++QcdPJX+GggYeHbd85NNnm6DIvWB8VIHqipl7dL51Pw9h35ck+7CBUZ
FvK54EV6glBhcElMv3sd3Hd4OQabCTGa07g4t0k7mxfj6Cds6OUIjAgJcK3lnxKbr14RafgTpci3
+zrM04hJsi2M4uVu5nFArOPD6t6/dMNxrk2JXLzxllsJy1lCrH381H7bJOjqeMKk0ZY/0op91JBr
URIIyGuS3zzSGK8BaQEs4UCxhvbWmYPHDINbW7f9dLQlbyeRpudttY4bq1QqYpHUK4B9/3Ws9/PX
sJvwdZzzyJVYR7qDVFQAx43AFjEHqdXwaa8T/mU7D2R/DL/bVUKVDzyOBwcVuZOu2ihyIBfY0LGN
0g94qkELVu1qMDwG+wTGZ0XoIQAl6BKBJF5NmQhdy7cD+Gm6f9+Kv8ZjkhBQVRnGtMN4eFsYYDZC
O0UQwzmKwmX6P2gTv8tGN0Z2K8cPTXH4ZhqRU588kpHEKMuS62r55VLAferwYkivfoRVJC66P25c
eBAAK0E1/28P5US6Znr+t8y9qmz9aMUiFCPk/pPaWdJcwErntUkVU8QpvaQATpy1LNBErThVDJye
Lac7tKxFUpc+22iyDt6b1sYULbs2ZbRyx+7ssbu9Huuwewy0lMRBATVE6e6sG92Kwwm4P5pXIHdX
JKT9GFZ4qAZ4WgnmHchsjwCtKL5l06BPrxQot2M/oM6q1GTI5xNs1e5MvcKzCDrAydggUEdOhza1
XyG0kiVmFRi9SsHIJrIKjohTutabT2GN05ZNK8ajccagS4q/aULa62iWxyUrA2aTJEh8O5yeXBci
hW3GVEqMrhGYDA5VXrnbzRmWq+85K0IFjH8QMICaBpJgBgkASR6OG8MuSO8AUeXgL6jtdmX8LWPv
nNJPQfb8pgirwvnnQ1PCmzXxzwJr85MimyPyqs0taHnoLljYUTlG5qceHkQHU74cvpjU/UwM7Rvi
fzibfMMS8x581gDm4ajcdGVNbhuB8XXbMw9c2mu/KkFaEQdRNibRVA8Lh15qStINXPfCqH2AQ+sy
1VZrQP3GDOGTSB/gq8dypvvf4ddRwbZinHCnMENbiFuvFmdAfFddntTLYMteNKAHqciM5sbhrQ6S
mcnxpU2yvGJWhXiFm29SHRrRN5JCgncIRKQpKS04gpX+vx9EHI3ZwqReGNqn1lFbthERSxo/9HPF
s3NBw6rPAOAg/2LUsqbz7cMnE9vSZgw6a+U0KTuD9IAG4zou9K54v/lVFONNasUuX5rxUGVuRM8j
UW9kv5xueHl+yXQ7Iw88GS2PxeuP1E33/H3lAxGaQW0boJhbcsJu+hN8NyfCOc279sHMx8dt8TAx
i3sdf3VjJwS+ArG5UYItglllvbaWecE9bsGHSHxv40PthgrIng0MwrFxLMfZBEDWlUgplxtwlIbW
Tv3zxVM9T3/FUyMtuNpRnr5P2BgHGXN8lKzLZAJGRmE2bQ+5gLhg/x+ZDG3RJR1UEWfbj7KNSe4y
xJXUyhqRlm2d6sQJqOEYbBeqo4xbZ0n/kqK3D+ngkcebZcH3z3A3E6Y6Gy3+60iSjmEV4jTCQpYe
txrqNmbUphyYCD9psAJmzMHjbkgVo6g3I3Xu33hsd/XumTAUS8+ZM3CIcHAyyke2AFvWR031hl4f
d9bRFxFM93/bpEOBnb3V/4vKb/GuBDuh3mA/hRhx5I/OT/sMwCzAnbs/58pzPW9ASn16+RjFJvlK
Dsa+VVBgcD8kq+z+QS1cJQpkUrgZ9uh8Lpgr5DhCYUzJdheVAS5BpbXnzePiRUhN9ulqMiuK8tut
yAK28JqW9tMSVXrmPA4o1W0twRqi1+sA+rSe1eojKT44unQSts31hngdtMlWGKmfQ3ihHp1UWt5l
unHDiDo+UpGSiivUA/N7ztFyADfUNKSMAEX3QL2o/l/qqp6S7O9O+gVbyvCwKW4pnkfEaTWTIeda
iYbnJjapUKsGtStaOdPy1ZIPM9DyMAM70NWmy7TgEow4roda3L4QvFw+0fcmNHIyDJya+WENe1UR
S1oSLZqsFQJGhKQ6vQqr3Uw0+0HUgPYRn4QI+lUmknqzup3MfGf0afIjcAp9Y0vnVwLBMRSJOOCs
G4TnpulbT7WlWAYf71hQyY/pwLKfDCDYYD38CuPubCvYwR2G0esVAuaZc7DFNNe5XGeKi9P85AQj
LOHgIjRok2tqOY+zOJmI/ecYug4Ku8LzOjCxxw5kYcf4GVV0WhE0CNZQDA0/uV+FhCJtSK2gKG+y
us8btOtmsrBoG3IjbLKKDQfBaxySPg2Yj0y5+d8VhEHeNQ6e17iEN3w3ko0PljYWEtYDDK3T/laC
nehgcaj0zLFNiaL93LnYKbWgYyw37ld5MZ5vROPtpyobyF//lc90D1Tf6xoj+OyTMP53MlXGq00i
PWrY/ue4hLG5veIJtlyKg0bpfh0K+u9xi/ZFcM9nfkzDRLPPlDOE1/HQS4NRzbDZldpr+2qVDRKG
Z2M/LTPW3Rt7FOiaGdkahsBg4ZYuDzVROPHCYwBT0Ro/qW2xAxlt3qFyjwn/Pri1ELHG2cTxFTxl
c9MsNFM4bwaDOIsvkJ8oiB/hJzg41gFmu4SXmg1D0gWevi9/VNz/FTKz4C070p/WUjO+Iwc6fl67
wjSlZwk8yuT6dwAZoJkyJkMeX/uysi+m+/0sXmDyms5ftXxRxRCUuxkEFmHWIcxdwOeKCoowyj4i
eUg7MgB7HB7P7bO+tjlof1ufrjQE995tkxalzY3o5iR9CfVeERi7CMvaNxXleswJ9kIJugwAGrDs
blaF4Y0H+b0mc0ElEkkhjKuhgvfC/lYwC57OBWqoVfU9VFPBQ7d6f2SZ0Kp+ta5u9xvrQv68OJ88
shzNhx+I4bQ3L1Hyg8DBvJWRDCBXzz25eoWmjmm3HAIh0nc7WtTgyvAKQq1b5UA0krcDn6FN+i3K
WaKwaPK52YQr8+MOcB0Z1yqa/JxZZO8qHSMmGJujLXQtlOIQBQ6TcQD0T+GkCMoE+TiClxbob4yP
iUO7FXclLgCSQoJVt4VYWi2x2uig2YKSN3YrnIezVHQGGtRYl13zM2J/tlW5NSiUbB+9j4HoDLC/
ZY5BD5DxkODoz44hKVxvW8G3Vbcgzri6EzfUC7IHMuybphW4IZwfJrg8OnSbm/UdP7cwxDE0GUiR
rNmZe9+c3P+NVocAnPgrtiPnvJ29HH4/J244ngDppdvZJsipXvu4T1tty++uATKpsoc6guvl5OrU
P/m07LBWrkrIs6+duv3reyl0RPgX8ej9N21EXuHK3aJUL9zF7/kkbrhs6s+OV6JIYeSZG9AleC4p
ZXXkyUZvr9RCoyqmWQtUzUdGelF0ebEmhbKYO0KcQvV44Evx/d5TmSsQ2apJdUHS/jwWk1d1PhWg
GhCj9jwLFSGNEj7G6h1xHxCr4CKogzLyps86kCaO8jB/IFmJ25hiKoemDe6I1InP2WVXRm0XVq7v
BKlRJGHdTAln/tViULXcVkYvBBIQDce3hE2fXTlSIlkj1Ef0HgywxVHM8xABn5KMMR36zYnY99nI
pu2kvmdXn2RUsoIO/qwTyyWPxA5u8RSHQxAlIu5aRXcYNqsTnwnFS5yu3TjcXnTlEY2oCLOyKWID
8x6MBg+oQyGiDJcANqm+m9adrWfCzOyzhoNJ3GYKxs39hRQfN10b7oj1f8NuutXJN5LQMxfsCxCY
cNpppWSRDWLoq8ZkQyFQC43O2z0Lgid8QZVTxglGtix/6mno8GrECf0kH2xGvBQ8yQXSHMILTbRk
5CtrNUQzdUlDbGlwzWuwKwnyuiPMIjQvTMqGjGyhJxROE5y19c7+aC5kCVUxhETnBcEjrjLYEGDo
HaMFBkDpCfwpvczoTHHz6ajGpwJod2le81ViBPJPPMrN+wJD1gmeq0gYsoxaM4rnPl8D+BcYI7HE
1oH6dKCk02A9sHUUlZ3cuNWW5ueK+Svvkwy8S0N/C5L7aW5eSc9a+qLNFBkNGN09LV9hbEgtBy/T
/6BLJ5r/8KKBkZRiLcAyjiGwECS6oOHupy3pV/dRjQ7xvK/8E6WUuNDXSB3mFnm+czXHA9GOMe14
UfEoSh8iuHugZ3oaNy0cr2Gv41LW8MEL1GGHZF7Py3pY/3GUhO54SOv5QifFCsisXRP47ayTTW9K
q13r80GZzEnpMvDaHdH6MDKqfNUTd0fu9UQ2qOBNHUE6ZRdFgPawSsSetQmi+kfM8z/akg700m4f
qFFD1Omutrrzop+Eoqq/EW/Bta/UCgyAIIWjYbakzQgoc958hrELq1zKNLzYvFXKKkshsAmpitkW
7vsD92FhNMGLCXJ0ckqsHGilFYENsNx72I6Kobsn+Jcws1587DLHXDKfcM8uea1BF7zrMoZ9augw
yGqLZK0EGppLhJAfeXaxSHyPkJ93UX25wOuz3Ae/ab2xFvLRGS9H4gpr1IumxAVcEiWAbWvwFIKw
vxMsLD+rBWLKU0eh36c0Ie5dWAFWRI1G3B+GPqhVLXpJJOMbZmJgkkksB330xcMcUau4WA0DF+3u
B0/LI5JKKBVviA3m7+c91yNgiFfg9nI28C8YlpJlwyomc8Nu/MxCusAQEqPCWztX8C/bVW0Mff77
kSwd3m5o52/8Sdq1iYUxST0UW10+eX4jyK6cnYYt3ncny51ZBXaHRf+hIfRgiIPI2rNnahMF639e
UcHa9Gk/qrZIwpBZ76LV24r8z+SAQAH36I+Ss9HxKvZcZGGpPvBOUoyFFZgDICarr5cTiyRtGiui
MCOMg0P0v9THI2vbb31fQ2BertFJh/lXGhVmwUWAWwcGbNzCGV0QIeFTxCc4mbD4fWKhRktf7XmQ
7YHS/7loqRnpmgsedE1w24GBAFDIyb5YXQ/jAEC4XCpi/tuBHX/GndVyAejXpJJFa4yTpZXfvG/j
4H3RzTiX1iFuJKrWBnrttdRIyzkMFW6fdJE/I5QScSTph/po96Ngh71f2mz0KyXtUxX7PkGoXe07
t6HokSqfvw8annxiPe+gBSxwLkkB+JQyVXmrBfZvWMAm35T0JMDDewKa397L5/7OW7zCPT1Zo3ok
gJ5WV07zpofxgZzSsbOiTDHsNUBnMgZ2XZz21wBippe8xN9Aui9qVwol0ZgUmmzHYcne6poNWQcv
UNxkBt4MotJl9whvYGpZtOVFGhZK3oQijd7rBrRth22DMKDQvwkNyO57KPd7RYThnjp9umPXkKCx
KHwpeAj6WRvobAstFv1Yf5kG1/QM8HoPkccn0vjOVgfbDzqcUspKHRcbJDxC8RHnYQLAXmWfUuly
aMizvDUpZTAh8yPskXxCmWARrWK661tHIuHbcLTWDAA5ej0+OFfDkknEb4g61ZXUcPO6RCkpE9V5
+2kvCPteAGgKXEhIzaC/id0tnajbomWQ53AZqcD+cqlBTnvydESCb+WOuY9iyUGxH4qpQHff263l
/CkYfyskMGjHRlIRznaZ0qWgCfu8JKnK7BVvEld2VS3T1pAEQI0+OTRXZrtmd3s8JmOzXnj9auVb
17K7MwBMig5SRByZgsTOQFzYUwsG1v2WdM0xbi0aBKne5Odfbtl0Q3x68MtXpoUsGqK2/gr6h8qe
gIoQ0apbBNnU6ThV0AlTBf0dXSrVvoA++rASsl0lal1cS6mkWqAqOoBkdPITsQdHxHUs1ZgaFvhW
kM9ZByT3Csu56d7+1Y/Xa9Wt18DzwcdAOaQ/v/4TroNIDTilIPQTFx3xo2jsi29xLin4kdOonNLu
XujAeWsBYLQIPpzeveQRQLWssWe0zJzOhPrmWFkK3E0g2qQnOP8VSRnvUfEselaos3g5tDYlub3U
oRvwsGFBYZ1G68O+ibAU9Eg6E1lNvoviPIo2wWnQg30tuI4XbZNNNaZiieWY5McW1VmkBOQ5oVkN
3PbFTlOM/iMYnNyBEncjgV9Zk9mMQZpo4YTGrYYz3K/BSWpm2y00JOhG0zczblYecJqOjpSnfk3R
huEklwJZ6rDc/+mpA5Nj2Xh4cVCTUeWX3Nd1lZbs/gZaQbAxn1PDXhAs4JePYlWxM9RJ190HwdXI
YxWL1SiOrafKGM0ShvJI6KFa/9NpUEdrEinqkDACZ4cOf/wub4bwerj8RvymlMdA7XvEYGW5H0/o
P1oTWgsotel4TxmEdiIN3NCzaK4up8/UoV/jDt1PT+rpssGUYS3hl1x2hDRuUVQnA7wRelmS8SJA
CCOavlIw/2ZXVuVpEw4P3tkorziiOh103Bfk05zpdOzGYEVEi4SI3SXw+foGiPRM9PUvcFYl82gS
ZJ/ZZySkxJayelzP9wbmeXlvTX0+SfTlpmqfCaoisq2kT5WcoIRQg0iGGx9uT3RJtsdIz8VetuCO
ZUfT3PlpN9otPDoBPABykAeD0EgH4t/ksFLOmCpX5dOHJlLZJLWsfMiAHE2NoRY0HfsB4sq4yu+9
WwDGGY0H9HSJ2+Qn2sVEtgDKmyAkaouUJOAh9WolM1/uC8+DPy1GTkEO+RFvT3HLSFaFTGJnl8O8
+FFCAiv1DNtMCsOxOOMzryhqnro538oA+ggBrQM8hcT/BebGNibOFZ870ruLVJzypxYX1bobIpVN
quRD3NtZlQ/7zD6/JfDc41+b3IPCSyDX5cDM7DVwSDdDpWcUS4d8B9fxRjRc29UUMI/Xr5XcwSQj
k2Y1U8UIUwnMJGsREmP/Ls+HemeYnUFyy9BH8stzbaaRndRl76CD3iwz6Q6BQAhnmgd8eWBvpiy/
VWvpJjS0nWOKUalOBfzOCzgh5FidCwNcg5hgST8Re2nY6LAB/jK/AfOIL7cEKGVAsim+iG2hJ2v2
8K5C/ly0jV15oFRIFWT0tK6nQMymL+wToY+OWJv39m+38mbDYN5C/7jkhJl8Je94zUF7fWWxzOHv
66ztjatg0U/5Nt44UkeGkFYyc5y+HEd+vCecxeft/jthbq2L3n1aW9opEPLyP180ornghKGA1tb+
YN4gNECDACepMd78kSQOCwcO8rtuSWDV6lPBshIGxWTpYHx2Q6PSVi+5nkJMejTgegxcQ66WaHz5
CHZljIIkV7Ggm99GptWvJSzr2mO4y9VJHD4CnFEk//uqVX5ObM9SmETukBLmz0F6e9Oe0ZvVKH2M
4zMRypk460NqJAX2ndXccMLKyOzNkGllUG8wj4AXpbWP3lBcd3AgCgWW8ab96qRIf4TfqdrNkRhN
JV1gtpmJ8H79ovkokbQR94L9f5OrBGQ8nQHIkAL8rOL0KMoUwlkjYJwn0WMy+tM6Qx1l29tGmQe6
mX0ggS8DqDs3hnM3hBE8wJpRGcrMnwmuzDNXMUyWKhq/KU9iEg9fPbHWIyufwcJFsmOlG8W6W2Qh
clDHrQkeZK56bviMXEpwzdvc4FFSn4lCC7erVd+YNSGgGL1f21xY72qnS9YERfv48hGz29gFIc7+
SioCA4fiXWpz6DHfP6PqtFVNC+sR+dQl+G97WrK79De8Yb0P41ATS/PxwFkpDKjCdSRAV6wrr6pc
/8U90deCLO+6f72czULmrFjXoz+LgGyTgz8HidHTYxSjcaxW3pkvj4knrs40AuRPFRFXNF++CAlG
+k9OYx7kKy/Z+pMKI/iF5fmABq6MVxQG88c+AXCPQispuCcfeUVj/rE1kQs1pHEgLVye1NWI9li4
M3DH/0frZ5BaS2SUxyjvNLZNe0R7k+bANGhQ1paIc/F+QIatxlpX7wy13VU0ihBkLFkZ9eEMxGqA
0KZ9fVOLgDelnZ9y2PoLgaBExkGucHd7VVpVl5anjQfimUxFECwGChc6INKg10bWaOTvjtkVKbgd
ITmKLVcxEH/QNjrOzftQqcg8h+xJT2MKsb+rEDtRMXZoc7H5qX3aHCNDZGI74AqDk1WuyeE0x4Uc
H2lCXUz+8LME4pFQx2qIKjqui03RfGI2LE7MWqT7B8KqYCygWJJ7NXIASqhZ5ePWiMArXG5U+82P
QDAxEz+SxVYhXCtPZiydjNnhehjEozHOltQOo9vw+NyAxUJw4v0zMN3Bg3K67Epo5+xWZHrNUrNd
VzAkZauneIkSjCUfv4pof1ZCQG+QufSoQ4nBDX5HvOqYaTL9zw/FdHx4dI96PnOpcn+ooYxHvCWg
vvNjXFipf4e5b33eADmTXbLd5JT/YmD/kWoBQKXXCgMX5peGronhD7g2/g9DZdtmm2K1DuXqfrJA
gu0S5kT0IF48oeqjqvJP6+KQKWZp6NXPKWGg6HA161GA/e5LLZwnkEzb5CbyglJukgvbpBSdNFAy
9LP9x/CcnopM98d2ZDb3Eq+1PQA1aYbVUsodk8Lmh6No3RxBCILFDsgFxEgDiFbXOWvvfy3Rr9WY
N+GdYznlJQmVZSuCl/D8XyZWUvzQWxcpis9VGt5p+ApZx3Pfb3wBD/Ynxk/mRTMH+uEuS0LpoNVz
sCM3VHzJRMVew43vMKZKsvKom/TpP4oCvLKhxY2NxY/Haq5pDtDOocnSEUbTfA85xfYg9Im0vL6C
xFlJQ70bxe+UAztc4iF8OUnceZTuDUFpCtPlJDf9u1I3I0FYc84KrP4nHvfrrFkeXi4XUpEJ2wDc
IcpE1hI4+Bm3848whBjpQfcoyvTBsC7ZJmn8vhPT5q2Ut9Lfgknm5N+vYNxcstENoUCSzg4gZ50D
DOZ4lnxOZ53okE0AIoYObl5tT6XfFJNRDpj9ZGIkK3X8/xozLti4d4PTep/FsTMRBr1AGduB7c1L
+asKCk1xc3D/r4BgSO2lMzux4+zaP28kVFaueB5hrPSsPzRNDS26LdiNec4CIfKQGOqoi1usgCwM
kfJ1ibM9XFAzGsZ//eAxsYn9puW5LL5HxnN+sg8Ou8ECutMgv3rKz6KGCqDNbQWu9B6OR5jCvcSj
j3t7jATE1rN+Mohv1ydcW60Ft71Bd9YV2oRi50oWGvjsOYYKhygZbJUMxKXM1S/136Tuyw1hHfNX
J9HlC50nDhJw1782mQFW6Z0d90M9ctGgZsvErKnBTFn3o1aP7BoVtdYNsMrivl+2JcO8q8vSAhZK
2MMj5QpnB7KAGLpRCfn+JVH5IG6HaF0e5xRRFe9HNtirqzkyWteIGXXguoUPSfcv9c4A+7ON00tw
9MXArUzFL3JuZgjBjLGwxhuzuehSFLykZT0BELF/jZQ3FXH1CmK+I52f2oC9S1DtuvVahx6M+/Ma
Cz2NKbQSouNXN/U2oBPWv7UaDHX5KLR5SfYI4rnv2E1oIhfkRCjSokXrHitOuCJCS8yDs1JBjBqT
7d4UmM275lCzDVaeelzJAOb46/WcBmdXzHzbJRREphHZi6pTGaXuuvE2kcdocnkZGWOio9qFtYpA
Brgv/4TbCGhhFwb3YCRcQB8eDJR0/Imki4NPd8S0+gnYHHiYcqH5heyg9Rgf8VJm6hs6adjdIES8
YLHEYu0exmvdJZF7iFmPFYR2WcndxvSiyfgV3GjVvY/6+yhAvL16JVbpU31F59l5kyJ8jxqxakHF
t80qdlobqL/xM2KbwTuaj9Gajil8zb+Gog+mUb2WGQHwqWIuGok/fQ+4ElVma73wlidQ6aslCeIU
u+Zuq0iQKnq1m3uuwxSrce+Ta8HPIyGOgT8n9fXF7NAxbPMHxaZYAJYb/3QBQF9ZfiHLr78XGPpH
bM2nYc01V4PT0hCpH8nAPvribqz2WHnlEIVmUKASaupAPSvwt2bMaUpzgQ5Fh8rdmNPEBpGRNO+t
F7SUXzyIqUxS4nRI7UD7A4BV/a+8k6NPeJr+e8SO/NOgmGEk2r+I0vG72qi2CwNS2zzk1VlnwIQ+
lfl8ETUur1Nmyc3hiXrSNMcvOvs7JjmkinNW0phB1CTec3GpMONlqc58ED6w4MLObQLhTHfjnf4R
tP2V66zHwHgT3LX+XioXdAYVM85vCHug2B7GRRjUnFOcULWCGwz+9n5J3vpqBgt3TfUBGV8VAupy
eAaCmbQbEb/nLaUDUCYqeolm2UYvld6tqAyjnpN+pI1qT4qW3Nzg3b6RTgTD8VQ1us+VXfiY9B+b
uUGkgjQ6ejsoFtrv6QOltc8x433FggaNOoceRr5IHvewAyd+HI4Dk4w3jO93d/76RSnDmt4nfufO
wqHmjGIeW3XFzgNRO+gZ5PeCnncegZ0+3fbjnly41oYwMpZlTgGxL5xFP6ngoPngkd/We2sBnIMM
fp9lXloMy7okxrbdwXXJRJJmdA5kmUQtyKTiKSWnKeXqPN5IAgc23ebJ0L12kS8shijeBSWjLAPU
ucmtPrj2cRqgGAwzxXHQvybOWF5eTI//1vd57VEqHvaRH3eYUhdybSJ8QHbVXdT+J49JiIhGXJVL
Qx/VOXnLOEk0p1ZHKbGE6Ii+jx9JJ+S4+5IbSDpLxOG8Y9zSkWCC+3gDawWn/KRCVqklHBfR7sCj
VEJbQLwdOZGA38LFuhin1KeB6Drg7IRBfV4eqKzuN8UGbjXHWRoxNE22Cetaot41wiVYqbzXBfQ+
6Dhq+6EccuSpDCWNUmeg7PeI8n86XKhlSyjB3smpmx4IiC1lZjyVjKd3CPYacXip4RobmlbYx9vF
lzmGtytPFnJ8cMwenqnmawbwMl2Nqx+Hbnvy7G21yZr7aIHmmI/IXKRRzOquhHY+zMcGEyK5t2MC
eqJ7xIv9tp3Y9rqkNaCyX4wN0STJ1o1+ZOyKA5DV5akeQkzS1u7ME0n928LIVxZhKr39O7HM16Vk
wFHieJ9qCi/Jba0DLCXkkf/KpYGnok87VQnV1g4+ow9kk9ckroguyN59N7EZlfmzIVOUXKttcejS
OCQyusdb0anmfH40IjHLMw8lsJFrMgs85qA8jz8q8zmQpmVqG9rJG8czNf5THX81JA02JkLv3vzm
A1JvSbiGPIiNl9WyMQtxsGp9Novz4P8+Dibz1zgDN5I+9hxQOljK+npXYvtXimVdFyeWTUCIFvSl
sirepLzJVvKRESJOXhv+Xs2Ke4GPkpkXw5Uif8URIc70JrcDimB44CPsA52dInixMBvkCrWyBiXI
wq+deS9DRaMWzMzVP/MwbZT8NOslfuQ65PwE7MKfTvJ1epk6r03Nso82YOo+iLuhxPAmGBO/y6WT
0Bl7omK4poHJxwX7d6XWH8UQbHNPMA0Ro1arxDhSQ/7y52maHwpuz3sljf/St1/00uJn37PbPlCU
aCGt69JV9O5ORfXqNc3tWpQ9PYYmtvziYm0ItHLcv65wFzxocQo/9dOer17nAWP/lm0RwXMD76x4
wsGKS/JLEEV3WbayDnGZ8cS7LlRi7wUvL1qpn8HIlIrHWUC457bK23CQAqwDiCNgkH/AlSJJBPWp
dxD+CmAqnwJLjTzHhVybKi/gJcUIEuos7VMrhEUhIdOG+Mi1PwX2meeSNnl7BEd+oPrH6CiTaQjD
+CldgOowbLVe6logqK8Ty8c2W40shUZueTXlQwUuAzsTq7ZiCwY2G+9q7by4b+KrGofoLPDd0T/a
Jpng0nKjbXXPNluoisMj5MOHDwpL0W9pab4SxjA2TikATGrNsYE/mXMhVlUT7Kh8FS8LgtVa35+v
2tEXUmYUs2uVwkin2pukBVWRhIpVWhmI6R2Ab+YqUp48udw0Y+K6Q1W9/40QNh+HrUxhHZ3uZATf
MMlVp8KX8HA50HsE7X+ITO27hzYuPan5QDZKsdPn5XK7B3iy1j/lIb0tVCL70Gl+0NXnGjW9CGKi
wnc27bw+BYMhw1wnxJjCeYwrdtbT6iEUKnU4wuyJJyq+PLxu5C7VDlyQD6gF18ZXdaDy/UDqF0IG
7S7KTKlXvkRpNWoRnPXU9xjLuVTOsAyh0ox8GdKtqwEP9Y36r0RiXYyzjav4VCkCPDznixpZJf+W
M8GnT0ZcRrkOc+Y2GLHSnzorhdDJtkeAhWKIkAQeO7IAYPYgVwVplUrJkd4H2eNJn2nflFjhrPDI
hPJEjKLZxM9LjN352X2BT4Uh285HYxxQkXNCgUbk+eY7ATfovdHjbWh9SJ+DGH26M7w0CuQXdSAl
dZYrlMigvAp/nQvAoMqQ2iu7/+tSFcvDOblVCJnsvPLi0HoQf/OVBFp1+dthxT8cj0OCNhhrqDEB
ArzNoJRYnwtIqnJtjBbUVF9sZISH/SownXdeK3Tz1kRDoxAw/MRp5JC8jsmaR6XDqndjI5EgIh4S
Lw6L9BiqenqLemdAc9H2zYfvY9bO8ZabbsfijNJ18fkAp15NfrGlfUtAnQlK0zPzPkMaaCYND5EY
LjNeUqJ8ZoISWT/Re+rBMYPNAevx6SD1g0aomMm6XBgwHRix9LEF4gPETef52+PlNHqM1OYLy7mw
6o12XX1LdcURcz4F4QeB9UKwPPSR1W8ma5e2EAb/ftod6ybahP+WHE+3ZUsbNNF9lYRcIv3crJCK
6DLCKeUnIBPzZHWxLFB2wkMhrC4lsfM9PL/HMvaf7mTaomuTnbi7LFGMil3Y21zgAh4qo8JrXGfv
7+mhOPzd6xQ6QZfP/wgjJ8D9+e53B5Vn+iS7ey0ydbqgEAFjGtTjb+UMJI9KVWU/txSnXZ6Rkc0m
W5ncxRq9iLhDGGjriz09JWBnbLVXqCmUjUcYzlkO6dMP8iFwFuKLhPv/7dUvxOgWWAPkSGNtcZtc
rIK4eKIZvh4ud7Nas+hJ/U++MeVaD3KtwEhRlZ0EFK/FwFA0rDVOy5vsYmxjAk9N0g/QOyHCFDbH
OH1KcfywKA8pee+NElYh2HX/vPUGDEF8Bllk5qNyNkd9h+Ggl01eZp57WvGqeDDbeAfzC1gllrnb
KCUMYPfxEmhQOpC+SuZ+UYEp2cfna8YAm0uaMDDva79cTRt6XUnKXEFQCuFkX2Mw/MVd777VsuSE
9MfL3qF5kGRMBDTb+e69G94MMWaFNM7e0zISFqsu1BcNNH7kMqKW8F+ghBZT28P+5GgYVAJvXJzD
basjkTeJP645UHdgFOmEdc2iQz1p6C0W/Xi3Ucudwaybc8rGo28q5NeK0E8L1gVkJq5WjjO96CbV
6S4woaBQr6rL7BUTj/hNQtAu7o1rXc9rsMVgPGBFGpNRduThIevIa1AHhGM3CfsydN+1VjgL+hWI
nT1HtVHs7C09aScHmDxidTgEQibZegkZUDqnZYjYc0lbry9YorgxMInSqSfeF/1UO0Im9KGcsEvs
ZKKiL/TvNRAvzKnpLVvg/6yv3aBrlS741VMYUI2Rxp54/rTKTB8KVt/7tKczX3b8YdiHujznFpii
YZyHWco9aAH8RkyEwQ9tvvQLHUOS7QjI2wwFILtvxTh62pX7j3yK2PJQrfPso7sWMfnT2R+V34es
P2hqTteQI3v9wm+VXkujvapnYDEhXEJ7s/VanFz7xt2BWmdHO0iQE8agnsqTvCDvbGO1mWVnJ4GX
pSG3/RNO33QhwaGadnVkpL5SZ6AdunBOmvAGWrON7N2rtL8aaYJ7aUr9IeTb/zdJwFfnwk/I7L2z
pNDN7n9NevbLhjH6DxyQrkLw+G5Wr4A0ejG/v/Fz8fQiKVH1N/7Ue0xkEVpW3zV+Kek1uq2oU4gV
0cw6QSAyOPH5csBoggDAD7mJr101W3mr9TlYnNZO5A2zmw3khM9Q6TgZkWCGhpfpyGDbZR8vpSKW
BGOwP1phi7znyWNYhxNlCZTeVoQsFs9P1O4tOAallNdFM878g8Ha/bGOi8u9W3IZt/IUhN4c2J72
7ZMXhSTOcrNeik/nW+A3TbpMDJjpzY3Mke0jMwo8t1r6zBRfjh8dJLQucK8KXmcA6yJ1retIfX8B
r/yIXxmFJLAG/JHS0LNGbUY1lE4LllfSFJYOoL5yDcrvBsF69YZPHcvvmwuhh2MZ371bliOZrvkW
DsUxlcHsEVCRRYZZxUYBeMhx+juajQWaEEveg4zg5ZFEkLpAdND/2CJMAIBEyCWPzPcljzc0yA8V
XrW/xCN4qVVZP+zWvLBkOP8qpKiNyesvurEjfo4//gasNAvEJp5OZj+3MpTLJmN9RKXcPWZZ50eM
sNsU5Tk5YHQNat39eKzTLq4+mZq0lcaEPetbojI++WkcIko1VHwM/B+mNalCXtG2xxvHm496D63m
Zj/Y9qivGiHPdER/QVxSfhluC+8da8z8OsF85VZAgpaty09o05Z4tXorFdu1M7p4HK+22NN1jY4b
wSXcRZB0zoIBwrIQphyxaMTbirM1n2gbJZdjZ+xKVKgoaYz/Qy0Heq1Bo4tBRAw/+8RA/cwZCj4o
WLSIS4IjcLnYY5Yfofe8kLFtbLSXhkR1fjGyRyZFtKdlJoGW//TmoeyWl8lVVaAvingcGz4/9h/o
MOzpfel13AD6akCDlLQUg/uazSdDXul/zot+16FY0Dsapb1LRpnt9NI7xr3XLUerSkgd/TPdxhqe
TScGGLjQqRl7AcHpd2KSvk+yvSwPfKlVom1OiD/o2m3nFzJExqQZ959Iz8+AfGm376AfJsKUqqTy
h0kgxH6isKv4bpHwZF+M9eG3sL0Sv4FDJ2ZlqJ0DmeVhI5KDZG+SavEHCb4RSE5RCHpC/hwlZR8h
SGt7WHCiRpFizqWJTCt8VwHZib8E14Ce7CZCY5PRESCZ3aXqK2acjrS1RIsyeiezi5d8mUvzC70P
qzj8Ff3vhgTJEQ1snaree0xh4v7H4izS0f2DHZ1IBbLhXSkCPSb0PROSCHE5SPVkiuGN1HsuGHxf
DRNiX85lLu5Txnqrw89GAq84f2CypwEVHSS7W7o8orZ/VU0sFosNtpCyZfB2Im9GtIVbxlsOHX0y
JG/0n7m+Gd/iGRlaHQ6wSPJusm3D10PLplGjS+KI4LiaHEHwXnxkOWld6NyK5Zm4NvrQEronFuJV
4vPYzbmaxCNPgO5dWU5hVthtyXIxwzpTDsZ0vd/HwooOSRrsBs6Inuo/2QQkF70W1KSB9JtC1yWW
YwI28aJ0pb67OB2Y8VS5UniFw5KXDbl1y1oa9mMLnFuyL8o6nf4zOTOXo8KlIyvRCS//pnp0kOt1
n7lHKfhzwg0K1iiY646e1JT16NJNQV3nqvBzuXn/hIpNVeD1yNDbx7FopJTlE1u9skJD4TuOFUD9
Ur5zOKVaKaAL4g3r6bjyhrEWGGUeoN6CxvG9qpMBHO25//1ZlO/77LPm1UVoBXGDXKgwwM7SIDO3
x/z/8xr1Tzr6CfWCCn0RzAwS7Th/3JX/989hm3Ho++C5ma50neo2XPPZ3hfcZgRoB132jeN04r/q
RSANlOigYyum5wQjuwGLeIy8BQ8ogS6RGNpjG96ZCTJFVOB8TzIs+e6hAFRue5vSBxysd8sYsq/N
Y8in3yr/MswNo+4rCzHd8mYHTdd+k5XMOG04hmuTdiw1ChuiT5jIgrIQF/ZpWDmrvFVZlccRJPN0
4P81Rh3WlmO/Ikj9M5AtPGVvOmAAtX1V2Lv24IVq1PKAPqoZvOAiFu7RNzk/fJyr6TD+/sSyMDtv
wx5cD3jWZvb33YRAJuNLwBBBzsAsi6aG1SxdmgiM0dFthT0yjFVCafAiLHLH0YBi5WxWcxTg7v+O
HoI3pcW4XJnOSGmy3ss9A1DbkfXfB+rrpu/PtT4DOWx/ahhuK5uefjJitOdvoRaFML5jOQxT4ULc
Phro7xe47GpPYsPykEOtEt+b5a+oJdSjjwgIvIAIiKP1lX259QPYl7xlYyG0R+ceR5T6v9uPYbra
zXytcLPN1Repxyrj9IMwtcibdGg/pim0Zu44BIRewsdZjIGz1lR6QNGDrotbCdGRcUcAfmy+DTac
n60JEWxj9NyQrBz0+OO2a/dRQPTRbHiJtypkWhzdL/RhWFT58NFc3W14BVyps/G+w20lXESMRsKf
tOZbNRMSaYWipYnhCk8ydMMv9y3SXYtLNls+NN+exq0rg9+S23A4lFCsG23I+nQXcKVkFd1ZQDsV
XlseJpimN2YGak+qYlhwHFELMwnM5CnnQqxYODPSHyBh8b1dOpj9ImlAlmnHQj3vgO591s3G1MuL
p/gZuPEwB5hS5+RhHlkvO87M40fhdDUXf0Xj1+2znGhUlON7/k1Hio/myq9NiL655AuA8NrkRfjh
rOns1VrPGRMPE8hQc7OpdG0skL0MbxwHitLN9v/Lptr1Xhys2LD+FDN7FwKeHvLJ7LBxiYRZiO+U
6fnfVH5kzkNDYx7NE/Sw811GJZdWYyUWXC3IioBvjoU4oqIAxbVOoULjxo/pH6P6hFZeNkwHZ9Rz
cQ0aP9atUwq46I3t8ut0Dgj/WiFitXsWa2sxKJVOHkm1mdTSDfSAFHXtySnFGcnwj/FphcveTpnn
ibRtpSk5E7AOZ9rYt03Xiav1xDrggEtVLZqiehGuRqXd9gs6lPBfzxq897/302yZ+/jhDSw2cVmQ
qXmJTfrCChxllcKpSgTmcv/0KS3O06Z7cK3THdXeMJ/f++kl2aVdqFODy/vaTfmuWthFSVwyZnSs
+vH9m8qycjoHZGLnUC6HElriepoHPt/sUWRVCipU6MUCEu8sv37nG5jBHP+stxoTQ0cxtQ2zKuA3
Mo4clKCVjveFYRUMbtsadvgiuvB/oB6SOzBUi/nioJRlrx6a0q0T9w5tMS+N+fDSV8yW1qKg6l/Z
BQGX4ukV5oidEYnfcxNi1XoBjtfA+WDR95XIgz9bj39AWW6Ir47okfZ8n99+fFLcxZKVwpGw5MwO
asCHyuY+tc2e9shiHM7fxar7xleJyC64A2Lv2zOqcv2eyvRaTvtjHOs0i42VC66681t4zxYa5M5W
PPGJbupsLlSQA58YbBvi2d0O2lr4H9QZEJoA6S7GxTpYahslZlukbs2MPMy0OzfDmwSYZ3cqeweV
HG5PtE2JZziUJRP4SEJ1ZJmRdH61SaFgbBdudJak2Pn6QiQKiE9RrtJ8mvfJF+sV+/8a0T7MYz+s
gP28NTovgorySk5xCIQbn0a/5GFNwgPn2JU3iCjfp48KIHw5MBfHtyjZgJkd7ss0N0rflH+IoC8a
dnaKIL9UQYyCyinFbV94Qe+yAdtwbMjiXLLq8d6mV/e16VQHvR0ByPgNyyFFkVuMykMLOFa4mLrF
1ACoAyU0B+SRJCr2Kj4pncJxkLCiaS6vOIAZziBEtuu/zRLo7cozlmF050M/gYcHnp8EdtD/nXuk
PPLgWLwFCN1g/JiGzJR0i8AJlhyVhsOvF0UMzubBKACeSRASSirZ06VGwbHPquR2las97hQ8bTlP
vsvrAFtSAnoHcfyUlFrpdeRvPpRB6NYB0/rrTXM9tqCCDWE/YGG9rRAU6zk1vLdhz0XVnkxM4Q9C
EUm5GXbiquYRhOw0BCf6APgmcYhL19n1g1XaP3sDU3gXMYKAgswk/4n9jHbryq3pjjZqx46odFO0
mbVQF4VufawcSAD2foKPJBdCDmx5bKacM7Q07hfWEmRxPbTwq8VDEpVd9IXEXtDai/gPWV9KJ4LS
ApCQMXJjXCjcM8p1WpS833vVzT3ko/mMt9/WX9rtC0AjUm+6uPsx2ku7rfnOAT2NoJ9lpW/8iJRm
oFwX5AknEI9jnmKoh8Qj1NYLLiTU6xn9IrMxIUvyG4AUb1WtIRTfhir+ACyd+YWYerGaF0DiqMgK
EM+0DTudzT7AIDNaE4l+EV/9mFNKWhf3YgV6WQWUDoHDxUxD3uAMrRb2soD4soNIC61urQPVrcoY
/bEs+0pqgUis/miL6/r0k3S/RYD/YTC2SXNcmYpsdNBuI9yormz7/tkciQ9wuoeGjy7XWSN1cx/Z
JoKDxHFnGrD6sb+vOqVcBWurzs0zAW/2e+YhxWxoyRntp4ZeDMu1nIcfboBalaQke61R1Eeid8Pe
LpfctnzvdVperp/325fkhjy4aXNgYW9xwNNpj4iv3uclDU+fgZOKeAJm/iOVS7e++U0jvDscXbQ/
AfBNoMpNzTf1WKjPFfm7fmf48q+m2PVelAtTk9VoV5B9WE9/o7rhdrjcxRKC6DzjuQQa0zeo3X6Q
/0ODFDKms7y6J6A4fBi6uHs+GM0F2zDITVwB/wPiU2hYS/6Ddyq9sSVPv0Ei28S52lG1Yi8W3uan
8stxZafSsbpO5PmiuHXY8qsl5+nrD1nSCelWiHdTBIK+beSUbsh4K0MdvTkhEqhDKZZZBri2bIH1
CoxpM7W/0v81CopTx3kBswxkWAjWqs9tbxgGq+qc/2W+Dtfh93gjspwCwZ1ekZ4wNnvdVpc9apXq
UT+aoFN3FnZ37jnRxXmVPM7j5ismK9xwMdFDEiL/fI5nDVtGOEVnBEb/OFX/Q8/q1zxL6YYAfqYT
8sRaFvVTepOjPXSGNwRbndeJg0ddjDAeW1dC2VGC3FteMwA4GZ5sqQUxLfpYCMU5ct5sVghvsJJH
RIPd+3jTEB/YCLh+pWKjtXQy9CwITHykXe5KJbHou1ZIeo1hNUN8ML27Hn1M5lY3Ly5xUyy+tUBj
jgWK9LBckuwEW3jg7ynB9rzAn+gbnvA1IAc1VAfX2OXzb04c5PWvrwNrXsG9hsfce2XEPfYMOjuQ
KOdhvdeK9F6XfrRoEtfBJKK4mbHVge540KXMoGZzCDpdUuMuSG23ZdUgAvpzxxidw6Rb5MM1aVLA
Z6rl8RQ3I+LIeXDptbV3u69Xchk8Q+luvvJVGRVzdeO3IzZouYaERc70hS3wSOcTmZGplxzPAom+
i+WGs0/6CEM+K0jyIfu5UzVwPmSepwswKwJa5EiYLEilbnVr0F3v8DpzoZdhE/WGRmGb9r4VrdKa
zGvx2yNpGU/eVnmMIgaUPThEc9YfjnQoDknTJOToNwyZyFZ5BZ1Qf3OgIi/6CmfxKRLWqkRIB7K5
/v7IO04v+mo9JKbKqnSkkekuTfd8rAz/JEXyNEk03aLSC6DBmWogZihl1/jAQLtrNGjHtfT2Aqt+
uEDOsV7cwkAHwbgcicsMtToZewT1nMBYYvpbb653WZFYiRxXde/Ajtj9Guu6pfLF3lvaZmJPfdG0
2ZNuTOQAAfKbq3QFRxG4UBoroq16ePIjlwtfvjCHi/KvX/kWjtMkStqUHqdVfkmQe5aePA/n54xg
0MB4ydidpq4LU9AUV6t5l9JuMFOC57yHFuW5EJ17QwvGWof2NA/sgrslW4w7oqUNecwmAsqWfLFS
UBSuK6TnP85/qCSegUkLqhJRqFHLRSyFQeT0skI/pEu8/tEZEF1Cp9sCcDQeJFNAjmLKWConbhhP
ibm6R0VQXLai74N/erbECyQ6qDCb/9umw7YsmmON6YRveULaBBklyvR/GifeY1hAoZmbpSnQaK52
ACkcfDDQ8zP/lEveRuMp26D9J7YLi59xhAyrnrlps2zAWNhTnqzLR05tY8mSUy2+pLQ7uohKse6c
eAzTDcKHXC0BV/E0b7/TVW46Jflj1gqFFVZ5paTmOTAD2Fh3kjwTlcuXlzs8MRGRv6UKy2puJSTL
6MIbWgH7BCd21PA4J4mwbSugPQzTi6NkzSTaROBApPaCwjQIVxWZktys1juP6hzNd7l7L7pfOpxz
x8+WjsnOUBkhZyTMzmrKXAwrC5/XZp4xBa63e4q01nEMlOou+vcbMSwp7au+Y5XpsXyb3DhyrS5X
1N82cD/uhz8oYqo/Uh62bWMMipHbqEZwg3lbqRJKBFCxA01oU3ym5/g6kegn0o2ZnKVpeARhXm/m
EcHObl8QPAap/AwAqNb7cAlKz104zMEKtcu7Cao9BpvyDi0EahbeUMlkZl1epglf047xbuwJawk/
Vc4W3O1aOUeMkgdI+zbWgdag3t/MHgW4rPFstehykBGoL5Q7eW3qL2vEVYn/+6/S1XzP6L/qUKU5
iRGdHHA9UPF1Me4DF3P0mnMYGS6vLwxCCdg4i/Ya0tWTKdgd7Py1Oq74cx2oEK3SPOYyuKiSJBy8
yX+EArzjWrcb479gwDL9iyeXSHMNCZSVs4vpLR/B0iow8lRZ5zrWFNaQuj/Zl1s7FfQtHEu2/QYV
02yoqBXnHltSsxBuoNlc6sfVMkbhghn2YB1pEP8pIPMjTJNfzs3pxVX6nC7v+bZ5kjWZ0IKLY1Bd
Snkum6no5xssV9vHUBXIWeZdUzsv2PuqC9P6c1/a7NmUjGX3jPneiAUrYRxhjaBwui60k6hhyTc+
TB/sMF6bl8XHToaRB6W12sqvRPsRQL0G3k2xzXVgHUASmv6YGayLHjribzG7sbbfGyw7v01hYrRf
5KeHR4ThXZB9d0m/tWgqN63b0Of/mzzCep1HpyZFsqFMrsV+GVcKAzZJbnyHnhac/8jo7EYSEafC
+/U3aRKfs0izdeRpnG6zfi5eirQeryZV2f381wy+fv+qJFwDUntjDUr5RwcnhvOdwDBWNDyS6OYk
GcU8txxhxP//aB8GfsPHbLIv4bT17gyoLQUj7122XKoehuukGebzIk2PI16S8WMKir2r7M7E+ke4
OVOIO9mAs0zrN4VTK5uqNpsuGOaWF6YrKFsbK87h1lueYucAJk95U/0iRRKmUg1QTkouuoZoExpz
ty78G9g+/sapG+aj0cMmy7LnwdxH4ZVL7yS2Zc41ZQ0lgVUjPbL11mKG+eudjZIcaP3Sb5rAn+lJ
PEM8Ic5whkSPRwiaYbI/zaDjZSpmnPAy7509qcO/vdHjS23Yje8BP0K+OVt5iJmVJqNmEhiFGwMN
B1rEa2oTtZt5w/yNiNP5JSL3eP80f7yW0cvLhFpD0xtjmH8f8tyT3esiWGmB2O8/yBxwUVtRXAXg
iJz+zd4UQdqXMN6XXpyIlgz5pwVS7piidsfpr/1FDRboLqAPIZ+9oH+a3QwlD8lge6P0HCmyu80s
to425PmiaYcFTfRSOgeWwWkcmF98pqv4cOVviPd8NPmdEYi1TMLy9H5XiU0niG5N1Dn0K7f5PA3w
wGNCGrX7PzohhTJlr3meP0386uRNORj4NCzwqv8KHR/GfgEQpaHg919RtSMmWoATrrLZO9KuaaY1
T9iW2KDDyKV6f1hNAYsXFndBM/LY/U9T6FDoiqZxqEdMY2Dwz5MJFLUUJ7TdRYMWe6HKQKfeyg4T
lOVbK8U1HXnsq9vS7QhSbDg7Yzs/j2MLpdOjgFDemYs2W2jDkBZYQsMzSkdeFGr2wqg5sx3wTVPa
bTk24kilzIvWuZu/1JcMdBqARcAESpbRc++GrOF5CZmGhuPOvuZc7c7JB6sTfBQYb9CCfjC9Ritk
eHtj4tgTLsqUjMTsJlJNllpADHViKgbmHCPOqONLYvVp36qPrp9XKzpYgxHr8ZX+jsfgT9AD8I+g
9CoLKFyuUI78Ol19vv955/Uqucbqe3ovntcCPR3JjkGct+AnNRWBtVKE38qhwkeiExMH/qt9+fXg
WJl7ke1QQa44zxjBdSUmJa4QyLfxUVP06Fnfv2djO/MaFh/1i4Cb4tCecDojVk5Xt4glykM14j1Z
36M2PxCXqDjnc4Jk8w4wkMogqNSf6+mtZjfO0+ze1Gcp60HDOPsAdSTp/06+aJDRWVerCzD+QgJZ
q4/qBY/GDM3SB6jkkXTABCwOWro0aUikUFLDZvHSE73QmaRZcHkxqHWidhgbX6vvynTt1/VzMn85
1M9iU0Oj4m3b9PcHATPPdor4DahMXbiJVpvPod2iEqPZ6+P4pfWXnUc4vxOVWMxlSesVSPlmVu5f
n89TU55JET4CVeE2OKOJ9PFrj5hnbOLFi1rSrRX/NASN+kUngAALUuxIwW3K7MuzRNVLoCkhSBet
qDvbf7joRYNG4HMrRlJ2bevjmD1YMPMXyMztVJCV3JQvVfEF4op5v+3OSarZ2QZ7S1vfzVZ3CgNa
9va5IMQHDYWMvmVQUTxYnJV8uUrM3nxqktLQIsRzYWilbrMDsrPJK47r5e5eiROBWTvjk4nrpD+0
c707QNCKI9jVn0ZKsSJAUDvqZNCdkCpKeigozw20nnTaNnGOBhyyjgS6XxRitqbAsmiOpKJxODmH
S2nTRKJF0Olo0ullSSJqJLGTNyckjQn/ZV8HYed7w062ur6DIG8OI6a2kq94VvWAofflaS5xO7Ro
cQadd1X9i31Nuzw6VGf2V9Cx0nZX+CyAX3q0uDY0/jgYqCGxU16OstfV0e/jflHBMGyeEJZ9cgS/
y5hR+NNqDPGDXuVYe1pSQqyXuV7GGg9k9hEu5l/yHsGQTxVzgHi1FakVYDs6zXLLJ4i/u76JY26/
1RuBlirIZp7HQm+NHldT9omuJsHIgG8on/rRGw88zy/TRl9rV4ngOW3F2seju6+Leeno7qk7Ivkv
jYtSVnklFTXilW1rRw1CKy9UAd9SDeMu4r57gPG9fddsIqtnJtyQ0w/EtvFY2DUyJrun53rvYv54
gsNX0aUDrBGTs2I0SVMvvFmooIbSvtrVyu80k8zsXiip4W44fUhZ20jpaxdCvl2nhDVrHznS+Gj+
BymbnGplPH+GQR8ENuW4XG8izx7KLx/T3nOoMczQtlKq1D9pdXlUm3JIUZo8EkubVGmElZakCrbx
oyn6VypbprQAnRW3/GHAK0DubaLQQL9K7PzJ2qZsPyyaAXsMMAv3HuME3r4EmfZsH43sZnIsEZxP
ZnnkB4AQPQ1QJ+2mk5NK94go7GECeb8SgSdJJNmrsFPmmJscrW4kJWJvZmecT/9wAQrub+nA1EiL
UXuKQnP4A01fqkd8ZrhG4T/eJHgE0NODHZIDDi621bUoeGGZxFiMW1zW7mGid50ZUXNyDhDCAFOt
26Ra7n+FPaUskMZZRSC41+SpuoyxTkysBo91RwgAibwMHu2SaYSxb9qsexCcmYi+Els3UngALfF6
TtxS4ArWAXHclKIQC6XV2ue/Yal4jxqEM+/GtrR7u0/Y4btBwSvltr1PdjtA4Qbk3a8zSNUO8UkU
PLmBzybdIIOOaPlMKqbn7IlEu+TePCqiR5h7s5bCHzacQ7qKKBJyUohCGQucjwHORBkOSouRE3Ji
ShpNer1x8AkoSzB03SD/l5f1EK1pDrUNX+6J2bzoRKoFzl6Aiq9VJ6yzbfu86eDGsTArOAgUgz/W
Ve8h+N2Wml+K8COzFNA9YtRyKNgLqKOX/x7RfWbPYF3LnUiyyFvWGHduEwyjV1rklaV6e04X6DdY
39AE1GADVjOcvuBJHkWnUr4FymMkvQKR0wMg3SwKjkLHzLIcgoJWUbkdVk9Ioq9fdIOlSK3BN3gS
1ekWro0jxum+9X8U1tFs3ICHgCdyv5NFUuI4mvtZsCcGlj+vTYunATN/pQmiQk01Kf0T3r1XuIfv
84YddSu+TwO4PpO1d7QGKPOeeBJfReRx1qWu4mDaoV8yktPz6z6zyfWvoOCesWLiThnGuPmdCrIZ
EMSnQ0KdmJ4YDYt/34Rz2823OLKvuj7FHPHkF88BNUXm25FT43vqCdmCl9wFfKkjfH3U/q2Px72m
r1vsKmoI8SLhbHuOFaCnU+Twp9f+P371MPtEsnu78csGLeu4zfqQXT/SXDHrWcGCAoq0qRb98z36
V/mgzofqxXkwjzQ1JI+PUTONp1G7wQwhf7xKdvK+ulblXJ1YKT51KnqaA9IQb0iUlz9jBLuIurRJ
mls4WKZTYyncJTQ13t3CuZO4vHMy4NJb7EImEhYjNQWa3B3bWcxQ3NUf70aiUKQwOd8pJl5yM5ty
M9Vgzcq8d5FwjLdliXO2xMiHxG9uTW2WhVFU9JwqJZP5I7a+GYiMvIRPN3Jrz2YFcF3iQ/uQOr3v
T0pfDQXA+5o9ZtQTqPVY/CYwjkInF5ZnuDEKBp6zGNgz5BC4+D/3OsJ9HySVXy/86It9OGDy/8n1
aWeRUIYoJ7cCpNfLeopjLI0a7hitsRx/9mTi7qiAjLadtj5VLlLVqfQTbawdwHg1ijLBEp9NNuVH
0VyoudY3gAe6TfD31SFcry0DLSeznI+g309eAPTVeQhWwVnkHp+B/tirTjabyqiTjxs0tXypcz6m
wTlAUGBxkugQqzuefb9PKTxTV61RXKRrYxVxMikAefT0VN7lpZiHsu0ATIPSwtCuTAMPJ7M6vuOZ
9+DfW3T9Fbb3W2lRfspCdmiT+RN+aeoy6lLy58af9psI1cwkdgN7ZmbeqWdlwCyN6Utwm/vsq1Oo
eUqLC8aDnXkrC3C5BZlKjccYMhw5UTSmg92IJ8d6RjH9J0aXtSpfvsPpBTwZBOpzyylvqhvcAz1e
pgOmH3fdx94VZrLw5IeOCYpuHIYhqo1lTLX5UhZwZNjmT+fTvs1Tu2PhY6/d34nwmeMTO/ZpdxPd
RANW5qmuJzT8ewB3xS3tFtjgAyPIJdRPNNlJFUmHny4Y7nTmWI9+G+rXkqrLvCFvm2oOmpXue8pq
BWuPYruRZrQlvugKLnwdHVYhB2FvO6MP0ObUuwJ+1h35ao5hX1ClkLQksLpwZRUzPGluDRTZ3F29
dskqKglnVCwAlBPPAP5xEL92TTbVfEziqbVfjVaRLBfjW3pOQ4bpumrjvoOqObMQOtBe7rAzfoH6
CyxOKO96SnxIo3Jft9QU4f/JlrA1dQr8Trx4LYwDL76Mf6QpiwqBQ1Av6NkNWRJxIf6PBbanU/hA
px68ylAFUVyaNbSwgddcDRStGVal0SjGnf+jdz+1wR71e+nHJC2q1qP4zQJynZ+jnUBKmlQQQ6gl
UltTWB3BryWFp/6i2f9xC7plr9/ImZCiulo/9ylfLSJeYYCdEtfWm71HpI3VGle3ADMDXlb9142y
yH9Qn8OcWVnApCtaDJm+VlpjoMosBlFq1Eq0XFBV3o0bK/bB27H73HawpjGe2dJNFVJ3Ao/57VTr
NXwTHyyJqWbIPbe4pwQjBVvP9gMiwzCtjVUuuVWVVLzf/0AbRawIaFoRGlmngIglcFG+PtOsxwBg
YPiUFhu8iGKXP4zpJ4Ck/khCR3MWXZg4PH/vTtGrwJaF4mP1cP+lPLOsWyBF/PvTgFJXErXrHQH6
sZvny60BbV7JaFKyH18ezJYaEJyOYRcgiLLYeObEzex5GoJvaOAFzx/6lzEU3lBlDfAc11Q/qRXa
Y2bs9P+LR69QBjwNiFAegkFU6sMGJ5mPiqNOvcuoZRFzEoFnLuHvt/yKuUo5yljH0dT5U+P8GfqV
e0HvWnXbwbuIYq0MHVCeHPN5B7Q5/hwDOFRAhncsjaWoNSRuONmMsIjV+IT9OiRfnk9+zxullxi3
xl0/JExWeN1mYAo56LlvvH8psWkd6gCjujHHdLSecyJfFpxgC+deOCPNXGAOu6v8lKD0FJdvU3HJ
Q6Ubki3sNsbUrc8hI4Dl+yKcfD+EAYAW66NRxgoOSLcSEj7bYtbqeiT/qlWYtKpxcHOFMf7Gr0Te
UZsHQSZsYUy89dUr1ewByzXynIM1xnHlykAtAv9Z9u6dkDgIANF9CImRu8hpvXqgiv9ILg4rrB0y
HHmdvV00cERRERuCD/xjmYfCZkjRJ9ssc6K/shxcbwl3K6R6b6YEkAPVY4oz66PZt3q6ZUXYRswD
Pk6nezSxVK7IDgXSuy7BiJt95IlSGcPYfit/8Eb5pBSept/k3wQPZdYLgvH4iC3FjJe/a44BfFZw
TOW/QnQGUY3lc1faAONtT91zfCPd5AxI7JTl24RXhJz9Sfk8bnwZwtKIiADGThmNN5VlwBjBMQEj
h5aZFySzug6PbAlgyfsVEf9vcMidctQE/WWBl1MasbCjHCXXhWJxvk7xDCEZZBSc4lYdr2KXXFzS
zDke3Bfux5F8j14psEXAPQTKgdMEDdoM2BGunmqxa+swSpmw3OKp/D1URcuFQ74GBwzxx3pftG7K
b6eTgivihtmtezPIg0JjjTDJbDvGoHp/rsNM6ZEGQ6k0byHJO5k4sV7zlK0pX2nqaGqCVn++3woe
e8rQamc5x7RZqmXcUbxSDFvUgSzkqdMgjsrO/xA1Qg4Mvf0bGA6/zAZadE3jKhUEDifIMGKCs12i
Kn5Nmk4rT86IvNJjK7wr3424ucEZTy6ThmxUeBQQEOop++XQga0WJIplRi/ySs8uzeH3lLlxiw/V
6x5VVkiA8Uy0yyZV9qWD2rXiwHo/yzgGHE7vdv9xdJbFzGMfFed6Y5hGfkJpoYSPpFT0UZnyDPY0
jnRT5av7z4O6gGShoB1Sk+dZWsYcMCIK+WA9BWBrA70JynAUgt5D5GqaJQn0TdHCja0/GoGuScs8
G6seyLMhDiFzYuDUAk1Il1/dFHy+a9Jzs7ibCzPH3GujS2qp5xcYn3qzzHfaJTYUCnZOjC6PhNtY
7IBEME9xUk0C2VyP2lLIvdCBQ11QuwieVkTWM29g9ICsgahgO5N0DP89GqcOYun+EU/Dv9+qq5LN
n9xTlJItMqcaKEBs3vobLQqVvAKBLbCKtpvCbiZpE7I+8pN5+lbd6s93VXw3v+cS9IVz7QND7uKP
pRomy2QbQ7CpXOYuLGiXL101msADUKKbBwI4r0vzw5/aE06G1KkBfenb7bzkX45AGrDFa4SGL8wx
iXJJHK/RvuI2aoeYXlMSmG+4Nv7Mf+jinAsb2UDPbOWHtNnSPpapYle0HqNbpvibVSqYQmrJIB1C
3rdJkGvgYHZZnWYMm8ox3hwOFJKKzGeCgrC/FWmVf2xwVJTG3ExKjFrLHOVtiSov09an0KnqX1La
4vNbz2VKZksI+5jj/SmMcxSKJBTdnLTL6tk+B4FdIqYsNGbnb+FaHyCMT0lOxJRTC+LutIN79BnM
ppG1VY7EApuOeCR1l/1gZOb3+vxs4EJNXEU4dKWC4G20l3ASVcQvttn+ax255flRGNCjY3vBHyB8
1akDBTBtChYmfjMdMDq5s2mPFKQLNIAYvgtueXOULM6aSvZQ62eykOMCkiHuxLwXJhRt7ppIpod1
Ag8XfPZP8IsDpQBXqKw5C7mcRP+9kl+f7mOkXCHDFHmlRCe0k5LYVu6iF8FJGa4P5ZSB3zsBoTV7
VcuXC1yiEppytQjMw+ULCe6l0lDFnPDACgvFP9fpr6iZqECbsTNFJq8HgIbQA+pBH7X1qcumOFWS
n3FFU5rI8zxf0Xdye3F6TmCbYbGtuzgxz4Z4i1XJzLtltN+QwawlzTPcrqnCYlsDeBvGb5QuiMRc
4dNCsVvwINi9gpUxW+cMA80bE9/ann+iwaFlBYsOx4uuwZ/GG734Er0uVLNES0dGqlxkNN58RgsR
7g+Z3JweF8Jxmjn0EOEg2OGTQAIKNonArHooq31/eK3ZEzABZuwzvzMCwmLFw7egc8DYU1x4nZGR
YjdS2njNPfp7IeDgd32/tplFTXK3eu8Z2LYTZykDsPG4ycCOApLhzqz4EKPlNp3zuNXKOAxFkFH/
gKUzRT9RTcPrOilllTzU5N/qGX24aaHKuxZ/PCn3PqGjy3x21a9/20qzt+J0GlYS2lqn0NMyI10N
Utydani/pE0BNby/yXHbnCZxv/24zlZ3NFg2AiLhwqiXy5BbnGWs86Jb+42iFTk+RI6/vRqPN/n4
5Hh2yBa7Fsivtm+sYrwnVY0AgI16yj/2iPukITg/fMZkpTZnbt1y6UfBOy3mC/pKvs7gb3gDzaWY
rczoxJRIc7W73dj8ZEN5E6YtobB4j/MuPWxbv0/7qGRfYHtJXF6Xlcg1s7KeaP2FRtB43lMo7YWL
T2erXyHNX/VoSzneBAr42TBoXos32FPZVrrf2+Eg4t+CmMNbLPba11Oz4a+6/ixAuwijEtvHTGL7
BanmIkB6q978AZBDUy9qitnwIwVuQT1Pd/peYl9gpeRiMCIDdCTRUpbrz9SIzDXmRrE5Ep6zs4Ma
iMHbqSGOPXd4ftTexBOMrihs2tKG9iF+EFX/Q8hXGG/IXU3KBJPnshXVyvAvUTpIyopCw6pBs1AP
8EviOjJSJLIrf+72L2gPND00vPUbdi/MDvzdaWHjBMrqRYJQc4vXADL/qPgsOusWLcRx1PeltrGh
TYX5W7q3GCmlMUAP7SEs4mlHVfnEcZio2O4ldCEuvUsc43f1YRvl0tFJMy/C93S/AkyolbdH4qqN
KuJolbxipimmQN9cEaSR58EUB2al5W78yk+qvIsosPvyh1oibZUczUjeRK8MHfktlt+vcpy6m5Mo
6tEYrfSyinmGzf6OSQZ3I4peoAaqJvPsw4+Y530Awp4KbbW8YDoNsmjFpAEVI8PERFv1KxJD3a/y
1aIejogziofoIcN2rbDLEX/SVtPJgY7XarpfED01wzEPVr4olPw/eeSv6pIz8nZ9DhLGH68U2iph
yFGIcQXkW7nlOA2smRwHwqQ3NV4Ru2eQNPYqvMNQZwqgup/5lcxQyYbt8Pcm/UkDy2AdTQ+EfPtd
+nmB6qdQDOcNrmyvKnDwz9wheLD5OOjO3KJuhAxeiyIkKQTFbCdzQDLD6/XsZ+fhn7s+jYo3mLG6
lyHEbFEt6zX0vNzFYq1D7Ahcdsp659Psjw3hv5wBVjTbUhOEPwYqreAVhmDKNARBjxTitReH65i/
B1DmQ7e6ql1iAaALA/Xkc4Jr2IUA18F4udChQFSHFnVbmmfKFOITOzdIAZUTkMFANtUFvPqR47gh
5PpSwRoT+w9NbAK4G3LZ55F2zUUrSPQHVBaQy4W8j2QdBWvsIp7wKT+t1pa53jrN6byFZ+HKMgW7
oFTV2U2jAN1O19r8QqfHFpiVOhSYUbUDTYpj08e0164mH7zd+QrgoVL5KumFByzH8mjxBGVuvCqK
s5ZqG927AF95tV67bQsQs2V4ob6vrcEyZFnFHVVP62VfjXlEQ/1FeKVRrorAHXcP18bzcS7/dJJx
AjW17olDjR7NQ5mlOawBJos/BokTLd83IMks9i8GCOe8E9XBGKhRun/7jO9+CYXWN0mrxnqn2Wl1
5/tu/5RSgG7KBrxrBd09Tk7Q1viRKcBjIF+kJFcHy+HuGzJFVEMQ3l90PyyrXZV9lvQJJBbTkGr9
fHTeu4/v9oNJ44ZIcoYUEUxYq7IYGaoqKXjOdFY6Zz4TpUhzEMHw0JcCPFd9Ms72qY1hkYz610px
WPS3BXftRlJW8BKkjckWGPZ9LD8Ty1SwcVD6CTKqGEIq/qPGwjOchMCQ2RoZulSuJY9Y0OoJy8AP
SBLrQjZMGCW4eo4UILRTCSBwyqn6zDZlA66fH66PkEArkvhtkv0awJNmi2n4Eoym2wO7TCiDNeri
NxVKdY8hyi+ol8p9A+LRWP1wwWyC9tmhgzOtotW3gufoHrCIglT5WVKuYIdSBnMbu03TL12rZDnU
v8IMI3YCJ2YvTswnW0bS1Xu+hLeHjJSWwMuIJNFzWVVmIrW70YUmNORMnzCWAWb8igkzXzYWWXA2
ooyuMc6vZ0kupUZPyPRzWva8Llr/hg5dMJZAWmok4MrkiaNLP4ixOhfYNVMl4cZlFn8JMFNQ+pft
STvSvI98AgieIEKsVizfbYp/BFytn4Ln6ipT7X/BbNtzmLK+zO9oQ16k0TKQJdQF2J6jx6daD5Cb
R4EzM4MDuMWqNq7jFZSQf8yAj/521kOmRZV6KKha/3sIRdEG3+0r1lyUEdjV3wLKCDTxSq6+vM15
H06VpBZojT4wngBxrPkPDlF9xaTFFiy22e26RMN43h09Ps/fm+LTJv4ydcBFgg6u2z/WIC+EqRWS
+qh0U4Kn5H8t4zLGCa7yLDFpZLV6YUuVFRSkzCEd84pUWi6t2B9D7BTk1h9PSUA8XJIbYnygFmKe
p8LtGeO6/dFmxLIiDz3KlvxL1GzwN4yw/gggzfUcCZIqSe3enZoVOg/5Lsji9/A6gQ47O+M5SNmd
5156x0HXiTa/xxcxhQVAZ5cjRmnFy1VSowlYeCChCBkNEnfYKcexTrQkRxsxlz+fhixxI3i1bAUb
n+HDFyglaHkZ9MdeOhpB+ZRU24nsJNVycKMa8UM5qCcyLLofhLDJXdaxcjfy+gdoPVV4uRp3RhSx
pm/C4TdLmhFeQWAYQtiJnJHQ4p6BWRmMEzmWCQ8ysnriXxTjMf4HQj5JTDL5DMlbqUWIhF/ddILI
dsQS4aEjnrSt5g8ludtUl/1txt5/2PVRWYvb4RIQVhoX7AddvjVFDt0XbmsoUmsRMHcFjIoUhYRc
uc8dTUa/o5SSg25i/mczkUphjPTF1LoaagNP1ZDJLh02+vP+3yxwBImbXmUA+KnxfDx6f6EpcZhI
vKXrvJRkOjbFXjgOpIG2nkXRUbsFv/mvaI378mpI+Rmw4oCM8I1s00oygZ/QTADG7Kn4NtGkZdlz
5KFhenHNJtfV0J+njAYEZeTgBQiIkdIkGWiqv+I+b1oJKAqXbFxN/yBYs7mOkAeiIe/EMw0xpuZ+
hx1O2susAJJnOBPpEjHFKf2sfbPGCa+/GG45tTlkfuv4BUVo8Ry/WiW3f4yScFbeeCAFngJ7nyIu
kohOjjrg0MuyYZogNFlY0lEx4AePAKouLX3g4wyw1NuxERtwhi5mzMpVWkE45uyAojXzgVt4KQTk
6J8KKPFFdf9MUkGVYfLhP3zdhw9IhyqGYkomeqmFSe9R2DmwtfCgk7I/RDtI2qsMdRN8X6DS+dw4
wY4XY+dBs/y94va6vXVcqNEa9wXOL3v0K9czSjcqcjkZ7W50hXJfMOs5s8qdVHbwup6IzBjMHGsk
ciyTCYzmfGketRb2d2L2I28NJ8MGDZhNXKYnyiP9GUZvOrr5F5NCG9MP6HOe9YHh49N1NDE6Y8L9
6Zk36WjsrQk/JTpcDFBVWDLk98+Hfm2IwUzirT2o8w5P/igJio7Y1IGHZQoXX/ONBCQzJgLs00Fn
+sC2LLQ9VgczZlNlXam0mVWX7jj0ZVFS4gEPehpV6o0/L1Tvex5BbtNEJdYZtMkI3ws6YrXmIIDu
58pSilLQ9bCtule/qQ6bBd2RIgJGXqHwLZmf+K3lDu/fzzOkvjt1Cf145VcZmF5Bjgno6c0x5bup
Cs3ItBTCrtwiUisKGQu4e5JjKq2f4L6pIha8VgvPa/PXDyxBI+wG378f4ePVywjgx4SDMse+hXVq
cD6Jlb55qV0CljTki9g+0VKDHLw2L/yvDjANCA1vQ5gLYdmyI0JrPNh2oiS97ruTvJ5Cwa2kBGQ/
jBlihlOaIcwXovd60h+Uhq38VLOF/A7er5XL2s0xxQPA7fpJHWyLIyNUdBUM9KU/qNnsKDrzKU5H
3uJ3IIjqdhQkSirBe+b3KqQKjbFJh+ou0oqcIlQqi/DbGT9lN5eb7lSp4mBI8dj12WVhCnzPFEER
Lueml9wcXGmwba1w9UTRDcqBu6lsGuc5XdYM9WS9L0dcbtEkAXEQNUk964L4ZR49UAr2eQiUzOvi
VvmzINc9smotz39peyJ7C7330hL4S3yUsYKOA0a8Rcg5x28zZq7zjYkcy8s8HHPcIa1XapiuU1Ky
cHSarfOESUtoWu1fRkmg7IVM8gYL8qKsckUMyBTw0nNbWKYCPudhgK3XhRZEOYdt03IgM1vnMEsI
Ghxt1v2KrfbXi9q31CZO9BJEWhdNe+Olq1WN3QfuxxyXYzkWaR6NvePF+6Q+PdI9BeYs/NeXQAiu
YIatxVAHyWTobKhjsYQJbHy5s41TvnzEhgKFo3svq+dG3+TMjQ9j8z34aFp8ZpLsKh2yA9NN9K7F
vRTPIaWuTOlwvfq9gmvRYItoFD2DCOh/i4LSOU4i2mLR+IeyEFIgWylPyuKFdaS1kVbXw00BHmQX
46B4oHuiPjoFSIiEHuSDCsD0rZDd6Ocb3R8ihLN7HlIV47C8YNWRFM/LZFobwcl/XRV8PVGZcrrC
vAo1nWFOA1mBtN2km26p+9PWd3ZPRugtEoJ1RQF9DWfk4qstRvDSsk3SXYwOXLSheai68EOTIzn9
9NU7YRv84r38Uu4qwf43ygo4W2TjjdaVJNTCcs1OYH6Mz7xtmuhz/l7eNmsFmCdfttSeD5DlGSc7
VXsRpHo41W/92KHTrFF2/rPxcSDu9BSnvRVoqdCC+lSD+uv+Zbj5Xwkj7EMQYxoriBr2qzUns7Fm
3yB1rstlbSKq4MQdrvXMX/rT9RU3JKE9OfG3JpjlfNH5PPi7r6fRn/wMVYTo7TXEZ/LOBafpmEoW
EquLaisTGEtBvHBRTJPT496uW06hVZ6MG0IwbxaDvEpRenGPzY2UvF3gQoTZzMkHqUMvblPExWIB
hz7Q4HVkVH49W8kQk/5CqhYn5zUbkrAjA6l8UwWWGEd5Ne3ycxKLFqvg4nnwg0h0bx4jbT3OttEV
KyFIK25u9plEsAfdz1O9JDl7IJNkWu+lkA59uSH146Vy5P/CMxzlT9G5TrQJA/RYCbspK2UBB8qy
SeSCv4lwd0+aAHR56/kiwy+HgP/2rwVHISitECuicxN2GZGykqT3ChaeblQNBJSqhsO8gJ8sXGay
nyLuh0NO3Qb4VnBGMI1eGFTN5X6nm3zOVlyFIGn6MajE2wja4X0YIRc+tJqiZDm2xtsNfZEVrQ7f
8J6PuYw09+Qk4Y+VVJYL7ONp9KScNBMbi5QH9yzdXoHqwmwXISyL0Xh1P3MGWfE7l5Pc4Mf7rUMr
6jP1FuKXd4hkoiicN4oagxaUUd1oeP25x2sTNcsLHtXtz14/lD8EMdmM0tKqomgY+2ynCgdmGXan
GGy7VjzgpZtPk/tQxxNB0GcAya/8sEM321CHtsNjgtJF9To5cOgGey5QKgRQDK9m9I1VZBXxV5iG
aAEpbS/jS39hqzdtl8oqIO7Twk3OMn7g2sAc4sqixOZHgGb16sFfSt/WW8sDdRHKdnFf2W/HS4JC
qjA8lleBRuyRc3o9mX8oGvZD062+feTkeSS/bYWaIhhvHTzbwO7fNpsH8Yanaes5JCFnlBlBSaRc
3c01nreMwhh6PSLRTa8w3uhO1dGG8PynN3ZbsbPyjCsYQslcl3FNGxUz9z6pGc8toLs3qU/W+XCK
URU6GvOi2mQX/6cCwKAUHEdgL/PvNu/Ezwxq4Z0BDlagbrljDMVpFCqjp71kK9ZESnrGRxRdYyUV
YIGfL58/Q6QTz3+P5tkgQX6i40/wWsKFZxNF0bLxxFX2BDf4avppmP+osz2gu0FCCSI4Fn3v4jAI
KlCBsPuDvV4+YgykkYyusYhn8r/E4K8fH9sGqQdpSddbO4D3HExeXskHYlHZOnwlyBsNzEmhAo9K
UZacTXPacW1SHqB9ge6z1heLJeGmUfb6dRDj7B71lWkLqlx7ajtAzSupyZ91oGASC66+Ou4UklkX
vtqeTYT5PHQQcO4/ChaAhY71hp/r6p+6Haf4NHTYXeHZ2b4ECFRxh5p3qTVm2mgyh21nsimMRQB9
VfeHQYBtN8Feg6zkj/4UCUBxHSiwM0eGtjetAIlOxiogi0Yg8xlCjctJVEQOFP7pDudOKQHjgxJF
GuOonCQF7LYBLsxUs5dzbktelP4UcGWh0Th7gs3C26PraP34J5K0LgDKC6qOiQTUfpMChLzW+KGQ
JCnsZZoFVWTQ+XRvbH/1S005/4kvpLPVAaa0q7d89yGDiPyNmo5uWHBXNM17LObkPvOaT12ulpX9
wIDrSjDcxmr8NMWK6VpUpGRm/eCLnEldrYvvfDp2rs0t4hoetlr5aAgehDlLPk9UnCKK6Y05m3Fo
Ui2Z75tfleT3EA8q5drFC7h64rpHXFCi4qDxjtprqR8AYTtfk+HFSjRa3UWfDmkvajTFn7WsmX+R
bxNDi2EIbzXXBGnJNU3rbwyQuQC6lpDhx4F3744gDx8fLvPGtYIULotDC+O+EY+YJ5h6JCoAwYKq
kouVEgYbM0HskgwcUJOTO+5whukogBaD3pYwxsLbbURJyGch3nNiEj1uWIGQJcgFlNGUmZBYvELg
L08nfJ0GQ/Z1h2RfmuOA2OSttKPyGFoUrAoxSLX00hMWumqbrJ8oAH55Ye0Ti7ZmhQJzf+646Qb7
Vc3jMaw9epht8BmDVzxDni5jfhqm0kZ9o8cRCPemLg/+GjJqAIBrv7pv3pAyxyrpsGUXCzVIqee7
RXIIw7PXh3Sjogwanr+odMsPeCBv08sL49eLgxcpr24Ehvpd624TC7Rp2IjlwIqEdhPNziP6B0Fl
jpESCPVHAcrwibAUm8tdwK98o49yDcLz6H0mNzcmCl5F1fRyIB2IPQmrdHK0NVUzoP2eaInHPGG6
6PpGnOQLGnH/tbyXEDMOI/riRymYcW382R6bt5MyJj3F4bnAOpTDAHRnXYT0he6fZEzspwt6sk/W
C9VYkaizBYpbFOlhL23Ro6L3tvSQf987k4kxbJDVEaUJQGo4NMuJBcAx+erv/dJmQHRpS2g8JRSb
yx6ARJf+rcnS9mrlZ71OxeGyPe/klJfGrV9kcUJPrTArwY2cEYkHsdXWaTy6EuhkYLAMsN1bWaXa
zGtIGsqCwr0QF7Qy8wvltYMF7pK3c68Wx4h+P2xpXsTdbwWwcC2QDEVVyvOrI+KCKEvvLzHsRRT4
KZorDkSwLhQq0RE6fY/X2HCXrW3FlW2e6o25M4gfaGpuoUeFXgdz3lC4I7pRVkf3Eej6JG43T4hD
F3WAp5rE/o7NRMwUiKwcgslAMPXYC7BbjXqf4GXp/LzRPlN+6pJkfQzzhHci6avL2HdXUkmE4/S4
SzfcoBMSxLoNZynFV7XjBfZ1Q+u2GsbfvdHqH2kvEItBLN+pzXCiDzilKotImTyJw8UdFusbvUlk
Vos6KrJ0mjJuUvCjxhV4UcczRmZ4VOTqu8HvdM9CC960dConoTsC/AENxHYmDGpf+5hD4m03bKva
8voTAxRWfeQ92xaGD34Ywicu0FAB2XBhU/RnRNsxPNIjh5I50JVdpQdVdADy3OWjV+3iwcO34bOI
GRYbqbu7/ZequBjS0NjQXldut/j3a971iZUNvD/24HpIIPukTquXASccCbJxtlhehTjZAESL7NxV
BWzcnPoCxNfLEedI2ppe7xwcd3Dw6MB4TTdYZaMc5G5DxXebpbbvVQaViV4u/BgrSQuCaofQZRCH
18GoEWanuOUSo5phF0cOO6fCsCRUhhEzKreHWVKrvHokrxKdN1C00M3LNsLYXljaIu46aXY4RbK0
HqthLnLm/prbPGN0WNptvamopZxVrYRNcHh1MUzn5itLscSAqT8hPOxsca6rA6N3oM+Tgpxsd7dD
WsfMVPdU99jl5EvN8h8KLDRd4DEtdbIBcSe58IO6H2zDXzCEBgtqKgijyLJjsMS1exqTrwGzwXbn
g/1CHkgnSt/9k+esBWIbHlXETL8wpJJRgXsMpPJYb8lGm3ziTQECkvKF8hwxwxcWX0m0n9YHp7/H
p4a6yJxWsgNrHW57RtSgkthAcyejbSyAbhJlCSv9eqbC0fcgn6BmbU+KgrVuz5ZjyruElpdkkhaK
wxnNEVqY8T8h4FO0gkRQmEKaFzn2eNQAirpcI8wLuMTkOZeBfFqEbN2khVvRhHkEFjSiqfNoXACj
0xfOS4xWcQ3wIHdci3tOHUMuLq76txie1rCZMXXU0+cnT7yjKMB81QzfnIwbno0EtPKPbthaGGc4
+lwehdNjgVvuxONNHG27xOBZdqkYJkRxigYYTpv4JJSOQJETydi1j3JvK8yhjqx1470lNSdkxhv9
0EdRC4cM/qxvXR98ub8r2grEtbb5ZyQAxcH2kQLZkulMS9K9vdGm+HWmnV+nUi15wLdPnzT1ROOb
o6vvBEAnoz3K1vhlIZr4aJjivCJIvZ/jrDJVHVNfD+A90UaPQSBFIfhJYVv3xnnJrtI+U7XZMtln
ZarvoRvuMf4raT5s60O+u6emzEuhSPfT0rjCy6+DH9DTuCVlRBUOMa3bcLEQeCRngsX8MNnql/zn
umtm27Mg5zuCAVKZyf4kQECXz6x0kyHNNao6hHOqAaO+qNqPilusEvJbMybVomPOh+7QacQW2Cee
WE++6tYkfcGgJ4hnty3JgxqhRR6OFB6+UgHy4kPXlHNCjRax+PzF4EK0437LxtUNtvWLWAbe3opz
RtupRdulSPs9IlPtNjyk62CCixzyz9e78G9SCNjFppUP37/QEUJtJ9bLm4ed6KrZM1w2I2Lgn8iN
bMrnqh83ZkVBU5SXL5Z6iymb89fIZNyIsM5vA/nYekZNRtfinNt2zzLSNhBnT9E8ysHvA+yloRa+
tH63Zsxl8kDpQYmsYjEPYH1CNIBTsdN1hRJ9Jf3Kd6YMAYUX8TVXeuG5tODtohMyUhBawsQtzfnA
Lv9YcLAPG9x6psdkn8aofb94nLsTXotwrI1TobQSNcD+8MeCw58RwWOJjWGVB4N7sm/U6u+vm8qn
42ll1C3Ydd2GH1YhG6KxpY+GiRMEOLOiszB5NvofgcpO2Q2vbr3uHK1N79DS/Mu6NK/0G6d0CXDh
zRm5v5ZOXkIO1F2uoqQhllo01znM+s0NjoefMXzaazbJL+0kyfPX8J6tuZqq9nKR0cyObbzSbV6T
b12gLtInLJKUzSRmo32CCPhI9sfpa8h78q0mYfqciFeNGWCyT5sqMwaDcxwuO8I7joq7UG6Gg9Un
cBsnnNqQyJlvs5zcX2Id8RnuqAsp2XSfIWyucqAWJ7NDQqgwv1lYEuo3VSPhpBqm+/D8uH+UJpv0
EzEJLNO9l/EcDUTAFI8PRhw9a3DMfUvM+VGOXVr3/cBD9U0+Onpbfyf912ajLAaT9vxu+MU911ns
pwT8gFIwFtXt6pCamYrVhE3cPI2eew3J+sVTmxYiU0sBrl+TLACVK6UarrpW+fXQ6/WM+CA5LiFp
L+KUT5O/Au4mPaG5lhT+5XY2HGKhh/ZGq+Okzf3Rgq98WdEJqyOubHoKZPOYjZy/WPp1HB2FHe46
RoDQIp0Ga7wR8MmpYhqdB1rjUZlwytpyyKPsekFQc/JztFXCBJMLtU09FPqhdyKFh75CAuxjpn47
38SnIIoFHifWLaJoN7G3oTwoith5YIKjgwPtXiVzyRASW3lBwRlktYjHro9iQhumemlYFXjH3sfZ
x711323odN+yRq11bbT6zEhMOeJX4vxvp8J7mQCkGiBvp14RtderBBIzjduOqpTlKZ7nRkYg4/DL
vi1ZpzQWcS+5Sl2Nui2fUpFJXmYgS3md6n9/Hz44H3gjDAXdcERY+7YIIz5zxYdJ54r/YgVh0I+o
l6foJwYgqJjVP9phopPopl4pN1RTqZlyZj0zYZJBNqpQBvwd0Ap+9s1SRUjbIEZmBih1efqEsoQ0
sOjhLwj+u0To/1ZbFfhO3SQ3pKQs0u7OVLMsdBP+adDs7NyA/Gr0TebxrX32znzdElyVYx1/3TRY
5/cQtEG6mEatOj9zw/Mt2GVWvFTp4sdsIC3hpjyUVMznEcf2Hc5Qcvzxcy7VQ/A1aTPz7ZlbSR1l
vgYyX1xyDkvOTOHF3jgxaK6XdfAxdGWYLJVe+x2pN4fTRbkdXeFe5d9V5MeOE6t0leuvGvRXapgC
U9yqBg185Osq6skNJuskSS5VDEZp25Wf6XFkaZM0vloOECtFjGWvNStOrFVKiaMe9nhnWKUEcd3b
f0EolmJwgJ8d5nj6E79exq3L3SWNWCnFSmQ2EkZipzwiXHhHm8+lbg4BemnxzcZnyux2Pvy9tWsd
Fqi/mBHzt+SDtqI9xGxun3uE5Au7V+xNlH6bArVDlMB6pjvYB494saXJYvKsViSf6HAbZy6GJsO3
bFtWFMDmQc2SwM3PGpnq12PHvy6YzF+oEEZF9HKy59EuC02i5EWAdlJtLwodK6T1kgNlaz1CHFUO
Gb9snxFWz0nQlzeMrQilM6ZESatkXpJljf3Z8Cywi56Ltrlcl6OZjOtuSITiL8fTKe6bUNr1VWFI
pCWK7+Q7WMr8/PRqs6cUdoFPmR+xuHS7KvDhotml8FSIbhfQp82XO25bXVthFXEUnHLBUAJna8F7
2THLW+QyhjINqepo3G5zejbXwYwbTPWenReI8JeyoVdLaK1H4Z3ObAaeVF9OwrZ3ApyVo6db+b5t
2EdkWcOp9TCNHYYs7RJjMvHbQFVn4jR3fdtKvjoPnXhH1xS+3ZCNCCv/BDiXxgnngXmsOSw0RBv8
ukD0V7oj+y/CB/Ac6X8uRbD7ne/oyy2U4DjGBKlgwBLyG6lHnSmwcLbGjDOfgMkikhs/B74gJq6o
yw6OzRtY7JVGXvLlwovBOPlgw6n5Wtk8595FbF6iJn6S6qT2zVhbQPAj6mVy4mt3LojqR3kud+Xt
ejLtz+cv/K9quh77GgJ6NmLxl29n/3ZQ3vPFrfc6m4Q2MZvpeFhkE1CCAeBug4dk+9j/8i2vmhar
Gw8W8rqBrHfutwpnx60pbaHzxZ6Sdpshkr4HzEf5Lo/aHt5arpRxmiY8RZGoFiOYFOcpg6bqo2Wp
E6FsTJUALaz48m5rlRejYoERJDPvkm8OQ6o0o41pP+qiy2X13lrhvaP/qFxCF0vYjb4shON8OydZ
uoMHqDtZ5eNyfZdhjG1oLBa296iVamfr9NjleAt3rsjqPwQnFws99cs1Mkomj4ziMq9ai7podbNR
eengLkdsv3mM/L0bQPwbJkWHa8reptzrTZwHzQcL/fXhGLfahEpFj27bC3//iWIGActVByG8V7sP
FBi7FwHK86JRaps/h1eeUNA6qj0tyrHazy/yp0e+m9QjRqykgfUXtJiNpYLJvQ4g5nOCblrKh6tA
qNuu9gdozQNskT56Z4Muo1ePka3RegKjeEKAyNvxDTjk/8JOjMEn4+5LP1rmCxCN4XvzqwBS4wLg
vRkArx62GNWvcTy2pEnsqS9RfY8smnn9qLIN26Sg0Z/r8ecwVeSLmnEcwbnqvMZpAUtiX3Y6Qi1m
zrdA59tGjDcZsIFZaNIU0CG92K8k4pW/qwJd0pGDqkB6oG9wLKlt0itgh/n5ieeJYvbapuT2vt6u
r2qclcmjctmTm/rfZYE15Hn7c7Vk8gCIe/WYZLu87tvKY3l97t1enIjih6dwt1hifuLVd4dBzCs/
7WHy4E0ZBbumJihAOt8t3IP8gPaP0WZG+RMAgvbt7D68lf+7X3B1EN7fqddHipV1zosRuzJVGcle
fvYlktp17mqar33VQULu9K0L8NYD1LbRhFjSrjuLaBw/DSlxrprB9bUm2SyEgAkVJjYVvz9QtZ8Q
g/MRe98iWeN95BZEFGle/d42TvNdZq4fkfuUuc6waLc156Hwj9fsMckP0DGeTkByzQZgkR9IOgLG
Vpva2GEYnKlFBO7Z/OhFjduXUAXekBZA9vArpoNGp/dUJgzKU4DtjdZDqG9nCWshGz+uwEusrjCH
Cx+lP7s/ZNWfWOLeOklChAxcPY8zzjYczGEup2LoU9G+XNIDkYc9Uaw/0SRuzdGAe0lF8cmBBnWk
l3mwHfnBtdYRE1Ed3cfhMMX/DzQjkafUL7Bqf+syj7/DD49z1XNwDO/QNXI2bgxJUwNRT/i2/0ce
JXAZpjEZtrgmR1WQ7lnH5q8mNjeD4j76Ph0/MH5jv03OSPQ/wnedpnZf38uC9toFnJ6LYFut2Jfe
gU0zn37qmtt/NIY5r7rTB79+3vzauEGOJPRbCzcd/gZGyVgaBhiQwz+Ul4IXhoO+vXNxdiZCL4Ds
QPcDc52nqeW9J5BeJi0VjUR2OrcHZK6San8G6W1k24KB4PTpLG7XubQHZUGJ08y/aYTYjX2kgKCI
96YbGbvIpLbEQNhA1ddiI1ziua5YQUFyiPe92ektJhWRzYImhRQUddyb5RzNmFCdCfh89fYirTTI
4LHIP4xcJZz0njt9m0kX4Oc+kkeT60YFU9x0UPRNRQV5q6B4vQOm/UqiTXvjbwxWuKY4ku8kEjMO
pICP1tKz2DxFChz96XyNZR4zykM5uySU7Zxb2Qdc0SfrugCje3nedqScWSr7HVyOYv2Ujn7ZbDj4
SdJek5d/AVvEGDar1EiWW9pVAoVuVSJFYtP5zpt1NZjYxef9E55Ly2By0YpJUguC6RjvAgowjPtw
8Mr8HP61ogZ/+a0usgxbrKdbc+k8gNousHPGQdaCjg0qOLHIsGmimMBo8X5xn6mXVU+DUNFEjhww
G9N4TpC/c5fh2lzEC/VhJUvOGK573Xvvh0Mo5DZWd76NtuMkajNYIzgKp+c3yphASvAnb9yONUJq
piLrLSo/4eLoQly1/UB2bnJI3/SctCzvO9LkJaTp4H0xts/fcZwo72BWGXHv9DKVTgx0ltuobZYe
yoQ+TOCYMHBOp2FS1IHiHo8nyrft3hRO8m1YooYMnsuiDAayGfDjMBnJs0irA7Z0B05OZExtP672
GBohGeAdOU/3v0sEeOSG1ucGTO8yWpsMOzhUPmVdT3ffqvKPh/Cx8x4PzqFv9NDzRdv5lBh+7aVf
+IgFkgTP9paXoFfqDTn+sNxUCUzc4E+jeG23RANevxZ7UAiGUF3SB5Hwr1gveGxLlpBsK6Vn49XL
T/cMrzfq2BACGp7BiF8jGry7V14oF4PLZi/R7o1yhZOtfq0rzcoGpU5eVKSOAK/eJjsUHSopH/3R
UryjbTgdKd+GRmSNjiUb/lIM/wysMd+X7w5Um6bbwEJXM/sFUGUdma4t1L/bvgP0hUGLCpCHiBDq
R0SD9NYD3+6i7FYWBi0iMIjLazXtWJhkrIZZD53FPQhSbezBfZoFle75H0AYghLfS829KZqaMbyO
q1LsEAo6nECzBnbzSTvUkrls9LFLiik17oSyTomUUyZSli6+DaxoXc54o420+IElFUBYXEGcNfNH
WPFrNX0ksBV3wnJcVElkhXrOhkcMgVFV5i5G3nVUkg0V7krrZDtmAaorbmxBA/np3GgyhsNU4G01
szns1/H8cAYAlpUdhjmIPAYx+9xZOIR+sTCH+qAFlJdddb9cDjQFkIsQNR5AfptEtKSEam6vp1Rv
JUD9s/276ZQmDJjtXXnpBXnHTYbBltyqpc+hxe71JFxBqUqoqkHd7R3vbgrGbB4NoVoNky+1x1Rc
X9sK7gm2VLBXGUaknfcavqo79Pu+DrEGRwxiht/GEOUOfPhvBgRjfO0TDj8nmSmsRU90Kc60mSPj
dJWC7Xr2T8wo0rtlKwHPmOUFSY3bOr/VqbO8/De5SSQUX6nJyqEge9mAGQiamTY3pL7vNsEQCj7q
iknO6XYqwoFYwXqOegJTV1rsHge2WWZM65Pcf7VHqYve+NxpZVzse9LmZXN7o40guK8rTeJNUael
Dcyk5xHFMpkRWgQkCBANI8LYrebDr7ySbL5mr9fjDbEjlPlKLqpksXaR00qTeMibdIFvob7UyBzo
ql0R4YbcZnGPH4QRo4nJ+esgQZLxY3ayQUUwWwoljbeEfNCOt8Xy95Y0mlDZo/B8rTB5SDSKR1oK
IuQducga2Rx0cRylxBoNHBrBGgkUNYRSlLCgL3YkPzfBPelWTkxh4ypqALTgNEzgCM6atvQ8XGAs
TYSsPlKxIlFIhHm9aAJ0mg3AG08/hxo0qzm6FNt8p/h5XvR4RDX8gkE0Gh2Aq69IvmOMSbb897LL
49y54Ym828HzXmwKTMvbrM5w73k/Rao0mgJ/weZVvpZyib1gweTy8yK8jLnrw03W/hpbDyXZr2as
OPU4cJHoY5l1favdWbVO40T9ptVZbp8MXk5XyK75cIMlydnXIxD2WNNhoN4trIl0m0g9uFRJrqYO
m/jztiyPT2VLCc0VuBoPoCf55w/fdKGCfdqR4AN8zc1lYu166ode4wy4Kv1swg29/WpBKbN3fX+H
Qefj3fmE4veXTkQSNlQuoPurRKIj3VK83WX0/AWrey8sArFhiYCEI9Bxc8ONRnmPSw1+de9sq3sR
adnCaAu7wlEYw89/HVc6b3E6ZOl56ZIWz6CPXYBwccFsx6fAbuyhrKKscVWg0L6wMa/cR10LFNpB
50BYoclbDmnw1PnyTLqr9Ocu6t6dENvDCz1Drx0rvlMkyWal3ETbm/17ddIx95LNdkaV/OTog5cN
oMQ7+lcXm5tJqbL6vDNjLaV2kybQ11B0ILRp9Y7NXM9nT0isHfIfUa+vGLBiGnHg1229jgP/dMpG
y43ROL4edOLPod8L5JhVm7vz2khACesOzjiG/tioOoDlKg94yBBwHhtUoGNFi9W+XSR8dQW8g6D5
Px4vF3uo/i0viBOflB4Zq6UpydCE6Ju9+1dDu8bChED/kpp12FaKZnm7ztQ7B+x8k0LV7qrbpGgg
wB7S8HGX/9mKPwms5byj5Phll3Bv1bYF7lmr+kYWkovGaheqMAcYnDOpD3Me6p7SUgLzqkZ+nGS+
nt2J70eF/jC4U1ixu5KrCZJPeJMJffuAHhcGjEMKg8g0xHByszjBxMkI8UPbB5My5gTdoXHcDx6M
RcVG7t8yxhCNGBdq60tcqjgwPX4fc7Gshnr0MtJEmrkUpzx58G2VSIoeBroy7/uTLafT+p54e08T
Fp2CWGLgo3luHwt9QGmZqBofSNt1OHoJPVA+/1eue8DwHGgISljaCVfQhsOS/9HA1/hubp2MYHU3
jxm3+xq9c9oyY4FNpvCQw97/8LIoyw/reQEPj4IekaW/KPtIWmiiTyMnQK6++hRAEkLRY4oPmHUP
gFtSG1nOP0OKSLtJ48qIInfWRglvCL7WxImkw2U3aXUL7VFyFqKMx3vaAYa5KVXYQd8gAr6Ghrtq
A5kCmqudi5I/D4a1ZEQJIflvS+ACsu8e/qjMw32pij3m5zJsOT3A6sqSyd9CK054fOiPKw/yFet9
f/0Z8yj2gQ6zMwCgrODoEvvJgr8K7Ip4aU87RDVXcG8fVoeMvFlcx1hEkagb6g/vY7F9nYlF1mh4
t7F4DF7GDNX/atydLOq1B9TWLuK4VgmvHpFyylc8ZihezP4AEX/tftE/K7G/bkCdvdDTX1oGoR6o
YwJsR9+chxwGHC4oV2OwKMs7/zT5FqvhE0TNX8IhBPnTk7p1aZ11KzfUc15g0R3hmua8i2VXOpmh
YSnB/HKryW0k9772iGb6i107RTZ5BsyFDYARZdo9ygufSZGKwhu/Lpd0X/phFkKaz8ZmyQysMb9H
HQxdJ9JngiLoI8X7Q+JDBmwrnzuX2oYEYI41vef+OZaNEX7vT9dY5jrRZceAxH5GT0WbykjICGns
Xgjdz5q+MEE2Eux6LbRlZB5NlBdj+g9kkvt9K03kKRZ1Hr0Lb+PXftkEuGXAVS3RPcYWBhsKCVJZ
xGfDB3JfTcGPKE2Hd74O/l+Csrttrz0wRK1mpEtyhyX/qzedS2+5N78l7Xrr1j2m3qUEd5bopcnX
VVPlh3ag1qN2MbhtcJYneATzupF2xFT2pnVIl1ki6t29Q9JoEr5GxT/JNvz1QPc+wv+sB/bgGO3f
H5sJXaPdjYCrYxsbzVMr5FuvT6vxN6Ztx33yXQJSZN4bDE+UFqOtYSaRcPDYsAzwdjvbKE4Fzx5c
J1NPHQvf6ltprRv6uM2G+qzlQqHErm8rTjHpjZCFrJyWD9Mc3KYjh9EcWud/ulZ0zmxbH/hiAKGX
1rWegtupplfflFrSG2PndnAYbUodlHC9xjBqfGU52euHjcpN2VuenpMODe5pR8udZipSMWTuAhQm
vaqrDqVeg4zl/eDhlu3fvDsCT7VfIKHqCKNjVJxMpGGnb+8uOoDIpV1jLxZoqFU8nFeHlHhRiklA
JBnvgqng+xY6zvs/AQTWKn6uCsbSPub8AsuNE+QzymF3yd1aCfPnXXXoe0P7CBC2OGckiRckE74p
EjDcvIdVq4BUKw8Tocb00eFKT4nSJw3ofLDCI0xrBF+daqp9FTnkM3Q9Kb/1WFCqlu4pS1GNuBUp
EtTujb6/OPR8LhK6dUEIflzvNxX6COyAV05Lzjs4gkri5clT4oDDBwnFqWFMG55W1+oc/MePoHuV
m0wfjsmVfMxVpxDifGBqEzsFLCFRRpQ//s1YfjOu8svQrevAqpiygwNM2KSiJS0Ck4H4LiKH40JW
BQX9c1oblUzdkb526l1IwONI78iOwVEZ7KZJMOd55puV3ElnpJ/QzSe2PqgkAn0Rd9VYcXITP0aY
G3eVw7wWMUk5bKPu8I59Fh3aDmkrMdHEciVs50U7HQ0ngk0Ef5L2kNDsRSIPdrdIxQvxbF6W92MB
q4liNnLuVVBSYGlz4w07IC2E0a1oAwVmFEDUjMdHTziuLFlPvIdNLQ4+5/chplwJi2bjFwpAEf2M
8hxOgiWFGz3rcnJC2NvJRQARHJLln2q5z083NmRFUaVnvwTzR4f/Gm/95AFzdLFUvF45/iyTWCfO
mBY8hmoyhPBL7w0u1hskONGVcQiQcFZiUJV8GhcIDE8XQIPXvNkAsMrceEPpedjEyx3wICa/o4rp
Iatbx6q3+w7xPCF5qMNYbsR2SYFrOqm5/ISlnKGK6Ckh9gcnouk+F5PogM6zyJHNUTTETerq5jmm
eV0NASAkxwPu63RuX2xwKAv0hgjFvZNrTvrO1pjseWHajTcSRAvRy0SLmM3FHiCz2yX9YzE403fJ
MAzTf58BnOAGPnfnNGptJc68Lr847kHD+UEN/C8vBaUBn00XQZ9QH7FzVrReUo8tbQIPf0ALTMbB
HqwLgrLuZnl+z5/BN9nCYiEcVZgw2TbQPzqgFjO09uwy1RDgAy36eQR0KbBP2TSZuWSBjDVz/dik
hdti58qSiTX7yz8U3U0z75dgpl5cnXceqVz6RIafdL11QdA+XM0TCXCU/vZZTeUVAeNOPvGn1yo3
7agjD+oV+pdk/a+WHzRlrpPdELyzEbbTH8dmRWtUlRnVH3Q0uLBz0iqgZZvPYitZqSEbCxxK1jbY
hcuIz2QEwp9dfHwYSEpN2Y6pf3eR93/zDCUV4vb5T+a4PQE4STcuCWen8S1kiBF2b0mVEHhjqRcu
USm4AmnzF1hP1rO9I4SAUQLn9xOJxjKgZV6MU5VF8XUdIMXJY5k46XxT6o71ClQIe2Xxs01isrRh
cYaG1Jfgl+DYXbDAudac3KSIHlJJXI8mfZpcdqeJhLeePoB91Mnfq7k9m+t3EENiIRLP4yPRxHNK
NlY498EKvpaYF0yiyT6sDuyMuZAxEoVROh7Kqwu7olklGCuHw40+xks3Qa1RYYculjiNCLHKt9YX
ph3kDKWCz/TkdqbkhIGyZ72Cv/8dqsF1Z4VXCMgjOVdNxU4/rerf7isYH5dOXzb2WHeuKuzPNOl0
Afe9gUOXk3mIutwu977c7zAsjncEFIymfvf/WXF9+z2IdxK/cV+um56v1ReE83JVjllBxLTFXKPp
9ij/hulPqogP04cAi99XCkT8M9z8JU0pbRYLpSgG9vmV0YbT3h9hHo4341BDK+G/IHlUSckX86n7
lcY3f8mBgwdQ498+hRtdFY1BGipevR2A1bSNGpXdIVgSO2SICdkCMlRJo7XmCqoPfbi4wFlGtB2Y
BrAxj6tSGsfviqrfWKszi73e3QVxYPx0F/Pr9ENbioJ0MPKF9hyb+3IiICNDaSS6w3aulLqu74Sy
4U0if8aFuTdsT8et8/WjvetdWmYb6CHBIdDS6iTjoKWLB6IVvDc5mKIRpcWjbxs6Wzsb/auB8Pg3
mxM0ImdOv1MVS1O5EW3dk99iVPM9CcpUbuCobXvBc2BAyNnaqnlvkm7kgkW/A+JbuPVL5F1buqsT
w2+ZPdDfj1RQysrYU0RU8iBw54/1ogSPZO7Vr+V26y/pDBjhCL+hAR24DWGqf2kc/Omf+ypqLQgg
ZrVC73Bq1etYbirUiHaZ6WPW5G20m41sCxX7c9q0dbTSY+xqscE9SuziW8PcRQq07AkqR4qg3wii
03jI4Z3DX8OfHun/MF2vfwlz2lR/AAgyl9pRfR1qfAiCne/yxla0rsS2CPbhY6iuj4kdr7Ymfww5
0VTYNZdHFObUS1WImnJaAl4pq3RcuPmSxwzUuSmrzcsEasve/9vhVyYCZifIxk96MPjf9gOg7gpC
5H49qJtw10OFwKg+IUEnn9UQOwqoP0Uw7qu8VW1U2SR8Excx/2dQ/hwlEwU8fFSk+pTE1aL7BwuA
P1XRUpZH1XCTMe+if2rdKoB9LEi9Tcb4l6COEOcj+ePYDNyT4CCjddx/HjadHEv0C7lfpCGMSIBQ
8un/n0VRezZdgD7Ihwl+jBUB0fEb2B2eFIyZ8woEg2DJ7qtr3472agaEY5YklPyAIxn9moAP3zuo
cvj00S8fokPP04RMO6Ofy/iDexMhYqyREPpH2VxieP4IvCvKb/9V1zfC5hPRKCCHRhaykjIYYsRU
zbl5gtsIiIodur/Kf3L0h/pJBB0HsedsYpUxjQ54enE9xwXTzS7UpiKtGPFhBM973UmASJ9aAxOc
vMVG5VhW+w6xK705/S1all80oMcdzf+caZLz6crY3H8s/786IswoqSbnV2is9uFZVqkBMganA6qe
A/nF4Az2XlqSpLQkRPjCuOQmUcvWpThayKmyAQdvfrb0l4k/cnx7cpA9RBnQFiBvrYPD3zeOFxnv
P7OHDJQDRpcQEZbNWdhCu9nOEESCQ0g7dGWZKEeOnnOOjcl96/17kgptwwHYTModxQV6BE2oBsyE
VUwoO4EIUTK/aAJ3sRIrgUCeuonFYlNOD88/EjvQDvPzuxMBsSDW66auTvgtM4R5xtedESropyHx
C9C2wp3EV0cSgwarLHMUxDxIYw18PcGaQfCcVr7uzDmKYm8a64H3LwLBaH+MZQ5ORbvbzW8QQNJY
L+P2mWkPQW8g12O4/ANbxF+kqkPzhJ+vNonBd6aHP65MuDzlWUZoKwDcVDoCHmIg64okGyGjGngF
Rq2iOAiJ2s0ymxBL4JPyS57lmPH7bxaGx6UBVHThRuRaNaXz1gAalz/vHgW7l9ANYy1S3SrlDj0g
RC8gmipvix2X+crGangUKxzuvIorCXpNqlAge5nlO8HwiblidfD+jOv7Oq+bVEtl3zCwZa/RlMOL
nTCCrapH9WDzTrUvdoo5qzO7LJnxd7Q+aQr1k5XrWFLD1Hecl+8ZbOuWAiewgp2CupUkWroY44LK
9B1P3hvSvuqpNoLXQ+jL8Giqs/SkZpVGAm9xE8mLCjE2fyIwfZlcf+R2ML3qc57aMdijfWxN53wE
lM9ZzYxS+8oUJyvevpmUjZiQCp7D0vPqsPKUg+bLfHjVeymYQHbP018/iw1ynB/bMa/fAFxrmCvA
UV5Ju0YrisWV0FixpZUHimnVu8XyzjcAF6/uUWsYw6AsRpe9149DtyuuhAI3y1Bgk1U+GQ/SB6Eb
kRpq6SSLbVoMxYgDvpoG0Vq4NpJQYzjlgcTolp18FZuZvj3s7buX9YupfG40UKi1ttzOfjI7wiSe
9jLPpcqSgXdyamDvWTmG9FCsKHSc7lhic23wLB+1a9YU6U+6YG8G5AvMr3j2fXYNigjBGsHhk8EB
zH3mh+EiGVtxwal4sv+KTCNIZekpHx8a95nivgeeeuQ2S/0ljIn6i1rIfoWtqgs30Z7So2AypOBl
NX11ABY4jYkIPpWrekiEZMDRKVGD+VjJ9m2E3oX+OjsNanDwREBMsn+35OIL4MCCTFrEGgXcZyWK
FmaItE07r5NquAjtQtaFNRdLa1kxQ/iDaotnVk8UOqpesD2TogUjapvbYAWJJifXur5WoIhRjFrh
j+ZjZAih1p6rq5S3RQNQeCq+LT4jIqXFdtfe3dz6ivyBI3VZlK6yxljrOAncRMcyY3OxQgwami+k
80WKCVLzZSJXy92ZQPDiDx1Qd9G9Fvln3EyZrh0lHfaIivinTkkszNvg9sZnjV8JRNJyhkfsi6PT
SYS5r1v9ygVW8ecznsHEr7MvrX46RwZH9ytNG6+sGZvAOIclsXPDcFOH0UnnliEVpDox/gXw6Mg0
oqNVL38jENgpy1YyCcaQt8ABOq5bVFkDNP0iIn0bbIoxf+Z1SuErsKwGkvCutRVJg5pxXbss/ft6
KLoUFIPyzzAIng2pgz91Kfj5OK0jo4rJRTcMr1Sy70UAvVFs3wUU+ZfKXwcCcDXy5M/T2vsmQgVR
E+ql8MuPR7gALjvX22NZpxfELhBXUhLQm4THf2iM5KQY+DjlHqwYrc83l5s3CJXjYserSOwn53jz
sa0fGse+01EoRO4Fk4q7vRhqPZoUZTlbhLW8z3hSQsCx5/puDI/xazkjfZHKQa529UFcdqeJjQ7/
J8D/Tkq/ArsfNkqWOS7gVR3dKNo9C55V/GeZ7hTPiEz7O99RNMsOuRva8aMamcLKiCqiHWHw897Q
YmynyuJa5LxoUl2i00j3WX6qW04RnvEnxQI5n4Xhuc4LVf3bhhV8llZVQhlj+hlxyXUU1JhiYKMa
neQYp+OcopkGCnXuOfrqIK/b/Sc7kvQI3HyCY54OmVIqn3EimAJpi5Jc0w3JMVG2S6vLvKED56oG
utCOzMVqxyqASuXfkNo06bNCXCOb6U8d6AIALZ/jYRuH5ZHOAwwblCVfZsDFoda0OXzqTizwmGSX
xY8pLXWzb0YC0pbByaHlopREUZ8AbbY+JHrXGMI10Ct26NgkpZ75vsigMjgHEfHyPHq1EpTBT2zm
qSeSoGSTcVkxCuRG7pHTf3vCclhF2I1gpuKnMHD9aLC4d3jyM9QDwah/9TwbjmADTQ9QPnBZTOeO
QBXz4+2SJXQ3xtTDgKIpwiTqck3EgngVqaut5/0D1UC/jBuU2JsIIjaWcmV7bmvD4Yo4w5EETBR7
x7oo40eKU5iN0P5ygW4LVkusF3pUAdk+E9PygLwnjHoQqKf6L1bQivbDjbfmMuPiZp8zvqvrmDuF
UUB0TB5EFLHQGC0zUsKLQR7cQfTOucOROpysnXfKQr6OWZXS45CuTxRitxj5l2/4SAMlgU8FqS4N
LKfvwghdTNq3Pu24+pwXhhF+Eoz7R2XAlPJgWo+Ip5++nGFa6gryClYx36RBbXpbA/KEmtQvTz0g
r8WWnfl9UWVeXzLrxubgqRdCPOoliOIDqKDQ9Nu1GTCTUjUuaEjL3YT/GUBDDwxXxZHvc/hRfD+n
FOMo+xYlYEvWy6/SPHoyg5XpIat0OY5sA2JUCyN+kcJrOERb/8jETz0TbAAF6QddQ5vLffV1lDHj
GP89w08+e0mCCy1NUhNuOn/120fSj3v4FYIk5gb/7ID1TvludOXWsJ5wqoLancDt+aerofUzj0Uq
EKedK6ZCYzVcScMO8QsYSmLgiHOcRwLZ8sEKKDEgfb9vl5/OoKBTaLtHAhCBoFIe4zmMcpaLnlrK
/f8TrpY8jRCRwriRMkDEtdwVgHPhizy02CEl3tETj9YQVDaB2YlhFDSFgEECnEf2lmJcfYdrmDnX
FMmY+4SBknLxjLy39TjT/7TTQoz4KaJxikYkfAds8TQ21uKNYBUq08R+BMpVKOnxhX5tbCv1dKUY
U9tYabmSiDZnZ0o6vf3D2jV20iGMe1HCT99z/uy4by9i9Axc3OM5aGX+27x3RO1ggCFgvn5TPUja
yr4nU4k408T6vdeG0ABHd+V9zqu2r+aCznDYMqSI4QYu5rT2Wv7NbwocCgfSmusdTlnZVdwPEIMU
Pa1XmVy0yD+y4QpXzpVfVW544sK9fnxqshaBeeLvbeahSq3DQIW97ybtoI0Bd2g7qmGPTa7n3Vv4
PkL03g6w/7EiU+1NmLZ6PyT6yWvEZ7DygAHZg469l3e1l72Pt+clOjbdVMwniiyKVfqTo6v9iAna
WsVGtuTFKqMdIFM1WDJFG4AiT2GTEg0wYjObWos+VWUJVcngCPKNKLQx/rzJKa2hYvkv82uw1uXn
5nmm9NEbN6n44GHFdMdHL/knug5tUB9oaY2hI5tVkH2ntg8Ou4g+WoTM6yZlZb2d9m+gHH6u8JsJ
11+/+QbOILk/s1aectjSztb86zGiqtc3EIAH0hos7r0rySuAtfhdozaTWZDiLYxpYwARNsefl14R
ZHK5mxrx7W0H5Bh2VOJAZCr8YaFmLUgBkUhODVNnL6YuhdxPV7iT+D2MzYi2i4P1o/P8aB6xRKOu
2muH0XQqvLJR7RjHCAvXOodjCxF6+RKbzrvqyXdPldfOg4TzmCilOPVd5wu8Ax2Gzqago+NDcGOE
YuByHIapJHqK+h9vwcdITwWK1RwxvF4fbK62oCnmH6GTaH28iFDkiWLURDsE1ywUQcb4rnCIhShi
8QxVxpMV28xvzd7Eg4TZ7QxBgwA71uE8Z39Zo0+rTk9rdzlYd+Ct1o9Lqjwr2YEJ6axZHoNx67ln
ZmmSePzUJKoPMBMXtUYdRzlxY2HVoqzHu6NSzOBOdbnumJ2C0irGyHfqIajgCM58+1kzSNw3wgtC
Uk+u6EzvHUpFGhzlA4ExbwOosCZl9p4/QXoJkNfAf4CTo1b5TynO1qa+WB4jCPT8diCI21BUC0eV
4+mK2AIQYZo9Kll/squEoUvm58pKn0i3VP1JY9iO8HitbBG0Cy7qTb8bTTB4C89CGYzbF2w0m7vn
rfBpbkzCposhB/q+9Oprma7wmBrKFqPGOnVKcWivK2M6utnzEocDt5yx9aIIx3grz8m7i2Ju2ZaT
5Kp86EK5QH0it05JDCXkN6muOoT/itPu7WnN/U7UusuloT0mGKVHFAY7KytBslNLowDj1u/xG7hF
7ojox5V98WGDx+/2ArU2iJZt1xYSzDUo4ahGjlZrGPQHQGWxaJDTgx5r4ODE4D0fYIIbZ5iIgvaC
sh2EGlRhP6FojndBiRYgJgUjU7drTdqn39bzJxwkm3psBUDZe1HENtHq0ED7/eiSwnV5NjRshqOi
7197ezI4VLvq+9f/oljKVlS7PlTYLa8R0GQXO99HIdD/BC6NdqxinYq7fdpCO8SyA3uLXDfrhHzt
uLMh0ChIZWRNFZnPeXW5czljVtxg6C9JQX+8X63mTihdVRoUmcLjs0fgrjZ2YKm6XXpnnUFdLcOJ
1WeO1EqYABUM3OvFN/MU/347S5uuBU9q80UN6iY4+b2ht9sAN5xzlhpl9x/ayUpgFr9WZSdORR3P
PrGA4dr3ggjMNPuM9qgMgOSCZhbcPDD+ZDzYd4wr/Gwpnh5BZ8p2qIhvs9qkIkdYp7crf8Tp3L4E
faWHHHZz2hIEMv6cekCOGQdetDTu4O2HbrXjfUKNq9JgCPGmd1PhEZdTELDHJOxEkBaaS9fxIlum
Bw9DyJlx1RiSO3M0lhFlVRrmUCzEKb51JFjGCdASIhAEpncx5BQo/fX3S8vfxCq+LAjympaw09Ge
9MHBQWe1DtCi5VGoUKFvOnkILneQfhxVzyXmyt28Sw6cOAKWlL0dVii780+dGwXmMoOkCM8hTjfZ
2ky2jiHncj0k99uieOsuMQi8uEE5KIi64460eGScEodLqdnTAOprC7i7KBFr+QeHlQu6zmD+rU0L
S2ElEqKwq8lvFsngTDbaNSNNtD1jd2kUjEmZlvuHbFI/LIjaVkG9URxn3Sq2vZmtq9KiyyO90NDe
8PKAJK7fwXGPI/npWylOrmXhgmTVtjedP+m5f2+bXuR/u02aDEepyLltHJgssrkCjjvWiK4y4UDD
5mxigDNW8GllfDlY1kV9yytkVL510I5F3LQ3Cue+cNtUJV+FRswyzYqOeffLS1LYEjaJDT8nu0PB
j+92dRT5OazuOfdIl1dBaejKxrWAQqaX0atpLAvOsHU3DXxgRhakXP/5kQ7U1obY3RaQu7U15Y7w
Rc1/vkuC4Sn7fR2TRYiyoW6IWfmYEnjatNgI+QUhHTeDQFMe51qTw8LzwV8U3Ms2wvCssCzcbArx
RSmI67H+7tF+vo+9evue/XYDv6IMS4tRVMJFu14mS6GVrRVe5OMkCC5zRCFFUWfifi0T71wz6icq
/exKRgN5EvkTry19XxsqYSHQbrx0tGrKRcfq9xhGr1QD2mqOLHNlY/opHxwMe+BAVGegOuoS2Pv0
sVQlKa2hyzsO2xWwDmZYN4jlgtAVGKg8eTY99KxjJ2O85hzUetsXBOSTLUzRfM8Qv7bui9gzyKI1
ZGmGEvMyOQH8qEU57RhgovKUCDzfmL/6J8mwypQOJXHXKLvelvBqKZbwccWUJfKsUqG5WErZ4UMq
PP8rnBxhFbpImWqx6UgFLUGwofDk+RkWZITdZ1C7K9jdun2hSWWfRwsy3wulQoLDnR0qxvw7+kq8
9zYR6hBlkgh1Z0SH5yDZ/mqqpr+w+knc2YyKePLE0fd3gZ3kknNHor7ORUewNfiG4iaoopvsVM2b
B9AY1fduayn1DhJ6EHOEz26NwcGDV/7/r33nSr/bzrKYo6XeFuB72d/CdQHlteo9ZVSCUyaeLIle
SufxWM0I6I74C9W9iuj3ipxsbrfukdWqB9zdY9KHfaVwCKigbxv/J4JRtmzhHj5f14zF0NsN6U94
PJIh1PbGfcX98vNkmdEsnyc1sUQi0n4VmhOIosnLh07uwRK+6RZLI7zDZdk/MTawYIP0Bh/yGU9G
GgVQKBjqX2w5dCvSiHZgAi1MtPux5HQbvFrpwW+m2x55tT0o8zJvyDQW75X/mjQ001S1dU7NUgtP
GBmr2A==
`protect end_protected
