`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qPo8qL/f4g8LOg3EtY31UwQGDRT6n5TVPPu0FjK0LpPPBFGSpYGPCVdE5KqOxmom/fSMaJK7szRt
Xx8ZuJiVVA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OXZ7EhrD3YXL0kEPJmQUhZlZhyAq4Af6/CMfGUDlMd0+WUy4CsD7XKVlEqLkH4m3Y9178ZVjItB+
n3xj4KORlh2mrX+KELVyVBvxGnb067jUjWNbMhFylmJ0MJ8j6amTkBlYvxt/tpkeg00kHygi41CX
RupkJaRAzFjcshT2yN0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W5drNjD16nA41IxVYCuTJUBmS4kKdd8rhWJT0cwhwMBwLE9Cq7seIXZcy7J4pCx3FBIcJkNlR6a6
leEKvYjFlKses0jbstUP8IOlzKcWN60fWqTysMNVI76izq2a7K6zNN1u2OQCGVnR3x3KJTa2H/tJ
h54G4m9eF+krk2rvtTi/xUIXbh4SgL/js92NIb5eMdctDwsf7/J+SUPO1cLzspQGoQvffKMClII5
B6aBwweOOZ3JN2Wmo9CpCC7LtenzZzd9fV7AWnlmHYlwzFRYNy7Q+VlWbghCdOw6LPV/IZob3O1M
L1L5T9bwUGTPla9djXX8DqMwUg1BVCe1bHYvrA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y1eyina0bo30zn23sq33AuWer82G7ckVf7C5hxQDTWOomv0VNEybhXnmUNuXYh7pzJ7W63u6mKZN
CKdPwmLTU1SiMXLrWXddvO9i8Z9oBcoel0NqI//eRpqqI5k8ORqsAvMQQPgVeCXiD7+vylH7vVOs
rY5c1WrEheVSyEY62Zg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tRj5rUYExVehnlsn6/y6040pKid0ym6A4AmtIxqT1C5TCY5Oy6+QD1++BM0jaDMUC/FJYzBLeYiH
xc+QVg5ZBsMEJk6yfiaNF8XnpPZsHovVabbrZdiA05UxGr5xWk2huFzsBKcmyhzYaww3s26UflPn
6I3l9IFLuvFtONOoUPMBRkHiD33dAw9byqwfunzXrR45w71W7vGMBHABC6dxmXiyNfDEkYwYAxHD
moUGRY2c9R/ZOYzN3o9c86CvhKIFK7UwvWZ6eO5uPC/3NNpVToEpzIyikJ/UysrxY73xEm6NvWoP
BD1Fc2gjSaau0X5E982gRSIAjgNxQ9Stz1q8jQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4928)
`protect data_block
CC0JpmmSQiO+xKZ+N93j9ql/R9QJV3bNLTBhDiJzp1DTj9cYW7gT9UlXZLblmWzlFOLp5dtVx094
+bLlStKa3C+PZfvC0kdDrQA7yAHCQFCX6lKsddiUiEixOwyCvqK9Ow/FoehVKs13z/CFe3sUMiwU
66NGwHUqXFVJs5OEArwKVFCNtXdH3sMQdmxG1nODo/0UPCucAKjR5fgeH/WU0R3D6D+kx/zsfU9m
8vCgNHF8OcYXBKWvdCDjJtttu84yTVb3b2Eb5OShlIISXUm59I4kyYEyjypJvMkMD4cohXC4vlR3
3of8lO6t++9Lg9ZM2q9l5Au/4UCZYN0dWJruA3IkZpYdMTfZAaCyLKgUP/CIQCt21GuWv4VPwRR8
mWbT++oWJPtbciRHvWHHxK/Q7N7RF+fkNcjfLNxfurxaMb2iGQCVMOlBVmV32OVxG+pFiRSWcdKE
bG0NngPGvwmV+FLBq2r1k81GODd1n/4l8kL+/rgSjnOQ7O6F233CdsL+MLSctEI+eR37WbUQSmtT
fJmDsciv699BMhS2UcEghYRfizfjTchKZth7NNqU8zID4bzHVBP+BliF75wF+yioqMg32hvfgiMP
JlQCEK4uZbkcS6q88eVfNDAZbwPseIoTNioVaFU7hX7fbzoKfb0VgBp7viLy53yxxe4HBEULxTiQ
6bGIYW7R6lhay61P1cbabvKmBimL+nxdUakp/fgH4At7iWyFiPE6050bZI9muS8ZheL2+qiLxAtq
SlxvwDZEeXBuVNO22PMYEB2+Q+UKr18HttyPB40ua5sF/4jUvJjQkZ9IO4lCrMs0gNPaH4EBAP6O
DqJdgN8XxhsKCKp7URzKjacFF7alPJun/ot5zgecJPHhJgdG1wRSdt1NqLjSMfz8vGpiynwENk69
vepYzMPVPfSDk+9555fqKqtSFBfmDRl80FIsBywqLr8KEI+LrGY2BLJdOqtvHeUZuNrqxpf4tIjT
YhwAqD4i5O6u5PCtJ1R3SpgNzq2CvMgdJwYqFNNUZktRvzjg6cGHHPfUtiqnn52xOthwXuVDRBPt
WnRzva4SeTXlQGeEJc7OSRq2IOgvdNr6CcizcalzaDXXcY4WZG5lNAesoAh92ErZ+a0feL2Ghqmf
t/3CeVMxeR/kffcOYIzREkXxrkrFKdXiML4JplwvNT8RnlcAla0md/AQEoyOJLoqgb1cw6cNU1Hj
4EBGpLXkNUkEoGHalccHNiY1deKJn5ds0cKVBVOG+p9tkatMkbEFeSTTx8+Sf8HS8HCswfI2IuuU
LycY4FUmA4vsmB/Sr8eF76nV/NoIYfAS8k6NTq/mIV71Q7HtvSzkpJ4GG6Gp0TtP/aGdwkgoVo1N
Gm05PxJsHYzVD8Q54ZzBAzuOvEIJFYWVaTKMBuD6QGUFPN2j4gIqgvEfJTOl6V+jQ4jLNeb/jr8f
tkQO51KUpoiz1UgGThc2gKJAc+sKUa7xlP8RLD+T9c9N9FWwZS+1HRSRzi7ZdFAB+zRJVMLge12y
mKlbRY1SrwcB+nemN+PBwLc0GbJSKL48TLjf2z2r0zl8gUBHrtWtdfFjjTbwIitAeFpXv7yLYTX8
mk4VwpVYQdxP0LuaTl9pfrFcsWzKiauWh43LgYqsGp912a9IqBhow0g3haR4zAkaNIKgNGH5MG6Y
uQODA1vMYMCPcjWLtmIY6JIAJ5RGJXau0XNNJsAN7KSMWGaVsYaLS4GxjW4S7RWdUM6omDyMjfYA
tBDt0OZwYQ4YXZI+3WTarkgppkl2zF9uMAxTVs3CWDvlqbookwdq5X1WfmkPqVVlBf7psOt6lo1R
FnFsKUUPWol/V0dz0bmqGqYjcCBehluUdllrtnsrBCMyXX04ag82OTv25pCZY7CXuGgz3XytQkHt
0naUu5owS2ZHiqRJWRokVx+0tKOIMFCt+UAdK9HJt7BArkYYYzb2hKrYIoh6L07pQoy52HmvYXYB
r5iurzzDXDpOpPCdA/uCfa7p9CTbIynzkNfkYTNSgetm6ICROmUj9V/y2X9Wo1wQ51r6DbooYhRJ
iWxVCuks/osj6LYT7X4iVKYSl9Py09BQtVfwRzm/r8K/yzjIah9uQb8YGOuierrpdpq/pCxasc4U
WUr7nlGYxRcLLCJa9uW1ujdwd+wJJcjE2/LpJ+4+OFQO+8HSEvfBAcsQCJTDLiSHKOcSmowzJ8Ug
NeD9mFNSe4tPUqoUj5J5Zr2DiDBor99UnfU1haJ8cMi0kR+SZi68u++KfM+RiaeK052Ac3hX/KWo
SpDb3IwnQUInI9PbiZsG/FcBS+HSqeGQo78idTeVuplg11sReWqTIxU4SZVxfSojWVicHikX/C2H
6OBiyBvShpoirH8Je+Wo2GGKM5/+XWuhOc8LUIgJ+DU/V4Cn/7jwGW+FzoQcjYb3VxfDxsYHx6b8
m7h3nhU8pHVn76M9e8JnC0klqZnVniuM0Y4CLMR8uZgwU4hIJ+8mSFPbeQBqXgBrzaVMi8FcPHtl
genPbhu4ijlJm0pjvKlXB3DDcgm0O5cNGLG5P5J2xQbRqTYUT4zxF1v8BmmrSnL8tVjusduNnckd
5tmKiCum0W5kdA2IQI8Y086F2Xiwo+6aoFPwwatMcB5MUgIR5rA9dsXcdB6NlUKq/PziPJVu+AYt
PZEO298GiuBGZ/GwrvHj3O/F0ckO5zDSxVQ7Lrozr9AFUoaB2yOvtWlIxZkb/ZOoECmzQE7lRAJt
hIh4iNbuTlXpCQOjNyEKi9sNXWkQ3EZ5tmqHz9j9k9yIJ3bMTcTHjPL6+2jcbSiAZe4U11B8Vgh1
RTT2fgsUAkbh8ffOXFOsMjexJPEh6f6pFFEJqBXNLxYK1DmQnKTTx6S+yOOR7AX+jKJ5rWNl3I6o
w7lWdmXPCAephkkXNfmI0zBLeQeE4CfkrszPJiySzwYX45d+b2XLMNa/QSVcBStJwtQtf3B03jV7
ZpHF6zLB/OqkPbQN3cjaDLUg2j7k76lMvU1QRmAcUh9jM0Av+FHfcz9c+zuUoo3aNCFZXIgeOXUO
KRa10aybXq8tSq1Nmo+1HKDG2JIW4VQHbwIzOqz6zY8cHOStlF/qxFd4QCHFVQAKLXq6tiukQGsY
gw/wNaEbOwiOMH8i8POZtwnOCTX4GxYhI0fshBqnHHK8zr9NkPmtJ6IfyvAxP5YaLfXlXUOaCjok
r3Maw76a4ftAvtTr+Cu/eXJhXn3VFxLU21cJf8zkhh5C25z0BvDsljFnvmBEnf5WC+SjpWuvtvMQ
GCf2nnQEoSeLgelS/qexJjwpeYwt+MPhhsHe7EJ5C0Klwvx48k8xBnfpZvv/NAs1gX/KRXEKq6ug
zOe2uJjN4u7k/rXUxNepKIHMX91AcmWrGkhLzbABOrsj7EOouDEKDw6WLjX8Y0Mnrg+wSf91+zpI
Nk0C0PYsDql3yf1f0fldmuGH7/GnqVtamoqGYklZdTv5haRvTQAFpEaytyhdRWihBtwwGE63esQx
cHgyFt9F0nmVT+k9BKxpZY4uRxt9NdlrG1HoXb/wG3JSnF1+2OcU9qCOo29cb1PYbMSLRWe/UJG0
gB6nSTRffdOHc9Wrcd2ZVSuSiXx5hzxicHm8NnO2gf17BhV2qOOm9DgrpHFZpqXMUQTHNFtzQU4t
p5GgCuKqXpGtn3Yg0WSZImNPMWMxUYKRVQ9CxTgyG+GU0KK3VMDYdC+clOedWtHv6GyjwGrR++aE
di7y+cnFrOoF5JfB2b4a+sq/k9lZQj+3wpJWVboH8632lDFRGQbUGeFiH8MLOY2BkmKDkpb3aoUh
a5cOSeY3mClsM5nPPdIK7joSpDbYt2kuKRMNbU/7TLtprscf7XjGizVuo3uT9t6flCr/sSAOPuiS
+CxFTrdqabKErCBPQ2mxEjRwEjEB1rSnwu/uNLqbaBC1KPFNeG0aeM1+F0KsvNvzTP9Qc5UiZYSV
L0n4CL5Z4rTLVOdVBFI8a1jGeNEqsgbiCLEMwqRB43jIHfQehMcklXxXyYk5qgxSr5TpOkcDf2QR
Pdv0v2H2GozHvuTbKBOzu5DTRPM8ITQiaQGBs3yMa2b+X966UQRsWoCvsC57qLtqqB5ueVlp2uX+
KnH9t/ccL6i/gYc+f7X7LM30OkTv7DjQSlL5++BGPVHyKmjJEowwBZdNaMH/CrpV6Ecq1gmt/7yz
rKoh4T1nfuAba073v4lQzHqY/At1Dm6u7X7rRVYsgeiUoIbU9BrvKWBcDn+fnHN8PzUikAW/IXjb
2AXViaA9v/v74KQVG5hpXT7arDbWr29A1sxj9fPjmssUo1UFt2MVF7YfkQG+oZQ4IEKCzNCOOFZ6
oaOuembJruXf/4aOid2zoJQeuDr3E3kJbho+NngR0e3Dftq0j1weRlYpTWYp3NwhF2fVayeJ5pbc
aqyySUqLtHqKjIMV924vNlvVBXFY9yvYozq0G6Wx++BU9ZDbsSlpV7eSjt+pRLVH7w4vu91G0ffi
25jW5EEUgSrFZi6ukyro2ycxediL1vwJTTyOrdtgiROqAdHDhcY2HPt9LoXBV8O9b57mfH5u8D0K
NQYlzBjgAuM635W6rCF8ghvku9wlXKGizTrWrbpImHUtCWOVdcBRzKfd3RQOPc73rkDvV57J1Cgl
maUYswPQsP2leSeBcM342O0DCzQCrx03mKpgUohs0lsSkcgpcipcb6HBttiAZ/vU36fWmQw74FLo
89MlIpvz7wMZOQ4DvheheboCe34xEPPQk4k9/Y+KadxDHgp+ESLEQlgtXGNCQjaf1exh556cYSv7
6jj05z4SYwfPI+b2jDxXo5Kt4XhhBvldPvDig9wRWSpSJePWg0UxCOWHW5HEjhO6uMMdbZDVJ+Vn
q0m3P3RVUy3JjubPyRBX8/Q4NtGmhsLxTcEvJILr9blvNcwaDbQxVJNviNdwHUT19UGz1z8yTRGr
vBAVHI6Qj3xvJEaFhtEFG+pZMhMkFOdwGhXQae8vxG2fZM4W3/Nvfy6NgeG6HIFmpdmqAI5ezZ9B
Tq4O1+sbc5HfgAe7Io4UU/B9Xk49wFQ66d/JbRQfB6W3oXA4dKQwg79u01PmbmGpJbCkTieNH5Hm
g1eHhjEe9sK8MEKLXB5xH0SCjhSRPcknpKFDVSC/WM5c0ei++jGPj3wzErAqd6t4iKsge20vGKme
Lv5Mxu38i+R1y2a288Luiez0Vp1+YnUyI2nYUXiH/BxD1LfNPfZimN1nqePJ8GlUuHHcc8XSeTz0
/PKMwSuiYymcy4UTFwI1rreF86vdDl8lSoSnlHxQST8qFsTs+Xj6OFg5LnQOyPcGXs4x4o7o5hvd
ODdYRMSeQabFFvUHNlomXacGtHf2i2gx008VzUp7qMg+X/TOqoOTilnMg2gEhUorciVV+lF8PjoI
O6NmEPIXfcA9SwWBbY5HGCKRP5Cf2bLd8tw4NeplZQvV35Or5MQZzLFC4ka+cAOPJNJHcdcmo5gJ
XSqOCavLseYf/fy6+dZX/Pbpl1KTuytIFKKWhWlnuEnS8udy2vcd7vJLxS35ePbggA40et6eqSSV
+EcKVSC2NsaRc7reDtcnFDaJ4Yg/LRRTbMO/DayBU4g9LrLtZfYcIrl1Sxoha8QMC4taTlkLHjfg
I/IN1ggHJc+lT/OA8KdXVYVNdbNKtmb5r3LldA7w7T3CPSGSsfN/RDUHdYK6kE02bnRa4QA00NCq
ufKzgOl35h4xq6D9FK+0+xJomxxoDg0Jn7xzu5WUpF3YMy8aUVvthpSBHGArGtHl4BmiIbTrx+bl
+OAOIpg/JUQMLx0Wl0yhAu8L7x9RGMjtWLAFQHyc0xBl0kCWmJrWPdk9fwe78kXeBjEE5qCwF24K
tWviqyIsQe66i4S5+K5jmKxjTKtA9hOyKKKNaogkl4tcnKv6DD/jSp4bmyAaPJz1d9S7O6R66LOY
Lzh45D39FXhb1ZTZF6BE3p3bV2+CawNWexMStsvqvZpbS4xaIUztzM9DyjyerzoiJHV3ijnY8s3p
fzuvebFc0YIpvK/kKkmEhNBe6aM2aChYf2cWTJQzJspT2yM7USQ4/7OzXexo1ce08UcCK7S0L8Xk
JQVIy//AMcsu4Yilt2UkhZgDYCA/KX64qtvdm/4VEmCQj62VjsDNWZIQg5Kl2so/KJuxg3tx/nxl
IuPNuWNrRIW5O/oCOXOHzT8zBTcxCMDrAaGAro2kQeHHlqpc7xBOdEkBCP9pn5zzppiZW2EdOQSY
/v1iwKAVunutym6KLBChf0DiabrnBuK2ZvzO436vHYQdLK37cVVIFYq926trGhrO1IRpPC3A869R
WUNDWvJ7nM6JhOPnGYNES1DszfA+vr4dFrpPSvhzyC8fbPBFXYMEwg25G90M3IuBiMqhjwvNFYA0
DZ3N5T6nkL+RzEgeO1o2yrOhGSqL1kfL7Zi+oXAen/HF46PPCJPnpC+oRimfz348ul2wYnS2YMsS
p280ClRFacGfwbvd9WHZgSsgxwYQisAQjj67rI5+mrhyyb9uYhthEFseM0JcCKb32kVrT3dihRXi
Wc1WTKZ8O2LXo20H0A5IyUvxPckqcbmMnuI=
`protect end_protected
