`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cGPwkHZDa5qef2uO5yzMDNHGcsIYvJuyMQRQH8e6Dk393WaSD1RhwPo89DB/QkIJLQJdgT1qSS4i
nAWNm0zJKg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TlTxZqy28617ZhJp7COpwklvzwTTlthx/X6JCUn+eY432i+gm8b5fbusZ1jLeXhns3G2NYBWs7/G
izghSFFv/5AdTS3uZE2OzbAr9O7GmMixUfqiIB8WobwsUdpVarkyjtIzMx9B/NIViR2En6WkkLvR
b0jQbDFCf5dUgeJec2c=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
A8UaAtwt5XgQxdxL4BEWIi5csqIoSo/hVV0xq0tkLYaTvH/0zoIQo6WvX5yIko9RmsPg8mU6WN+w
ZABJbIdu5mf1Pb6wYgmeMCjxz757LI5DZfvCsbsiWxosG7XHsKw6iC6psbep8F8jIHtop4rTTRot
rk1Z3EWWBY2wJEX/l8cyUstG8SH4HGPC1Df31/sLRxeeZctca3p23BbC8GQ4QAb2XabwniisZlL+
mdWCqaoNyspEzT7IiOCJl4q/CaE+YdCOKz1UaOf4p3C++yReEp8Braexs79NJrWooG1FAT+7+qZj
v71Map0fZ5lEbOoCU1s7JZwqOngeurOXUNmiPg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QBQeN/IV6OAhV7DA5yLCkkwuiM3/lJfeH9S/vwfk5gtjKVLDFhZoR/qMwvqD7K8BaFvQvrWacR0F
rfqKYiCI9OlJQoD3yMhqdBjM14AZUZVz5ZwVnFVo+ddpUHRZbmqmJGbQPgYOoBlnYjLpaPlZAGUn
mZa/CB4eEE+9YtbBK7U=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Pnh37oICzWtm5R/oPDq6JoUuMaH1cNh5gCbiJ0BCpskwYvvsgI/j4r39E0AMstJIn5IPYxL6hLtZ
676C/wGbMcp4Xgo4aiV0Ceml3KOBY476O/v4EZly6wSo9TjAmInMSv91IWTkj+RgIu1keeiHiJol
SI4vpfa0QU7H+AbWGwp+7vP32hTh7u8kLly6edsRWBS9DGa/SDVVoD2rsLex4ZQa74pZSx9qS7BW
N5AwGMEd5Zm6xFPPio2v+V/uQZr8ayC4UBziNQOCHjd5sSCuefc6pnzvmc3ShhbGRi3eKnypShI+
owDcF6g8ABs08DCX2JXdBp2xWNLl+BV4MhRHcw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 34944)
`protect data_block
8N3hPuJYVUeafybe/TupM+HQhRTs3LsP3jcu8Rqph1q22PYrOywdH5tMeuY0gB3mdWyPQAbeLZoT
rXTABu7xNTSuf0EDrDhfYaCb/7GhJAUr+uI2CMBErKn4d3xDUb/7yx/KZrYSZ0lKL2QurtGkYNnY
/aK5j/monJlrJsa26pT5xP0D1YDy0VwrJzDQz08wYa6Y80xZ6fch1gaeZZnEIvPVtBnNYHBkewph
HiAQHdXGX3/ADPE3yy7XVj2E2axWTsRiNYxTZA2PxieHV8gcMwFh3vqzVC1453bkrrl1/tZljx7v
rzqwWxxL57PGvpC/WmWOpv7lgdiP9cN18zw6ZcHDdJcVehkb3gLJsAjgm9x109qp2GOsToPRVEVo
Cft0WWFr6WNTcUecFfcMOF/KzgFvRysJSSHjUw3tODja165XfPHws3Roa3Uai4EXDxewHXROCkqi
4LWuNZfTfTacIQ7ZXIKH60IQAYxgYnEkdgl6CPah5nsGxk4sGFfsOg1imYz2rUew+pPcU4Ha+jTh
arMLvpI2eKykNwByIb+Hlq/YNI8vLkw6GRRdwsbvprQIC/Aiu9PZMyy3q0H9yriV/Jb+UEPNP9Io
npJqqdcM1B3eQiFHTVs5SHeX8Mwlsgrg+pGrHjytUkbs12+w16EtWlB4nT9uUmhDz4iCwLdNrVGy
dSm7BzYIznL3CR6EGeIDSo7xgjHq7+GqiySmh2h89tgN9xNI7XDyrIKKUwQieMIv0tSG16WBb+QI
nQM2wl8BxfCepR6hG70L4yZSnupK+KSZoPyY9a+EjNIypJUDy1LTX4F0Iy1mMUCk/aJZ881QIpoI
/ankCaH+TRrCg8eCqBubCDCIfgghqHtC9zGq/PHckq6AQ6gdPfTTtQW9cDbvTMZZLjPrA+J0JO/7
Z/0s8O4F/8dS3QPGGM6J649nErRCnC8sC2tBqslNQMwuLSB0LirPy6KrZ6mYrlNeIL8l2GPDwN7z
H1/cNvi3CXBJTmeWQNmUEE8nbx9s16LqQ/EUpO0OuBtHjoNo3KR4SKz8c/e9zufH/GBL+DdHOOx+
1I8OrZqfVU8+tqsa76MwqsQ5aKco8HnhrG4ZA0p1PvM+fgCTHbetn1HRnKm5iYEz9MwUGDrgLERO
gAs+o40UP7JXvRchTf8CNBmyCjCHSTkJeA5nATN02lgegzBy5UKIdCPXhs3BtIZS6w+so9kYueYb
N0ZbVSCRZxEATeZhTaIChYq9tavzyfzfUUIegajJPpaeXsBuEYq6kUPe/WAiIJNiJeDvDacuH6Fq
0ds2uip78SWKOHSLLSimhSZ1liAdO6qkATJwrzkqbL7iN7YIXMufiSPooG82gdg3djtp1zAu/vk6
KQeaFjLrhcwCKhjE6XHSsTuZGVRvUC57VxlzcDhC1jw25wLD0bN8oDh8t9glERVI+w33lhl34LR5
7fWiuJSHrciqt7HCDaj9MnH8ktaFX5Qa9mAW2+/Y54tql719od1k7qD4+O4TO/NGZj0T3SyQSkNH
+hEmLAmb8EZz8+9//snJgE6LiljRZmh/at7c/Ls4LwDE9xxAj4E+EHf6IswF9zSx/XJMPuxcCCPq
MZiDMvzAn8WCLtUhdgzPISoA482Ftsr75iCjgYO4NUp5u1O37uIWh0hXA6QYSUcPRX6qSMjuCxo3
ASFZw9bZ5z3XLGS/OB/1w/RhWiHMjd5uUzZJyqWGKyiuA6XaVdOThIx2zU7+v6aBL1eW9EtCMHwP
wTXLY90uj/rTdwqknv2GYhDZuH3mNuDYosn2bjVJ6KMD1pX8pRh+xW7BvHdwDgNskZ7zTFljDx63
4RaR4peqkP+3F2VX+Y5s3mKnhq2Ij/12swNwXKsoKKMrfJpgUfnyjv4D5tdGp3UDGxthVZ3wNinY
A8STL/XB73mYpOnP6ya8P0v07STviDjluT9rqqF0OOWBKihlPhD+NwUaJumfxW+cSY/obINNHFwb
WGDMLavwYVnndMb/kuF9wxbx0kCO6m3oDAihqjuMX+CpcDrb/C5GT7+KBwvQllsZ4zXj7BHqk2vt
doe2nwuj6Bplxfi5YuLvBwiOt10TM2+aaVsBrgTr4j+jEDAL3WxkpTKwYdijnENRPCajxCS8Uaha
aik227j55JG8oiBc5GQpjMJ/7t+Po9/qlySDG7UIV7lQ+oAZ0HaCbEFgds/Ni7hSjnRhrh0+PVMJ
90rlyNEGTpVsOaMNu+c8MPoWcX4KdaT7xnB9JbTCSN9136CKsTPb1JagOqOtsrviiApgz3fesb4G
Aa1orIATOUvn6594D7PkThSZxmY4zjj6i4EtRb2JBHKFOWEHFRjcISuf1zrY041lC3WW/vGU7jD2
v6o+uztHy+h6CWFhCW8zZZPJxjm+O5z+xVxPJ+5mqWjz+TDxacPYWSs28ho6CgDIgH2ftkvfLzI9
LKEgplm4X8JQEdhJ6e/A0waHgq1AWBsx4XMRrMOHksujZ8sKltn9WMdFRSDk8PjGYV7rOAcL+I2M
rXWkKbqcT/3OZuqfz0NQayfj2zYQUY042cMwPrd4dAA7ifh1kxHx4MjxO1I6V+qNFXgCdR4l31Bh
ykhtXbh8rZdn4SNxPVESEnr9VMF1HDaPsE1J8TgGWF4/+folwITrp28AtiN0tM13LH+rga2ErTdw
jTgLqp3EsnERz63Y6n/v79l9ny6BOZL7BVH91hHAkUjiFp/8FLleOaoZ+vX58nMgF9/f2jm6P91n
F3kwbevdqB08x2a5sFKbYQQCbtAK3sgkZY9V62/sv1GfBQOkscT7cKV8sg1Nd8BNsCcW0yEF9A3G
+14hL7NwGcbrpmgKIJvzt+1ExiCMrsBbMhMAw53hswmBSHdhOeoPBM3YBaA7T8r8TdsbIgtAZZjZ
lIJ1RGpxfnUxXEXW9oGvdHknJpUFFJrlmxvV3p411Rd0xvkxX7+tTFHZsDoZQZP+1SW0Wv98hKBS
IE98dfcT8j6jn7hPURXIoyMKl63eIbr143sDBNST86Oe8H3g2XugHuPiBkaE6UzAmnTz6yZglxbK
U+4JJ6l8xc1JM9vcJNAkpnF5CY571/mX93egRD6rMpUDvgefQZdRCY30g80tu7hoox1ztAu8jv1J
EhNcfm5PQs/QD2ujiH/gwmMVZGOFRjbM3bL0lydDMzAX/p5+ytFQdF0Ln10uQa1tEHK+LkCLVZ1I
lDSUa535ZK+1U2sg/MZlNGzXPC59ZkWvGzBE6sOIVf+rOaLdq/O+XU6E3sU4Vo9p9/5fEikFjRyf
yX9Z/XOFXSSIwsBDNFPJIpheYTG1lP7NFoZH/S5V63vfc3seUr3BUPenBzlr3R+8moVhJ+BBIm+Q
Trk1iooQIfg8w7JLIMBqLYVXIx+ZkRsA2Z/pjazwpAgBrikMG05Gign+ODRb8wxp88v76WPLWSkk
IFpb1FTvJJnaU/QoWtguf2JsdXskbbTlZhLskys7LKW0g2kW9lXJUkyX+wSdjwz36pfrIoc+awH7
53C4sLyfp8rsVIBeKClyXc6Pvy6kWmyk5hIJepW28k+xAlYRdo1f51zBtxfDXYEy4kdEje2FXGm5
YFpPdm/54418mnbpT3WEgY25JV18Cbqrl0gH/3sWOzZGJL2xndBPLXLukfqabGw1Q2YKmoyrg3ZB
AC+aChZ0SpMpvdHYT3pZD/Y1FplkP9eu9qD4q4yZaRH7uSE67Cka+W+p/Jsew4NatsW+cVlqRcmS
8HMrKeH0WjbMF+oQtJ93H+F+HrUvXQBJTQlXOGeZia5FK7eGkXPBrJ3f1BcpswMwg8bwwMsHlKv6
BTomnlQq/VSVDDNVWSIjemAnyjUPP/eHU7JL8ECnk9x5+KtqEtXepEQHdORa/ZdSt+XHPEC5YWAL
XYu0nn8oaKp5rAQ0WNo/NpT1C1fTBbsxQ0ao7GCB6Awy2r2S1/kXOD1fcv93ljZ87ZpNFKlgac4E
oSHOQSRuynwMBpJHatu8Xp3NcOWJG5nIlJBWBlRtznxHVPdaiI0pDJGwtUk6K15KvhcaJ+vVXL09
gj9JEnK87jkzaB+8XxBjdtFp7Hj+5SLaelAXQedpL0XtQcJo065FCHKYvRZ/r23SigUEB7aq7wc9
ibDOChFZ5sbicGDwDknVkS4x9rtLdBM85ncdBadLiHUcIM5KyHwRTdPJCwd8nLmc/E8cmzIE5dFq
Lkuk+lS2/kG6nrUlflbr/5a78rZKeut68MF1AoOqtbxdmHKI+913tPdWjZPxGAiKtn8fEIKQc3ib
Zna3xbpL9s+L32e0ShQU0fjKq0CMiqaBUs8bPKNo/KP6V3eSWfC7hcq7mY9TOxnYS6WeXi4d0T2z
UL0UNEdg/q7wx47zuYu3pzIEgSwOXwACV8Xrfzmz+/9T2NlUzClK5qJLE84HPyhAdLV+oEoH2qgE
st3JfRFWXRXQXgr9vnPWVqemfN5RotYooq7f1yDU263ygMJYY1tyACos/MDGRS0dVsi1fwiyDF/c
9voeNyWuajGEdpeDfHA4Gy9p1v0r0TTHLr4IDM0gLJy/BtbkbIPfI2pm/0blPoW1+fmNJiGkIXCs
YGJGKDMEB7XdQ7IoHP6r7cHxbsP2PaK42YDSuWbNyDgdQuWs4ub5USH4flrODW4CGSQVipWOv73t
xI1JgOjS8pxn+s3I+sYP3b0MicfKikJB1yJzkcEvrl7Ucjg0ppAuodB3OkS2BT5QRl5Ueg37iuLc
cnMXv2m5ARL9Ct4NsE6tpcc12Ey5jqvCP30zAAyP4gqUu6p/7HNocCpQ7A9Nd9ynhfhGC/qWvlnS
bhZjuJQUb/pONDSpro7vavEE9KyR0a1jn78kbViBKRhvEgkHvZZoNf4A92J0AxB5vpuf7AtW51Tb
rJt6ua182Q5WyuFUKTUxhZaJuthtYr+bkbxMwb6gQK6g1/nLAK4j1o+P3lBgB4dmHppGitmUwyBV
XAsvrXZdBcxO4q2uZMQsOzPB4FBvpnpebYgFg/bnmDNFzbML87pYpEwBGasBWDckJ3n58SgCV6/9
NXPfcxSZ42CD3o62yoC/QWFZxEMuBrJUmOIdANIheHuobRiq1Cvbltkekh7JbBIC/5WL7IxVC7R/
gj0sMIoP9zdXPBhqdWhtIhsggBrOVW6xHpnkHkWm1FPya0y/jgihXOjFaMBoHtqp9W6sTpcVfVCE
uGn1LPSsqWzZCcWeQA39Zt/RhfgBgO+5DwK30Uja1Gsrg+8aIuDgaJqGpBoD/VBN/2mdWBJmKJ++
KfsJbMQMqswAeg36tuOFSaZmr23juzXxYsay8mU8GSWghdw9ldxTyE4BJP3lrNw6QJyqVMMSeqix
kpeA/8InPvg0WzFOdQ3URnpW9uCx0IaAN6M4ogF7ru66RqV77M0vU2j6qM+uZR2k7l1d32gb6Vlw
pvG1EigWy5U1vxurrFyevtKBFHKPQk2mhIXGAUCgd64TQf2JOuhrgVo1Mt0i4zYRWx9aoSNbB8si
EwkJvRayo0C2+DDAtaq979FatRy6DpiOIjxGcH7QRfa1ARQLnhlYE7SGxykbhe/+ZQB9RVSEL0KN
h65g32xNWsuAN65kGe5Rxz/4EjWsv3ltHAVg6Fpq7azdGRlUlF8yzBTcenLuoyXf5jUWffNCuuoj
0jVdC3huXIJlEEPNKJDW+/oWDG8J82nZvVI3FvxVkwS6aFgU/H2xPORmX2VG+kZDAOJRaZs92D5N
4lrNndqOO+Ip97jsnOZt5H00a4QwS5ioMGDDpPsjnpb5ChrBYyiJ+pWCVhQlvbu2QvWwrg9FIMET
hayWpL23pBv6Wo/nMZ+G7Yalp27KBCacMQAbexPYbcapOT+ESntyp/W4l+r+cJLMLdlT5ogDtfgX
LAqxNJsp1V/RCcT3liE/F+k5XfgNzR54s0YHUZNMKEvRj0mgpmDpEO1PjjPfoFep49QE+cNCOnWV
vJppwHtmOfMVt+gTWbtmKl8G6zGbl4FNZ8omxQYS1Qa5nvI/lZWF3P8OV1I3su2Ns825Dm+Rno5B
rEBdu+ifzt6ywPXVbtZvi4j66iHZKOOsOo7fWdAXi2GZPA/MAII0EgdoMjuJp2XXZRkMabniNTCL
e6extzLBzsnSYCsQHwH/IQI4ulnKnn5VTwpZFGjTPKr83yVGHTbCtNSG1odWEF9nA+aQdBtBaEEq
9crPt2rkyUVfxBsEgmYvVhOm0smuh8yA0Cgz9ej2VMvFJv7CcYAIAPETFhDkEXtP/v7AdQOyiaw5
N33TClihWrGK/zBMnOfVosu74LjvAQa2+HaZP0Bvt3QELHvHYaO6YutELnB+bXu2IvepKql5OSZP
D1hV85A4447jidX/QJ9k/+vclvbiNzjFDeFMKV3jZVmwg3XdwMAo/7rhCDIa8e0tu5N1lnV7FS4g
d99WMu4wbJSJvUbYwCTyoH+5t09jWMdvQ0kg6MXD0oLWN7L3JYWgeZw+8ABdl8DOV4bwkgvHy0U5
QNKDsOEM3xoXuzL9iL4EoQgepkiBQK0l/uWImBCckewZZhsjUCeF/8E1KeA9j3205Aoos76AreNy
7fdsjM0Cr7aFjQsNDCL4qZzjp7J64gHzJovyM+dGdsdv3r90mWLjY7gtqQoowrE9rvgadBIwiPPw
DjrnpnuKO+DEX6DCBkpCfuswkaIPBdT+RiyB33IN9lDAR/XM806KYARKY/tcVgvzq+YOyvPFb/9a
2ijXPsB0KcDcUyMg1mqidGmnF5+RflfkNNn+gRwkR2tCuPtvXXJLFT2pYt8s0ooAiwHQFzasO05j
oCD0qG19985+G6yANHIBsU32ElYzLUg37CqJ+VawE+SlG43BnlenHIYDj9rNZIwG2fp7Y6DO/d+V
UmgflzSFxO6/8cy6qCDuQdP6GAG0soPj18oTRHbKuFYCQ1RyL+U6HsUA9UHWmgXlphzag5JkYG/O
FjO2SOQQJZBNPbnWJwW2009Pr3ZIVYpqzR0c6KBj0ZpV6AlVCDUz4aMKAzkqhSbVLtT9K6RX4dUK
6c6jZIOiJT6quzG5fsoJxJlJvG65zu0ooq8EuOmuMVPFq+w69fNf4+JESJi65Uc+vfASL3UVp2hO
E67iEv2aXtgJ0rw+Lh8gm31RNjhbcEJC+wVXfsTEjSpXC2oHIPb/nf3dlbYsy1HocYPKHpucFMsq
AjxMP1O6SWVFSf49/IIMy5TribP4r7GcsKPkgUB0jqv8wvgEr4MDu91QR1BSDfmzssKeB3b4Ip7H
AFlg4YLXnU8OovdevnmUdA7eyNLW5B4IuMDQLB4EAiIvK3wmVoDms6tK0/YDgoZ81eQLlNjYfTOE
eoIn3YSufG+kcxw3VYwaHRqqyX3XO9fMBJYDAvwSnR9XBbxtJ4O8mWzJOkDc7HemcoIKFga5bGip
CycrJ1wgD+bP6eAtTftTFlJ6uNt8BbFz3ukhS7JhR1yiNTTHej9JYJY2/H+mqlk/XQ6Ql5akNnDq
J5hbp38PG+X5IWkxUVFueDec+wG0jlq6YLEz40OGrAxy1cJBIb4RKRR4U/tJKEOTPm2vpCGX2Es/
7jzbS6iRH3pzksz2+yC+5BZUC0WcD1UoT5WS8sHNsr4SNDgGLlBOY5nSpK6faV4tvHkVorSLxj0m
u7YhpWPManqCQXTFAGw3Y+NNKEQCOPBNCFGnhYGgjMwqpbhNObmdOz2VlziF/ChIehK3LKGwBLQH
6MqkTqiOPhtJDk4KXDiVQeBoOgbwb1a9ZZaOQCtUYVdScolfULgsnOjGk1JJZVKFxDn6gV3o7DEk
XKMOD3qt85H4uiVFQvKOhwIqypnE9NlW8Dz6ItPfY7tAYPxOIvGmTA/dECwYrEP6Q30wSucCgsf0
Jsq0irmwFyJA5JWZXbGzQwD0MrBzDMyOjtnukK6UrYbR4nlh8o2hvFSJz0/p7yBkhKPf1avp1qsE
Cy5Fu+epzZ7eQD3sn7mC4Q+WpjsESJjmlLKmxnQY+wRuKZUmOZLUbyYUsxS0PNDVXchU5ElPhYKb
yjpn34AK9x5cRuSLE34u+4FA+5bqi4uTdrVAxwG9VFrhy6o8wwQj8zbUc1VZjE7OB10+qiVkveEn
5+l42izLJ4cX2Xt/4Kse584/UzwCJZeRZ/mU5EuGU0Qa6Aod9VbhgQ5MQakfUq9N1GjfeZvJHrnG
wTKXJmTuTr3oWbR6hgARG+GwBV6oxJ1UwoGWeTRts0RZcEc+vPV3Ou3MVf13PuNr0fdNn0dK1cCg
jpeH5pnfPGNAH5UKa3sdD4SqzZIphjznQIzc+l1HoDXC6ozjmJwUZiAsLb3tqQghsJNm8U3yz+XQ
ScrSBMYxWOG9DK+41O71Fty/sXFr0saGTkoR7iaC8s3Fy/hTrCxsv/1uyOcWFqbqPgxUDjm0A5Me
cC9wfNcarHoz6uJbXSH4IrpTLGK+bmDsWBaJ/BIPZJ/pcFiqW5MpK4DXoZ2H+wWb5GjkZAO46Rlr
rp4xOHyNUcOJE1Ks3fyrocl0FlgsjAzv96Skf7LyOErQTwPWcNrOPkCmkhyuFg22DbcqiiVve4kP
cnSeK8JFokki14hOM0QAVuY160YJjaolyvpd8WuTGhqSoslubytFTq/j82dwpJCi1m9XN2PueQj2
m0s0V2nPz5tvPwgPTLnp2AvVn1VqFtuLtw2pq1+C+8tn64nVKBG/1E96ZXK8Jg+UMo/Aw/0jiKRS
Gjsz/cUqFupe/KYG1U85g+7cZTYKkkUIcZEIKk+ESoP3oQEF4wEG9BCofWC4oS6DaCJg8HyPBkS1
orlEBWmQ98oWi3LfTSXaeZvKMjpu9hFFT+cZeSUFuV0gISegmDXHOC2a14VbSNZ9mw9ODLB4+wuQ
CnltOqxNpwl23a0n4x/NKhqgqzJoFJ+grTTypD0UAJtBZq7RjiVi4bRIAz8JU+e8hMWJx9NsaLYj
cRLpagOnP30KhaOEnYwASkCemG9FK1V928l9mY6sMZENP0LLKV2VVw9nolaeGTi1UcA8o/QZregN
XLys9LGYxwpKBlBK9giWKyxGM9l/tWkiM7sYJWjNtSysFCPNcKAnJ6L+GhX+TjFThyGK3o5vqpt/
zOslLzFHGnM0iziQL6v9JaXIAeJ6zEu1cOMiDuU8Y+gTVtWEezYrieJCCK4qwPRXv+3yi26o74FD
mrQIygrYsitrcb46FZClmbXckyr1EW6xGzAEHOBw8hIZ2Z1dOZBsmvfD4li1vx1gC8BgpkUFZ57k
8KIHuK7DUVcmn7ZB0guOREfPccZqB/tJFdq5Sj9wkUMsI2pXWlIxJvcwCkB2Ve/dNOSBqlYNUIP/
dqBoUll16l51CGuFmEYA74nrlBlSxSZvgiu2g4RLEZKTWsO42yHhyseymxd6kmeTKHnvoynejr81
Om2kSykd7qa7/FLaGXuwvJQthR1OvqmyzqGZpapoFnju4IG2gisy7MiDIiH7qTe7MjR0qNQdyV8c
h7RkgFG4wnRIbjPTOzhhRQuP2RaqhyYjV0N3G+4HUbfvvp7masBDxzOil/6roVFlf/xJwrFgjSH6
6xaNagituRlQZQCPu6IH9Vs98TesSLgZuo+x6yC5P9P/IcB05ArWIml78gTuXbyqhVPy9zI8z7XR
ec0Ws9K2i+q2LJ0oT28Fc5/D6GtrFVPsNdcAOL98EV/PTCm2QzroABDU694seFoETBdKfBUG6Xzq
KDQq2UXD2LU4AHTZNrJak3Gn5uQ7nyofKxKfdwLFLVrGvsgDddYqlepLOk92jqZ1CSY0KV67kttC
nMtQHo/bn7erxGLPIizWcFtrDvDafo0F8f3ammz4GyXFQwJwd84hlIOxirq1qh2uoUr3VaoIo5Ij
AkAUK1bxH5xvbA56U1H9MKY7TGhx67rhi/hUNphCRUJ/3hbQCVllNhaJZI2uHzbCQeeTnFb1prLA
gidgmIXAdnWltFbHQNZUImveCqO1ZjkJR5f7X7WHmGiCSCQz5n1K9xSE5XvwKC2Hk+c0vsNl+ikT
D6J0VkdEJBwgCZngu0AlNoFY8oqTuIVSJHRn1dX9CGnCXHCwgUwiBdAWVUsMbJT1yt+vFVCgi4ue
3dCdw3MhbsMzCEd002Lb0poTRXxzjbtAcg+EEDxC18KXapOIZIizUHHvuwfDMEXTCl2jN8C/ULxo
rLjTbQSEYSsMFg3ZLG2vFbd4hPkFAQR+1fJ00wZxQH/7lkiGWejz+wyKpfZVQZkUagAPAoYGpeQs
PKX+pqexGUtlU5u3ud0+Xx0btv/HgEmf5tHwLjimgPWHWiLfbmYTcpkit2Xf2+z+y1hW18ZzXKQy
RUX4LM0KhuSBbsTfhRNA3uAcq8Hy0mIxbV+zc0zhoj6s0Ocfmd9o87ANyu0so7kX9l+tdrrM6R5Q
O0D60VyzdN2TCcwAL1fWzQbYlPH6GOwWwUup1eyk1QeCP0fsHMscmL2Dy3wjin7GzNpdgdvncl+8
RFrERF+zqW9dOM06HxtaLQzmu9bsPRkWxYGUN51qtzn3ygYGSqpGAb80/7OkZW9Q65tsfaRcge2v
zL7zAF+rN6lmVjM4klb7Y7iEYlvkwGQDqg/AzBa2pdJ/7oLo+c2QVZp8isBcrU0ECbkCxs30+ItJ
tMN8xrrVw+Vkd8HmvU5VVIci1RKGXbirNknntIK5K9Sp1u/tfhb+14DcPkO8AQ2/mGHmHaYvn/jX
pkrO8NnqGvt3sJgL5nZwUhWlHYUdnRLVPboePp9NP5hatqyezXDTRGhB74c0H42nVqbSW/WSIcjZ
8YoHVSBFqh0T5EMW3VKPx8gUZjPenBVT4xBR71s4vDOqwo/CwohKOXeM1o+SeBu3E86RsnTZngDQ
PYIfHIQD2PpQrmjNiO2KxNeLPdMr8o0tbgoyzhMkXPiX+r35G2txyoHYzxLQ0kgtAvwqumnRNnuf
UqBNQ4nBt317Ryw+jRJ2Al7PmiB0oquLf4CkQx6fAoew3Z4rxfWxOFkllvo9blKHTiBRpwnnRYXu
QM/wMpEhooxtdU/hZHeYjqgG5DsNNpZXVhwvGGRyd8wZb3FePe/l9v37D5PEmrNDxJVEqXsizmnk
NcoqKcj77ULO4omHVng0+4SIxbgElb85EWpakBx8d7+A5DN7zreht0oYtMxNw0V/45sJZhys0Ilu
7BACdMoorLKeFRfHyk9I8JeA9Ab95Du9TEFLo6hHPr94yvBxwkG8m0yTkwBgpHc8wS3HCTLbgOqT
TZh6KMY9SJUP6M6ZKhP7FIjyZM4PI/9TRO49Ma/zCEnrIaXbW5D2MCcxkZQwlcdH4Gs1wa+3O8wU
GO5DaSUbxMwUGHJPJbRT4vRx2DtPsRF3PpNTtpdJdVGqbot9+bAPzUjCkLPX6Eto5WXncVTY8hXd
zANi1s+hcSzZY7eBQeqILgrIEWDS1mWayrbGIFkNrWSA0eTSGupEsC2WwW7qg3bPjUGKDPSPznU6
SyjYiiEQemS7zsB2Qa43Cw9zYDB4wadmTISClrZxTxqsVizPdWKmt9/71y5A8U5bJC0qqIPt3/Qn
Tb4hVtCbAjcYD9bfPl3UMdoKaFzFOwMHAej/rcjQ0lPE3gGX7gpzaEysZHg+gyWrepZZ6KHZun/K
7FK1GfIX9XBdba+ZP8KX3C4uBSG6thRXj0CCU+jIJgrNtFEzjnShO+w2Qa5MY9fuMYpk73R9BW81
TAHPoyKHS2Tr5Lge8szHZ/2NzGVBN/BFMpcn1UZckv163yRqI8PcCFi0Mp+Yx2GhqP5Is7tuacqj
F5WVkq3rZheLrh7fM9W6ECrHYRBI746HWs7zByvHeDTEGi9U8n8HaoWu2+QpS8FeqhAwax15a2o+
wXwUtgOyEyBrarxcWwszOdb3yeKYKQjsh6vKoWx44Bfy35otm3guuDCcxQLut2fjAQtY2X6m45bn
enlvkQin4vX5r0JdSmzcf2V6dWb1XBClCqKRE5EiC4Fo2vVPcPA3W7ATOJTB+2srqrzI3kqZsbNm
hvblRSYWgm9bdDND1bgLzmR++dz0zpSllpiAEgx35PeJsItNuDKid4UUPxNX8G3jqQaMx+0GVfVp
gAo3PF0XS5TYJC7H8PC748rY4KG9MgTslzPtpvm64vjOhDZ4+b+rk0qivnxw6bDmePoHgQtD3iKY
x77OmNWrsN2s5jMr8ErBhNLUVQ/AIwVWIEIqMnKcFhxnJje0SpcZ6bM/kbW5Jc7p8aGQYu1srPsk
MCsi6HqAnSjH19S5w9U53GpgedUo/Nl9fwlSqUi+4ufYJoBgk3xVoFVcoyR7cRk0Qo3MuhOSsf+P
GKqzmWIVQjrA1CPm+O0lLUPgedZ03elxg7ILX5JBA2AHiorqMskj3eR28IUXUdsC3GZjok1DfCF7
ctxnT0gUdCC2bhKP8J7MC9de36lYeOnAvu0hrTM7EseEyDXn5mf9CVtRm4vXxCMY9jY7DRv+vxtf
9R9p1MrXRnLiAJJUmjDGhXbZ+SGQvD814PwbUg22pAxC8ROxj/rtdQm7Q02LqF3FdCkbcxkbuBQ1
AOCmmRrsf98UCEjVgyEGYrUJKY+uOAFvWh0kdpR+QRSRqqM+DZqaFwJrzUphRqVgYF7Q7xDjvTaN
op0abXvlMKOE9/wXOsipDDHbM+2RCevEUVfeJabELFbL+QjtOT02DFsLY6MC9X7JFrseSn46sUW4
ziE4XSg4udPeriwwJ0aFqrQls9utjlmVr15JrcmcwSzQVO78Qr+6zyAmfD1KM3znqCkBs35ENS+J
txHoXDrLzc/3TaUaKuusFhTcuiRiMXmSVK7hv6o8JSzns8YDVt+J/T4pl54iWpE7PqA54nZE8Qi6
cSqf99/nUZObUPeto9FBehCRjEl2PoRvjMSPy2kPm9pnerDAWygw9Uc0uHgafwcD3MYbnfTZGsgR
PfCjTkfJEnG2r68Qqewn25BnZZk7FPJ1cetqL0nXV52lGwhX31h0CgX6u3w6xUlFQlvj3Fu/MOCe
gBe9VQA3ll5621Q1OuY4+GUM+s79zU1n9pqd/pGkK1U3aad5zcsh0BMEefXQMNrk5O5/2fbuSBUS
e66NMw7NHVQBnrlng3mvQjFqdaWbbMYu27bwEeuwUa/R89vJQcgaAoa7TreeQ1Tv9O6ngkpOajwL
a7uKkpQRyaDBSNNw9BFRpcRh36AtdJZTLEpPpIrtZk5bapAwutqlMLBborCiVbAvQy3Ks69AzYWZ
tgYskEROomhc3h86dYPpzCcpLjpq75HgSJpe/AlftwVLzgc6OfgBPB8+nfMQ73i7CVmx3xALmE88
u1S8GI0GnrIGyjM21Fvd3/cYS88YlZiWNOU045TIW3KFnUor83ExHi+stK7MoTJYKyU37R7XRfHQ
Pka2NBfwn9+yoVllhOoT1Drai8ppQs0M4rqrvxJvlsI/P228hg3CO23rO2PHYHu7BsYCMnxfdu2l
RrK+m4N92aWqTwxf7DPQDsqEDrVi51Att2TEQe2U8ZlacUNP/2YViji2pgtqgW/uK7v/H/MdcxTT
Xndm4LBia4L+aBa9PdJsge9EerDWyOqdD6OKY6AmiqpN/94teEHNzoWlERSPHYFkdW30aAnnFF/V
0aFhJb/nFHxLfHJ/eFmYC1ftuIlEjMUrhhMiInUMfxFrg3UBAbCozprLoicApX14lZt3uFDmOJQY
08zcsOsy9zEwBmndTGgPpsHiQFhNrAacFmccg6zTJw+wlJG8q4wccoge2G7KhldOE8Es0QNwflLk
Y4zc4+4vrwt+iEU9IgI3mi5NYPLKiIFuwLiwqosd2ViinUAuvUARqnQuP40frgNrxzX+DByzCmB0
XxTLTy2+vrsDS/Vz6q5V3B03zs3Rs3d38/HqLfv0/KHrABaVcds7pKb/Ii8wQG9oKzEekhrFBsvX
QrzoxzdlQzJIBuO3RCPmy6327EkPMEOOuUvgFaKMq1wsSH68DoDLsPy1Ub9hdpUkxyfNlt2UfcHF
ajP+nmsw5Ene5ezAwU3RhzbM0EaGXaiSuGbYiM/nUwQFIbV0D/W3ZzGv+dz90wJYduC2NXdaR+8w
goTa7AaqQcssb1hhEBw6GEz9ZV+m63+N1Q6putRPFxLnL/04HQf4+x9OoTnGyb1e1Y5HJSLj3xd/
/r8MicibAyBlCLI8e+/zqeeDnCQrWpX9Srq3Vlr+W+/hG862LWsJ1r7VY18wUe814UgwyU7ybf73
Ufj/6mFSlBt8GlF6J1b1ea9BbGss/ac2WgfdD8tv43Ny+8/EP/5e0sYkFDKqOkgISCWPDf2DbQYA
6Ii3P41DzyUMaaMDSaIydzw12ESdANJD0EbXKarNScaIvrZl55NrczuniQ5T/sdHtHgfdg0CLCRK
sPZW/4FZvRXndlAbtNlFFZYQ2gzAhZMfmFGDOIyqR9n5lfG03hfoyQ5NZFtboHr+KZc/I9+oIXim
r1yaf4DfSYqMgLFBDsz+CgMpCUV7FaHXGLiX/gHIw1JJcDwPVZCnm8jenA9BFzHhtxJAe+5lQfgd
oCQ4Dl3m4XMDBwXsILeCGiULq4Z8D21ywpmqzPGEuM0YVe6F2A1v6cUnjY2OFXqWh4jAqkx/GnoS
CBGvN2i/KdB2foA8XEL2VcveFzdmwsr/k71umHT5cp3pePGvlv6vfHFjzoSUCcHF/filXTbjpoJ9
7O3tlF8IbHJUCvz71LiS5Zk3bZe9eGecqB6bEtBbgMNojnvX4ZYDPydsCwPOF93Mnhtw9cbWQNdO
1TSxZcxl7PyzfcCrnY5t0Mq19UStpW8rUsFiP+2NSwyE4SuiQU4dtjZCN+iNuer1jkN7gDj6zdJ9
jLRlDHjWiPgSpoYvIBwkexQQ6jh3Q+8QuIwDPmxX2lAyY12yEtvpX0EI0FFZqn1sxbH8QtsKqUVO
KHpZGbUoADY7b4MP4PKE+sMRIj4EIyMS3TcKaWyyJtzbJMBPc3RIpzv5hk0XUheItbnqk5z+K5+a
1i51mukv7/NgD3Cn0T3j5/WN6qzEP1rwt0BykTDGMi6NdzXUWKO0jzq91TAfiwKc70hJ3j8hWjAW
ch/iEcUzBJLl+B/LsmHRvXd0jfwtye+rWS8YYuTAv7Sj2+GHVAC9pv8/NIywI8MFKqNqlRZrst+U
YPCCAJOlhxjPr/CpAOLt3X+irXVZV1I1d/aK+kytaYFXStcA7xhDyih8LVPneS9s4k4fm7cTcxUZ
IaZuwdyX1Mxt/iHEgcalo4d5XM2lND4bOKuVzFuYo62ALI9qg7/sRk5xy5gcBBoe7XfOvOmMVBAK
fa2+FHsrlN/nDsO2fgZ4pAJ/GsEEBpxvkw+n/UOO7wT8ft4/dZa4d11LZuChX9p/ppdSmcYiEqNe
npp4RAoEm/qT24NpIK/ikUyOuZbHFaOZ/GfmXdXGIzKPUUBsLRqy3vtU3sVCIyCjkxpZOMcb95l6
R5rHkVds8ju8MvLOwiqUSaSf/hWyIoFUhn6uWWywHoEr+02+3u4NNf3Hszne6+dFsMSCo1KMBVGM
JM9EJpvVrOhnPywzT0C1Ma9utJ19UWBk8NVpRByflmQhyaGoJsAijkAhvYgHHS5eopjXSLsH2cal
019zLuq4M1bdxv8VFrOYp+xCtUqTY6FeljgVmj855DzoyNxhyoAYu2CapQHHDIT4SaOhAx2fyCLr
nEi2qlm1N8CJPDy9/lmA2QIPt/FlCffgQkWT6J5mu3OoWzNDM7CExkBprQlEXhyN/td4QwTBtunl
hzTAKIL+pcPl4ZUMt6DPjPFY5SnvayxtqL+IRsZmCR/s6FruEK9uu9E8HXBOYtvk4LUo3TL3lVRy
TvcxiWi3lNztg9+CzOy4yL8RyHOTiq56pHMFyeNdmvHP75giWl/q5K/84Q8Pl9wo8oTpwyYpOtn1
s5s0QV/oQ92aGCpolqKq6hkc9gTpL/50eku0D6ubsUauNJap3O7OytoFYW7TKbDI6JyRHpe45Ukc
KL4tJTkWE2AKih/ylP94HfDdLtWqPyg8P4QmHoAkAM6IXb2Z25s5J0x+u51MC9s50+RwRdZupyqz
8qgOvgoFv5lPhCMj40N1CVliFrQKjUYg5B56ZFBbSfOOuleGdy8U/ZT+dtJmEu4Jh2sEDS9kOwlW
5ij1oNDNOXkSe+TH5uPPxTVFIZBS3jWz5TpjhD2MpbBNAhV0/puD+vVm4H8akiFaBMgOyeeO8SlC
uXVDS0mPnfofDe0ZhFDBOrdcXCjtwjjdhgTo0ID59GdoQnA4mrzdq9c1/kEfLbAYjvZj6FM5NDj6
l0s+vXVYPrgCumoyqYEQh96WZzJO+tGMJuQqdJq8IU19J7PaFmn029ZSucDblrh+BwowDrXPZKTM
9YrEsMlWwSdwg+mx54CVoT+tZLOVedstd+tnn0gy8h5Hmbtkl/S13NVa35+eobpr056dzWLqGJRT
X5/bgvesXQNOKu2Y+IUKD/MCso32ve4nMB+TSVd1I2geSU55Qry4Lb6k4SeRlDrAcowD006VjDwu
b1aYrFl0FAHcTJ10gak8xydSmVMtmFTZ/7XT0CNpdi0PJMeKtPrSCf9IW/q7g06bYb/a5lUt0aI0
KKi9TKK/WqA5edCnd0ysW4EGVkswifZhDcNqZqMIisAmUqkzBBUpiXpYVDEQBCj1/5MX1EbmFNR3
dF7QLIaOtspGbtpI52FkFeFFRLCvKvIKVOv9UqWlmVItjmuyGNaR3YL9g8XLi+xG+EaAk0CIeRSD
40MffEd3m9nWFSG6NDAh8AevuzDWczzoklOhl5DaJheQvRoxGgNppwBOtchmZvfnJUFMTjw0IGcF
9sPHMFbIEvROJQdXiOZaaEMybcHbwWOAXcmHB/VsP1lA7wT7jve7BsdyG0hY7cwgNWPNqoDdCzlJ
GDO69C1xO1fTNBqNlOSUnTfgLUM65ri2lhM1Uu0Q83tayRhn8qp1XYb6wLFnjE5bFfoz1JYa1/9N
Dj7q/pz0O/Oz0wdwzXOp/wUU6g6c8YAciHke3bBOvQ/Zkf1P9Y8bf7P02ebNhcPSuoluz7NazHXb
fAaZJ2aPqG31rrj4LOM03Jak9IN9xQc1vqeTu7xq6EgJ+kzxod9J1yB2XJHXRH42M0eIRxbIUTHW
QNI+YiBvuqGkgbTXMDDnT9YKSp4AWvfbi2Kku3P1cl2I4eP6AW+/k2apNDWPWr/Bd14Pw1PLN3xz
ysAC1U+CVca7eiosF2x4T4pP8Vhk8Gk4zJCFll9k2XH7kxZF338qjvWou9El9uML3qbj+6OB1Bxn
0gcIQyPGFjomr5IEhDOgUOXo/+e5iO5o96F7lZ+pzH8VpMDQbHDk45aTxeuepXmCuMr9/Ndsdu3I
Rd8TMSWJO4zdM8FkggGtq/VL3OENTC5SThio2Qgyx+/EUQi5htICRrp5RukfNIdVeXJlzKlWmG+2
eeMYmZtowir6iHmNXwDjreefh8XrsBqFLnzPPeXiubTsOqyFsurShZZHJz5y0IN+aXmmcEs/hiZq
e7E4e/2sReNkSVyD0liC1Km++npXoXXzb2jkCSMlZsmWSD9MObzwzoLUH3JT0hObgWV2Tkh5TpeF
BsIB9Nt3oBzQgA8z3/exrU8mhot2Ig9tI1KUDr5BsXaRESkz3x/1LRy2DWqhMKPKiTlPAyOrqHuz
AXeUmMInzQuEyff9ZTIqDZFLQfIiDfdSGPBYfEmRqQKw5pueY8zAN6nzZZRMuL7tVqDxaF8nQ/0o
KpnqqUb/aPiC2LO0CZzX7O/xGBZEj+gAx1QrWhBIgMvDTppA+tl++v3EIhMetmyFZvKwCl+nLh6j
fSl87GaTJv3BkVBzIQGJvNJaC8UA+u4ZuSJ3CdWWxRLE079zKQzeh8uvd4FO5J/naVTFaUz9Fu5V
hdrqxlYPdwgh8p4KHsZDrvt++IoDY1R+YEC9X4HRkzJEy64hykOZ6HJCY+FiDWtgdleD/bYoialh
H1RVv3uoU6hOtPFoYQicqtZW4sO8xLte5eLGTztUh5zfPiw/Fst+jJua3kAIzYECWNmtIFDb5eqX
/tUHxzDr4QkVBBSioGKJ7djnK0e9b7AnQodt3Tgw/YrvUDjBoDHkIVnIZrZiIUaMx6CbWY/GjdJP
Ubq1GF/2y8AhPjEpPU4QqmhGGrxzFFslsA/i0wraPKnL0RqaOhwAAbsXGBMxL3hm0WRz/d73Kn7x
Z1Hph4aD4tEqpkFLdJ5nN8bbPPjDwn2q+hFPET/iuVFYU4mkTqJy1panVCVb5i0+ECJZ8dCXDV1x
9F4x6k2byOYl0lfeDCA0CFQXe2WMkR0z7Xf6k3/i27nkNzkr5GTv4rf70OQTqPvPkoclTaruOKlZ
Hw9A0yBPOvS9MKUz2CrfBvW2xLqhEEH8fiIBNPalIe0ljJoAjGrAjDl394tTsnO4B+j+Yg1PQJZD
f+ufn+XTof7QiwiHDeis8VQIYTSFCU4jSkaHrW0+zT83nk4OhYzCw2hmFGUoMYl0Eq+E5V781VO4
VXnmWn7YQaLeI4Cz+rLgkJyvU6diDXUfbTUh8uRuH63svPGSEL9iPeC4ywqkKS2YOW27lsQIHDcV
EJItO7d8Iq9omQh/Q/xCUJ/w5fCClO20E40yGPNR3v3bMOfd4MDJJr7O4jg5hDH4t62WJAb5DFQ/
cDsFUPSX2eQG8y/E14cjlfsnqvSPfkY49ZhbRvZBte+LWtBExLge399JcoHASWqN3aAQeAprcP4O
85FTYs2LbpFfQGOV3SvoHznUYYt4U778YiplojIV5f4yyqXU63l+N22UHluVw0CjQwmaTXdUPKho
oec8kDFBjRkcpXIBnHDFh9WGKx2AlI3KH3P12veZoe9ZfnnJ6iCO9l3ouYrcUKVUmOeqb0aEWRiE
kVEVWzMNPpRrJPHf2v8DwYHOFMgDlsvaHiRAlZYxTDHLBum4lTFLI/4bWasn+qBUDb6veKfHgP2m
Ryrk3Ah14Y5Uu4qdEue6kU8sNr6dhLg5KMhUKspISR2xgN5A1twL5P9+TzigupINDx76am3MhUXe
YQGubgbF+Digs0yJPVZTkl+eh7cIOfCqLx6o3jzp6i1KVAtoCCqhP4m9Daw4tlgf3lWJRlVDAGrF
BxIonmjGr7dwR1Qz89CGDUMqFm24KiFgPa2x4U/2eATsJtXgoG7c9/WpahZfShcriM4MUWh2RFmV
/MD8VgOvytGawYLzvRpS2fT0SO25CFKtSCLwDgM/Zgs1KDdJ2n1OOlftWZVHpG4EeOFy0Wa+Proa
n60DMGX6wE3WdBWsA+Sng30rmQ0hZJlhD0DRGFgDB3kj50RwXF6myTHNP6pnCrSl6+os3EBs7l/5
+ICM+Kf1ydoOWmq6Dn+wDIG72y8adV0mqrnkxgWdraVVW19KqjJ3qZ0m8nxFH8IoEh4KqzzRzyJu
2/lZcE6cP69avLNo/9CCiKlwqZZvsYE4PJ51jRjHu543XonlUDgTPSTZMjdV7p7aEPxEXt8mttFZ
9Uc07sDD1RDFVslmrZSgFbHmZBzebWGjTTdysOZuMC5LyvMbzOEB1vVsD4WmOwaEx50SKNv90Tk9
IPB2ThmwMdtx3S81zOxEr8Miy01KbHhBhh77dX5LljOYqvlLMzC4fL5tttGkQXqQPZRu3k2kuG30
dWqDmoJ65AW6aLe7LTTkZCYzQ4ftXfIn61Ox6hddKemGS++nucjdDUJtXXeHKpcERzy+gQ023ZQv
EanzECn3yoRwmcDPasd8Adf+AoNSfzF5FeqwAcGaT4EV1o3FQsoMRopuNI06bFYJC39AJAywInHl
lWQ8uuFBvebIjotLK6buXqAt8eP6kR+d+nV6sIb53stmjl3mPSL6vA2gFuZ0W4tLBqV0TeAuF4KD
O9VBhSXadtXoV+XSL5kNoUn7ShjCOXSYKbxvDhORXo5MyaXuIy65kjpfh1NFzVvecRVynxIQSdhS
E+86ExbyNzYyFDJQ/8yFPYTRF3CmO3J1Cp1/p3F7q8KeRXRtpaWSmv7+Qt8DsRFzogWAFSS10O0K
ZZ6d3TxHVfrS/qJiSLutmorTBq1HJdFPdmetjUqHKMh8TjhZpojSRjANLlkGcP340SdCRhYoL7MN
iLdWA71vFZ1OB2GKd7g5Ij3e4cw87C1IDeIODOjZwUX07ixT5t7ajVNSzgjhG0rEtzu3RaGhmSXD
vTiuZV2a6tGFrUHc4WS/zC4+BAlxDmrjpOuFj+7GfvbgkxrqNuws40oWRoiRGQbOFOa1APSOpCMG
y5Zl+LQY6angbHR2bgrMumFRteduu3cLmugw+tXnaj/Z/UD/YGlla1e5xporIWR2S6TaOeQQz231
MT4mYV8UyibcByb1GToHZm9YEG/7vRI20TsDA11oj0Bb1cOY3Hdn8+mHBNycBpyVRu722dFz1leG
eGH/3zEjv0YDokgtYXpstCvPx6o+eS77BARe3EdjZiWEKX8tBhigzk4wqFmctUuePsrJdQ+YJcFH
ZOxlV4bkqiAygGmTYOY4mblyS0VlfaeiEM983g8nXBAPpaidZKV/M8Rt326Pf/uG5ybAJaHewC1w
RXI63r2f6gn3KZxOZxt3dGDBM3V5OdrUiIeM1ohtQwB9evCVaqMDLd6A5191n9am2kX/BR3oJzlG
QvCtDhP/QHwqNtfygL/1++keza2sNp/vIiPyOCKfiqrKmKkLQ0I2pbpsr086kcJuiZ8/dA7RZLxO
dhyNMFBQI3HkqYUwLz6N9am4MzOV9oeOXd1wj6G+PwPM4JArA/ru8xn5HHVKDe6mA6B8s4SmYzC/
Ps+pOXpKc6RG9FoNdwt4Lv4ZLI9jwAugZqXXComVz+F7+3EcX3Fk85Cxqdz3BY/bhrzBl88ZXa6D
VBi9MAzILa0z273bmL0R4j/XLlv5cUgqdrcA0/x7G/8o4A4MD2KYeGuqNqGptasPg3vDtpang4LT
abFAeEH8lGyjFMMDVp0H06cV4rmxUIm1lx0kPQbXR+tZ76fAEQQPvEw4G1m2xrs5OWYN6kdbCcKP
gpr7Vuce4RCBZ5zSWxISNZQccI1HwC5iy2hCqEbRZ+SX8eNo4++90wGJJqU0Kia9I0gghsIigmvC
agaqKeiFby9Fa1/O2SFBqjx45qk556cHgkZHwonBzYsnbSy2yumXxZGtauUyydyeDmp3qXjLDANR
GC6GpFtV2BQbKNXPs+N6Fgr2MhmRZO7St9RdpZ1S5GIu1e6xzfqn9x3zxLOqHAJynyOly4X+1zfL
It9GD+xXUvkC8NqhYYLpgInm0k8+VJUGK1ZKrcq/jQtepKNWVxHiUTc4mthf8pWX2lN70HLHUXEr
MVC5KMsRlVxYnG7bAmUA+izzd1IXrOb1jyxVX7vpD8idiz3eZzvyrLGIRkirlERB5mOgiiUCnilH
wVL/0KnGC7lLYFJs1YdYrKs/qvKvPt4qIldrVhn0nXa3AGLNRvjuNB64TgNl2EZQEeOOT13imvFJ
V7j2Ms3B1jdi8zU6NbwxxZFC0npfK7RlVISTBiFl2lI2/dcuEvLA5Irpp03od5mJMLA+wAXEW1Nz
G+SHDTwI95oXbt5gauKftqifxXNmenLcrEL1LuoEpuFNXs0DSGVZTWZuaTgF40AYbueNHTy/KXXz
aXYox+MqJWkcYD4yqOUfZvWXno/JnGZQf3AFi9jIV6XlzLflfI83M0Fshso3q/fwZz6A1C8Tht8w
PGDAItqX5b7p1UtiWTPZE5IFpm/BbKgCR1GBUQk10jNcUK1Fp8fbiggznJcsWAmFcB8PflVGuV9c
mL8Wi+0+snICU0mf78r5Hp03YCSEWODEKJp7dXIIyyCLj0ubq4w1BXZ0cWlAXKfOSPaRCZNRtjQc
bbedk0Hf98rWXKjcqX8m+wj0st8xtivHvU3/kVyO3484JEzfHOzkCv3xNQF02Z7mp3CXlR1cOb+/
/kwd5FEDl7sfnB6ugOoR2nHg5En248rjpL5r8G25dWwgK1n0Ebr+ZXrXteyh2NqgjPXNkGSsuYam
+Dmg1yMyjfyIaP17sQwjbtgf4ZDfXsCQBtXXl7wHwzBq1naal2F4MB1C/CySYNwviU3XVStbvrYT
3nFzzUl6DRbXUv5tjk52wT3Hl+sSqT1duWnICGaFGA0LN2sqYCV571L8bu9CBM06ewpyeRo+Cr1H
Cx95OhhSBJPZzHQQ1mLAEKiyfYwcZ1I224Ykqmg8boVX452ucg5SJ2hrweTP8scOT6zbzMliTiBd
0bkLJjtj8Tb/vcIsccjQsLSCQy7ASdy8gv/xYgHGJensxmZhFalX9sDvoMjqtZS37nCMAPiaX2vG
O9MfRdMfRyhocvytd7BVKroh1h25q5MdSJTboOp1PnF2OKoZyZC7SiOs0tDkZ8PM0XzBJY3YTXPN
o2cwSGOSbcmE6Y1cdD1C+RPsIXevw8Kohs8ql/6gs+Kpgmy0lICCxXazQG2RqB/q6D2mdSgnCREX
zIuIqLGNOhXO7wP8TfNrI0OXjtv0ddrCj4JkxzVlry/e6divsOlJWi+wa329KYB02kR9i1WS9Mb+
UU5uBW+gx6F9QvVuFzNdInowS5Pq0OppvyrfVSkRxx8B35664Ffzak0ezFCCjJA/GwWKUDqfBXk3
v0/KVorqhZxh0q8FSZqxZUGK2oqP8JTpOp0P9NdGTzn7RqpOcHarGhdOeFYCNY2DhTUG2DLjuxj5
AOCWlvMbrFUTu2+DpE1cT5jb6SC1KpDYxj+7zTgaUZxp+ls1208uteLvo1tho2owj5qDniNySXcg
W3u97MHo/hGYNCM+PygCGf2HLlkt6+Hs5y5EqBpGe2pBk7+/qxrZtHN+g0sno/gV3CERqzH3/2yI
LZQg/Jd9tZrWxLnWnt7yzFA30yeeQz5UZV3PozpnMRn8F5QNitgJeCQCz6ay0NRjtuym1s2nzT48
/IvY1RyKsqMIR5f6Xub+Me/lGChASWYZkes/WZIH0kTZd2A+7o+Q7fawLcFNPskL/Xy62MC0GIy6
87DEYB9HZ0Sr67ek1WraCABwqWflppvZq0B7OuxdsR0w9eB3kdJmzLEuj9Zl3zozom2wO44RNN5N
TE5CGReOsW0sC94cLfjCQMkB3LgKRubhitnN0cxyIiZB2gN541ypetxDvQO2yjcyYQxJzkb3Yx61
c2kzozVm9EDCKgHGRcIUs7R2u8c2gcwnaX9eaLYszU3n/v4y6VUcolJk4ElKpBGGYZZmb5UMhIIQ
gDo2bZ+q8srOWvRZPceVk10kN/XSS7EXAB5Uhn4nQ6BBUVSgUZVzXNFdN53o2a1jLWfNBofJ8lqo
x2H4I6FyxB6dDECpjSsfxAX6NHmF2VCticA9Ys+SpDS0/2wB7Tp/2W7uCliVsZrtpEwpVonTnHuu
+Jc0Z2QbGPQhKkZyKoJa0f/H5QitfzVENmVj1YHDuHYm3qTTxPORKXkdG/jjvQeiGWioJQB+ErZf
gNnWnv4ecvYm0o8QX4aHjg1R8Ijut4zd7BbJu05W+zMQZhPYVhDkQUWduMAwscFG3Qln4NZl2tF4
icM+KGHoYyuti55P8vDsbopVpqtEeKxIeSOSO2ms6GLT1P8rRX9JOHAN4FGMzSmJ+8UwOIHkfWYS
UDx68jS5SiGHeXvmB+AyurtlnDz+R+LFwF40Hrj0HIntGlUd1V/UYdmCDv4Kv2f8hFPHUTc7I7do
bGA6/wbUFpGbBzixESqToY02O0nHdigudU7PBtIJAqF5Z9NzAiHLRbDIJUD4l1msVKJUnCP+/rja
moHrm8YFIaMT2oZPAnSMZyUWLY221yVlDNzqpn5PuUjT/Ccjmvo5SCl8/aMZmGGJUCDw6V0RRbgD
5BEQA66iuA2+8Sej6dperOwYOOQs+tFtxilrTVxFaHb/k5v5azGlf/Kew8OVXU4Kdipka4pbl6XT
3x10mwPZL7Yv+e3wsc5Hlj88cRO397gxMAoGxZ2sK6LEKvwuol65TIqaocBOhaJ2NBPyWPXu7B19
axjHOpVah0a6pKbPjhGJqt1PoDvtSf0XmPl6JOLPSc+vK5QifzxhZ+xzLC1va7N6UYRjQ7fKsT9z
medegpinANpM2X5aViTag5cLUgROyd7jZUtg2jr1EnJ19Bmc/3r/cY1+FqYZZtAPOJ+Ra8Ip2VsL
O7DfQbvmvz4wNtZKYyWGAgRGc8u83ZnfyzEFW7Myd1DsPBNmzG7K5n3nKUZxR0WxgFe1cd3bHzFN
LVJgWh9isUy6BBTospf5rljcUxFekKGvQswZFOTQg8MWEi8tq0e5689xowdeY7B7mqQ364Ukv+3P
j4CSZvvzxxhvE4WbAusl+m4lxDiK1TinZ8nbCYNdZFAAdi1lvXaWzdT9WphTEosn49ojBb7Pu3Ox
oT+s/UkVeBKuJ6dWrN91MQJg39VCgQ20ZABFEVDB1R1+Qn6IV8I5Hs9J+z9+ljkG/Rh7vYrGiGvv
X/On44JdiI6HnUQZay2lk8shyk7gAyixNJNmJqcb9xMys3YFF12uSnxcotx9+5gr0MuGxajErdgV
o9PsrAKwPUKqLnWRx8b8Pn9cKUrHlWyEFZZ3dLNC3Pln/+yhgKPENSRj8Shx0dYCVt8YuayOuaop
dhFN9QpbVUk3Q2AgquUicHnboJMsosROZOmC3BDojOxojvkTqCDZRwblCwC/kOzOY3C0raB22cXV
+dP6xf2zjLJO1+9xDo+rcG2OcUg+y9xNNiNHzcvrhs8ZDugKwuIF4lhS7f7YwtVaWWOediRkIkXV
EvV0vsVu/FKCUkXRNUypO9dzU5LbBNmWobBwuJYJIY132EXJqxvvd9R/Lgd8A+zZGFI0VbRrp01Q
jtSSYSL2FUJGJWUol5UTyerEzswi/WBnM8zklmG2F1gZaqvQ0gWHYiHPRil9G4Dz1BnZdsfcweMP
qYVBPjU8Y2iNYYzmq1Y/j+aiFJJRv/BvKr6y3Q5TvLYELd9E2uqshabkl+wJyiXyzlcag0MZ+yMH
rkC3j2rW2Y764r9iMQ5v5pYCO0djw8dBH1OVKOs+NfMj0p5jO9NlSDLjkfNMq1SQvHjFjkP/afYR
FKRGwqVR+Nnaoy+N5xy1Up9Lfj1R24d16rTHzgadC2uc+zQ+mrv3YwbM9tBSif7XbwIVrQonEj1l
HsD84avEqbmyMHbVYY1G9WhI6gxL1aigIZheHDW5KSnXgAyn8Ykr2w3wdRgfsiOT0JMvm2gyTQhI
l0jHpoy6baV0lwEAv8A5VvjQ6ppXwIQuD4+itiyW74lBiaHeiy1L2vvhWQFuDgVp3h6zaPTcW8yg
nVEfCPsUFc3cOYOUXqo3dHDdJ1Hbo/521sgEwhRnCCoNVwQoiAoPH4bU68ZPKtIe8vH1Q38/WG9I
tdmhlFw0BpU2SWD/IzWETfU9BJP8Sg1XLfp1upHjGNePX+qxuXB1+DVMcL0rzZG65EgJpW5eSGGM
d4LROOIlQswZiUF52Fp0KWssq4K9419zpt6Mv311Mf4KX+w913vFNIV0EeUh+0vYE4FAiJ1sWZBw
Pj5+k0yMQyxAFkw1t+EFFFmVUt3px8jy42esOybfRjWtKVd9TlsK5lD0vYvkNuHeUoOIZ4d7qRPX
0xxK7clYQU8n2KICm9Z+HgHhgHPga3hA8E0vFdro4nZgqUNQvkvb+Ivpp0gK+oy2d1Va5uok58WZ
9CPgjIwUCnGPLA5SP5uUIxSAa7FXyuqIM7XOEQlOWN7jvki49qLzj3qqDBAUiwe3BNIzXBj9n8vO
6qS6lR2AVedF9hGpOVRTs7gauqxSc8vMM+EbIpbviZBvqbKQ0hg0r9nlCichQByjX91wIarCh5LI
uOREnhsxae3AxPkN4PZBj9QlSGOrBduPvvc2wDSaFqKJzoPgwvsfsotBcYtLV6ls1dhYFeog5fS3
Orx6/7vJgjuFJzF+H4k5iHZ0CK9FngjPTby/kNL9CQEjEnbNFGn1PV6H2NdW23w99uPtfkjYQNWb
7RuPXsYusD1VBpwZlQjXVx3fR/HtTAS4FEvsxoEjjPGSJgQX7gmIzsvXVdMHjxUeVpKveI1i3hO4
6NHQMDL2VLIm+0V3w2H65bpdZgMyRz2Z9nMFb/8Vw2eDnjVa8RhXy0WeEmeGipHvRExyP77znzmS
TkOH7rrxHFDC72/JPKdt+BMttOncaaVUk9ecMTScF5uOKxp+QyF8ZDOfHDAYnAbEpiKDlKpTcNu1
KcnbrWSLKnHCxnv2gt2fR6NBI10bdhZP0bYQRUvYYNIIlpj6ftSNB7gxgCPZIUMl7IzApIjhx5Xi
Q7i5NOaSMmaeQMRBkVYEfji+ZrIF7o5g2XDwU0nmuHd2rl50runhVdu5GbuIjVWN9YTN5CZkW0V0
hLtiHwClW8h1LSur1D83pZKsPMA2iKvHJbRLI+XkYc+NTM8VGlKhlMVNNZDZtoOZeaxdF/J9Qcvx
/VyuHpGayLhpCe0hgXfr0EUpr7O9nSX4mnhJvPOjZd3xnHHGYvBkLo9YGDmCP1ZjBzPdibhfRSRy
gihQcNMxeGkqFUia1cu9zIY0of0dIpOhP7LO5xTxYFwi4gTLIErzVoceFFXVd5JKaehnliCjoM+a
QMfieFrk5REvtR2dMdwSFslm5gzwegmYKZ3axVyyb1LhwP7hZRejGz08Odb7C4pJ2gBxIIqO51Qt
M5oVkeE4gkVDpHXDA4pRymuXbn1kDzn+kTh3QIdL0D7kSHmJiwWCISfYGaPSDt7E7ypiKC4EWgCA
gOtdC1a2q8ENmMIf7JaRYqhV72a+ZjQx79S7CL6jTUkbkLECNfssGG3Vy+40WrdIOoUD/CgOi1uQ
XCuF/6Q+7zfhHEDx51dWF6iLXfKSkF7sTR297M9le9r5CnlhqadTxrcROlKho3AZ6X+hwdejI8uG
QCgU8xTleYMMZixHddfA46oCL9uZqIGdQ0z+bRsl163q1LJODlj/CCLAIMrgrMk7BT53yL/lweJE
hIVtw3dVM58/fv9oQzK562kMS7MsIQhJohl14aVu5vLJ368i2oKVhzDROmiWWIaaM93moHOoIlBA
O0O/gut136jEZM909oNe61aKFK6HD5FelP0KUZoGy2AmilpfqAMnLBOc0s5a4IL+0xBunzsxWCys
8+ZsSiCj0Ui6PMva+3NG0YvtQcXSKrfuCAudL63hcn5M8fcqOJAz3e3p0jUcHK8TA3GIosMmyjZr
hm/v7kOYne6eSrzSoFGWCLrzsom26KfDGO0cUx9J4yEUULVr6gSJJ/aTIxOOmdN+F04ne+rdEsSz
0ddaFQwSbxdSOk+oop7tsly1yNkNOLWqkKZkpsW2SgGrDD7ObEPhUEIcDGoLmuBO9GUI2JBrSSpV
EDxNrj5XdtXwEaO2a+LHPTYLcuH0hp++R2XS4kqv0uavYBtzpAHjlS9Io733LK1F+3IZTsCxIvIL
AfrTEEUh8XDEZR4h4SdcgHZNFsG+NEo/ryLgBIZ4vWqahXIvaEp8hJj+NCuBTo5Im+4UAzNPE94t
h01PgBMqkJOEh5h3wBkGryx1SmNpGUnOmnHCSQxivvWIBvrAj9AzYWae0RPjpSmRjhKFgvQlBm5w
gVt2QW0WcbFNfhbtFtBPWLqvuflTj3cscnG9ueiv6qs7Z18X78D9xQjp5Qiil71NsmbDpJ79yXpw
bP6hEXziBIMBh8cMJ7oYh/CU20CKaUM31ZJ+NOwd0DL7kNMaK2jTHeBMTJWoBBdDIv54aXKqpU/2
PJxXGq0yw2fpkrCCWGQ/zYu5BLaQiFKJgntRlzGHiJ8m0W8dEeUvdVyocHUnRZ5z5xcNA+2EQekq
Dl1eFov7YA8GnZVUyGSyfw599+2bAvjEB99Tcs6EgZfWo3Q1clDxrYhxphgFjJxrJ7aSpKHk1zef
lXIXbJGYV6cy3v4tBAsdXeFm4/8zxrEiE5EDnHyq87Le4Wei459T/qLkK+ubQcIKSIsRmGzzTxYR
AVX9Ez5ZVzZyiLr3bzpkyA0b6fro34nes5gEz1LXlxzEaF9fUivh8VLhlq3huz8LEAhSKp+LC92T
pE+E2LfbFp+Ouf5FnDgcxsYRPUWSkUw4ExDYWun5bBUGiljsh7cmtes9MM36N5jbiADM1gZgFFG/
u/NfjLjde3sI2kmwmtDej12oUQuAZElYT/rWrZDxP+xhw2Wp5VG7gV5QJqV3EJanC9a9EvTLVDS1
5eUskRUkHpy7ptBQq9nq3AWM2r3dhqjNss4XMxF4XGGCKeOBn9RmPECyr53LLERqCX87YmJf73oX
zZ/PIsZ5Cc8WcXF8YYZlCtkunzU+N+fNT+Aou6axOamLfpqsmmZRqYGwWX91HLSrHgFg3kBODu+r
QAxGfk9t2XWR1o+MCiqjEDffAkLBW0L1qQwkPsRIFKyn5vFQA2hxw1gmQfq3wyeZSvssrpKgJyLA
Rng60rVTlphypQE67v35mHaORNeRJThTqRBifNkwoSC65ECHOm1u5JtzGSOZ/kG9lZyMJBl4PsLO
LiK+A66kdm9y0hoK0xhIHWADeEP0lMeW67SL8g8FEnAR292v8W6HBbzlWyIoWmOe3JCWN76BSLLD
wcRcI0DFnU2pB7/HuMC1Q6nG/WLJ4DL/Xtyl3KlzTVKpuAzRgpqgTJReut0nxGhcBrZwXZ4BbzdK
bDwCEO7AsZJCjeWTBad8dl2JyXya12F4rsBgelIEftnYXuvtwGV+KU3q27RYdp9/XGVX+T0OAQLw
RqnfHMPVnb6NRh9puZwP4+/RVSbmTNH+DvH+Uz8F8EJsw+EBG1e0I5S+epc1IURAr7sy7wfzfs6M
n1rV/9/956Dt7pwcJvmrAxyRujpj37LFDTfvWwB4oaiUE0wnCxvbtz+WRkZynRlxL3zcQcizvJs/
6KqfyF+nY6166cKfD4mkvlKYGQAzvdMnGcBi453rFOCDgF1xEjToqR69OMK9zbtbRH0O4XRKeQl6
Ax5CcwEs2pqjOEJ+V1ww1KC/nQ2PK9gLxfn5VLsM179KQDEuyN3tUMyfLgBHixXbbsIW86ZcZLty
N/yAK0jGfMPP4su8VRaYvgKKNnuFxMso02RKgBXctzLACiFakYWQw5oX5tCEPz9ImpFE9MyoQ7bk
1v8BIdzbxdO5b5q84Ta1wj3KovBp6aIuTb//gqVxtw9KZwzhOtBGM/WzDegfma5HxKgUMMlF1DgO
qdsTd3cnmG0Uts9JY8LWreKN2qs7PAkX6RLGrZ4mdZZsT6kTN6N8JcycUXna5YnOxBNoE+eXmA35
3cF/lMFPML8TMn3WGKIa77rUpSJvPyukDdYFCglHdREv3C/LqBIUeSPc3W+Fht9cpVPGv3bzZAWP
owoK0XnlsQiZABbspIDtpH5Ddlev5srPrdlaO6+btOUqTiJmgZlFo6ACD4/9JV3o5oKgBRyOjf6r
oaRXXE9kP9RTfi8us5cF7PE/jSCkNM8ZfA+J+uwi1SRhSwxQaVBTYDQnYU3t78O1cXIxezLuwgdm
NpZzFiylCVzfKKnHN9NmTCbUEkrEOHxcScyf2nCM2zl2mJ5ON+Q7jns4HbOVU3p5gSE2o2RB4zVF
QdfzGt9BX10wPBUWHACrwo0mpB2aZ763Do+jz16jqEN0DLBd+yWr65ZflClbEQ2lHSLgfDfyfK6H
GtSSYeCdwBwrxiRhvKwG9RkN4ndKJlwVUthB+TMVuNqgDoNVH/JN7lgRYCAZP5d2iXWwW/Yvre9K
o5T78sFghVXmTIQrBFU6fi2TbEeVxjTmYHWQMy5QF/AFYdt3cC/rLD8WAsvXCMEXDCI3JOS3JstJ
43Lb+f9QkeOt6SWpJzqGEu/gRzSNX6rObdajdwJNrq5fOJDjCCYZP31o/Sc26s4CC33kRk0uiY/Z
e8GY0o+aldz4/mCdZ9qWLyaCa6R/c42rh8hbQnKg6HE0Jg7cshrYqEM4tdbzFE2zOwWj54qXhpEV
EyVhsWaCZ1gjfswGSOciVckBHPM8Dw+t4W4CuPI1MSjV5qcvBrJTWix0fHzNnsj3QB4AbSmY64je
pVdL3pDyLR+yQ+n/o/zQheOSg8P5Jzd9HctiNO+Fs2XbyPOsglG+Kx5GmiI3Y9YDLntEaj3tYIfR
p4dQ+EEIsitD/fnyZzMFEIE2bXDkce7cso0XWVI8TjIwsOMsRE7CEYT4T8XJdnF4QPfgBAdi2Xni
S0UOYn29SVKVMHg+33sbD0UToDdFeFT1I702EbMxDdFYJWN3St1AMndGUUAWCKIARdhb1woWWLK0
GJ9188QRXPmHfVGICPGFsK2uxFeJF95GTfrrbUTaSeDhFJqCom8jn/WbH4vAY5kjxhllTJkASAd6
qG0x/9D73Ej351oTIFeJGAP00E13f8AFJzjMGkNVihv/+8p0r81ALdo+tnpiuU1NWdIhwSMrrn2e
lIQny+6vke0q2TtpL910MVUFUkdw1gqAB/Y2Tv5NvrbWGUwM+qU2VQqS1L0Dg7tDB1sxGQHcFzLb
/+QV2Pr3fD4/Xo2eKkxz0qk6nZHsVrhfFq8Nz1VPCzU0iE8AP2vvLsrlWhuQtCa6NCCSV39rmTKC
9S6lrKCz/9AU6G/ing0z3fUWjDgKApAgihgLmUlhXMa6yckHjQyKn5iBVwj9Ud3qEPYFcHCRVv95
+xNalQhMlkLIYeAQLvJNiEX0CALV5hWiMaP2eZA14Ph8j7Ui1bo+ZpRz9dxl9VO4SG7biDwGovK+
nZ0XNLvNOpQJuFC9viCO88v3hcREErKmOej0KIeGlsb0LLYHq4CTlxLvmO2W5fcrrs/vMr2w7mf+
FqrutKRx2JpgLHkhXTpJmJThdQkuImgwl0hfCJ8IoBm6a70NS3i0xf/gNZ8mq2+6O9QJ5pp8Xvs/
hHl0qxO01hxfyLsSodvCJbq0DplwUTyZimua84k1xlmbamxmlN/sTknYUd2NtmqM1S+j1KxJYBxC
iHSR5iga8/WBkTYn2qYcboENMWsaqfdUZOPjznMozAtthEYmHHIxkjQoWOzdlYCdN3MjGG6GoPYA
WOMAK406ClqAbuq+uVjfldccoPRdW6vo1Wu19LVr9RCizAO1ph229zw7siwRoOBke0xi5vC3H5Q0
sz8cHMrTfl4vv00ud5y0Fz7nOwlnyE58prZB8OW+e6tN5QZ2UFoG/ePaTNrw7qVtY+y5N+lWRzQd
0i6sSzftXTkwPC3nTbv4UbfIN5llcIk7hIfXOFUG/e6AhAcdTz6EYLfIDyRzLOO4jdjl2W7aYGlF
sgQsXegeFgNxsaITx75oZeAcIz0+1uAvST3EmoEqUqDBsnrVjYwJeXLQIofVqWo2acvfWmclGXAn
kN/QE4PpmgYyAOfUedijgKSMBlIud8Q79owbFIX9WWA0JI1cfCba4ss/c/2l3jEVQFTdRkGZJzJ2
9XHvtf8e1PC6ps9l5BCmEVitD13ZGBc7eS80yPscFfQeQCAbWSykgkbnTkk8mYJYtFA0BW5vrC0L
m9eX5uJr1Z4q5mv2Azfq9SPIPY74kF4POQCq1vitZorwsKKXNLvuXnI8LZtx/M2i6pxlzDWPaGvX
Z64QaS/99tORG1SGPeVXcD1Jmg8jOXzZdDw8RupGHONnHNvyrkZChCu4VQYKnSzbiCsE+6tRfX6G
/LM0M3h49UC/Jr0BG/4UaXtmQpjcwTVMTymbVSOesUgthzuYwfuTca7/m5VbENSQPgkpqjzpaRI/
ieEjq7ZIrymGwgYkcAdyz/XgWC00qyei8TxIyRISh+VOKd0ADtbLJ6Fw4yjtz2hiQd4w8oOkb0d8
CBjvwt4zIOTvppOpTG8EJj9qQQwBCptq/3Em8nuQnmykPQDxRaazd/aL+sKr2ut3zR/6xJUjeiX3
+hHtH4nX3VUMttAY2WlihaPlBvt14E1T9KzPNIUuabLY0ejGWTJM8hyaYzPXFEdAdlqvytJhknvl
2kjvnyfITiL4Zi7/VlVZ6crKHBhMJYCaRQnkjfLtQ5EaiautTTx6gGqk0+I4YoFgAagcXSX3xRYU
iTv/MfuHQWPHJxVtPNIt7Dx9nKwbRuy39AwjjP7nEzFpOJaQw3Bq0nu0+Q3Qaa7tRpm6glmqELFs
3NxOnBsy9vh2nP59bLUgdhXyOralbMKJDk1obxb9t5GS5G4xPwYkgfySJiHDysm7iAWJdYoV+Bnl
5y1qvGTVimH3fLQp/wOjTlrZlOfdOodVEUGmjWEE+Ibnn693VrkSQzh/ILcBw/XYoJf/xCRQKm/+
uINiaf0lgitm5p0TDZ1iJvYbvBqZKmG1xqlZgedfIkpUJyf72jTkFjWFEzXZpIlCSe1ZR7qAOqEZ
w4f3m73Oz7V/PrTLJWC0EH2d3L462pIUb/Oo+FpAFn5SNyYDoQ4CldrNEYIq2G2HYnbDfpG1UyE+
NSS4A3crQV6AZYc/kNmxch4/zwqbAbbmN9jaLX+T+qTZdBvoicmufVRcXcFR07UZyR8QpOO/as8k
SIjnyejucK2vAmbRls0ykt6FuiaHgDsa6RpnRkBV/5JWRUr51VQFSFzjsrU8/7IWzXqAKUTcKlLQ
lQFQB5ojknTdEByQP2f2fg/uOpDXPctm0NCGINGgHJz6fd3uLOu7D6WpShWH4s/tCg/xWCRS9HMW
KWKZvc7wOC1aXAWe05mFtDIqwJGL0KUyJNCfotEFQio3FvV1R8KhhyhD2PvFX7c5zAjH0DP1jqiD
wAjqpWVsUTedauCGTX2b7+X7xXSzqpwOvdo0FhTt82vtAD83K9xm0WvYkiKNNK0cBf4RfflDTdb5
mT11kO1OMS2aLv3w5l/d4x5Js+uTYhwHH4fgbh+Ubmcvnx/9XtJ+1TDH1koKR72HeQ5AVoFOoMva
+IrYnf3ld3SxdtTSYmJLuQC6xmevOoxLIA7Q5lezSCbL0lwIOpHLGi7tKa46BSNv4N5YzVQbNrKH
L8IVV2C8EMmvCYpbKRp9+mf4vX30WOb4Vy7n9c1KCtd3J/fNfY7JLE852uzY8v5CYKq+gSQ7+kvH
5bLcorERDdEjy1HtakIwjHAiN/qVKfhOh7U0EjmGnFll6EIsNH79fTjzo83U772jLolPqs4WOjK6
1RvtiYSt9/4LRiWF2OQOkbUTkRJAyRp4JxXdFQR49wLPzGN4fOQhQozx27/zYo/TnYDDWC4pJkn8
XUL/XC4UjCT/XCNBUfoT86M/Hpcp+O+KbkwHazI18LnTC1xqBIBkGrrIziTdWo2UFkLWkigYR+75
bnM07crvcrvqJP1CohzzVennP35nSelVf9zPgi8dPno9R2TZzD0XwMIi1usagQc56hfC2pPPzW1n
6mqZSWV8ckKkrXI3yM2Hp3VNPoluoMIyIxzz2+pTdiBfz0mUM+F+XstNVY9uX8jQ9Ez7CTNAPFBy
z7gdn/Dg1vBX/9noaWdwftUG7BzRHgqAYsepQT2Ei9oADuFKwHnuPT4erGbFLCyjdO1q20mytoPN
yywhRFnNlsVIlPQD8p6F+onE27pa//onbR2HPH4xSTk9NfZ+6Or7KgtMJtmWa6w3+jW8kvLY7fPu
lQ8sZBw2/L5xTK1O8scyJzSmdttHm74vNCGjbAvMhdKaOi+jh+n7PmyfyUKFjXc61fW18aRcBtNA
HUSeKW1QCAfxNCh+3fTLcEccCEAzuKZL2gUcqILyv6VVoybHOZU2NjjEzltVd9l9a6QXXs0hcNzl
ryoCyKV3byR56nwEa7zui8uAnEXvTuXDFQtGwjdQb4nrq+QMFg+pkp/nkKpAVuUBNB1qjfx2GjLW
/eBmYk/x1HKzATlJNaj+IEfEWIOo8d2Qptc9BC+Oyn6DOX7crppApsOPxxb6x9s0vHDJutfOC71w
I2f21q6Oy+P9+wyPtpRLViOQDOK7076wD0OcYWjvlh+FNZ4sqOA5Mzy7hXymousWsrbo6z/V4qon
rjthbtTzc+ebH4xD0UektV2cRMrPf49OwFt7UNkHycDKerVU0gsl0HpwuWdinxLP5B08oDUWxRNQ
WjxPCpPhlJ/8QklLEhRRdbhtk0121Ht8vTQv9WI+QwO8pETsLl1TQNqLKha6ClgrjlUnrwMzes1s
UxsJ3B59Moh74H583bMyogVq+Ki84emUEVTkXYJTsBtVBNdi/zlnWP4B3fnayO0DrkVRWUQEQvYw
hqOyaZQigLAVXBZeF9fN6UC8F6BFrNYTSluJA26UtvEk3+K0hAZs/CF9q1bkXJCJs5mMwWSbfSP7
YTlPvj2e/tQghIWDQLW2RNaP51yHvFnDdnKAM1iKdb7q58amD2PYG29DX7dbn5V4cLLXXLgIfghS
MpQLj87E5eTqYf/KgJLKOCCqEzVPezZBlJlvHKhvJ4aTJ1SZl3sCqH7ms+kQ4T4I1oAn0ethoVKR
NzZc+tzMKOd6vL0gCERuNx2UboeOtDQhozhj3/MDJHAqyWXUWVvb/tsR8Fr0U0/Yey3O2Kn+8HHd
InLUKMo0U5aSoHe0yD4tvU+FFbbt1MMNP6yjM8pjX5FzaqTKGb+iAXiEMXQsy3ms5OcMwJt1KV6w
pEcooHojMhgiZKmi64ahZESRZ5CjjU5Xi1JrrMhNouvm7UdHpjxBzOh213g8KyNe/cQIWcj82w5A
xUXGDvQbO1VRpg/IyQCQP042nKJhit0vplII9TGI2Xr2gHb3OfCDfkNTqL+pRcA/+qn9geHBgHue
OPFZkHeFfjJocNR+2NS4c3RgQWPhi4APVzr2VVTWf7Bith8GIzwVsskH8/yjV8HZAi3kY9CbRaxT
f38CE5Nsfr411p7RUTlO9/5XTxuSSRhJzHyYuuQwDzPVnKBqgpqXimdse01Oz18GMcWRB4Vujqb3
4rtu7B/VLeKPkYBKivKWHihy504JgNFK/1pUwIDh0A3mtfsy2LZxdbTFMRvvpbRNCATV5H1Aujge
IHLj4fqtRX1Ne7mP7BVkqTruibrkzMXIbrhjPj8hTy5ZKQehOTpvtF08pt94TGOOHwNz3w9J6ejT
CQAolV2NshWJ3wA1CAVS6EK1rRjE4UwRarWp/nb1kt9gayQtl0VeqCw7iJIawW+6o3XHqqtLSn8L
qiRw9XVuPcB3oNkKf2hUbvxoBcPeNFXVRuJqTu5Ti+DlwzRgU4L3GRqgzylnH5HE+4swtxw+RpFJ
P1YRqrLbPlpP3+HVDr91B+ynEF05ZY8WSuThbtgQnngDfMlWhYvkEa4LfAbMR0veaC0NYo+bH5B2
0iiNQUf/WS8dmTqjsYCgNZu3pXieUWUEkxKAmgWRrpPpmvxkZ8o/tVcGMHy4OpCUEu/GCy3WlVOQ
5k/1e6Q/j/YhPPjume32gI4t6A0akrTeRp4JXcBnWUlyLhXdr7N7wVXWoa/MmceOBgGNkMGE86Dp
ryu5+cKvUiZIULIcg0l4MrJIKX3w+P2gknwNH8py+XvRmntFiSZi5E6pnDHfLrovb2ydXfWa+GSf
ECOxb4VQH1uVhO0zySPsLeK5k8lRVnvQ9lafWhmEwqD75+XgNbjGwLzMPLxqtoIqDPX5JxErAIrO
qvnPoyIY/kbo5n5GLzDkJEcgz76KeILY7g0fp9iZchV4h+/x2Y69isGJ/PfLkEVxf82IXh9KOQHN
/6KC1LzRPg0sqMtAk72gU+juO+F8C+RPc1u9FKSK6Ky/QKlvqPZHIBs/q0l4P+f+dWIdjZ/xLj9d
UMnYtTQVtI33wuu/jYXghFF4KuSm3ukDgOHBS6MzldOegAd+EfA0XmAOf/5Yllc6JFR8rYqDmD46
SX/+A/581b6tNCgHQrvnG7s1Tgsn8tmGUkbk/Gqb+61OqdM2zYhvft58a3c9nJtvIm3HKnx2JzLt
LrO23R1ggHxA2vq3QYpRwcBHvZ+lK84S/k101uHUnb8yZWsncWZ7AloiTaLxpOfGwbLkz81XV3Qp
hQH5I/ljkc0N+zYFpQFbeF8k0gYx5mjneGfIWPU17xntaSmOK0ECwKp+8I3Txg0LT6HX87C9fMQK
ty1lvrKpKm2Ck9iXML4K+SHldw7CVEIWj5CYD7MgFHSguonzyPZVLMYXvmjkOn4Dkfs91MzffEXm
sCGIUCFiVR7LV4FsUx1MZIcNHquHq2LdErIKBvnjotn3DAR6fcaBnq8fdUCa1kjd8QJy7xagF4/4
QAE9Ja3ok+hyqca7DIOFSc3xD0IODUsCxTefzG8qbgfDY8M2L1JkeK8vFNKPiyFNg/a7WtyYVa3m
lqSwm4e3MUiV4yUXNyq/2LugBOd2AnEJnBnyq2B6F1lBwAGalgUchuJiTrO+EN4vRk8eD9WFxwII
KY3e6+BdT7Q1RH9q2TsDPOVOSwiF83WfwIp3/gPJMn2FZNlC/AM2p1+ChkpTZf14NWwY5tPEXxiJ
i7egqONM/DhGAOQ/Io7Qc8ltmWn6p5WhL3RuCYsXfUi7xCpZchlz1NEOeXmGBqtlmqCTYvHYVJgb
Vi9naI293wU5WvJMUGJXo18cSIIMNn7nV3EVZMdNbKZ6ia3k/3BEXbyoiP+UUryPtvd7PpTc42ON
OVedX6v+Z4VO/0UNmSwTG+dmOyQTOXppC36FsMh/cAdEhy83QXiqyOZWrPVln+9Ug10TI5pCVAQS
FBCbHMSstPlR0Pyao0vqMEIYdkwBSfIoSDt9LR9mbGuPah80EOsF+UZKExQfz9FX9Rjnz9xwojIQ
J5ZlD8Jkh9SwSEzP/1yKTVohcuA8dZIKLFDnskIzuyABE3b6LYP02sNuuRYBgfNromMgQO5ya/uJ
qPL90VCFRxUZaI2sy0/jJpneALMy6AzC8p2SPSTm1VtyuO042sJ3WuD/mEhW2PXUTVDZgOwfZ2O2
sFwLgDjM7f6oqHuZvrLELeKnaRTQ2mISa8V83Srxof8IP/u6u3pg7N4zW9Qvi0NqkLXepRn/hxqZ
hxcwnlnU2pK7DUpspqXb3Aatt5IGjtrINSNKl0yIhMo3e3VpuKNf1HBaAuYIv6exuv4cpB7q9WtH
SgldQBuk3AyMd7/+m2M1N6sZi6LbPPxW11W8wZpPnAT1ejq05VIN8WhpDF42AFJJ4wf8rMyWVuNt
7jPjj2KQoKdfxQ/hD0qlwMg5Zvop8uPE/tEPpb+6d7n4OibeSg/aPqtalNZn48VlqihvwBuv7LrQ
CfLTODSfxt14Gul1x4iY+cnlq9AfMJnDXzlKtpejSvCn/EfAgxaHAnQbQOdSE2n4Hgo3cSeu4YLT
SXYs/XJEyAghXF7AKeJrqTHE5hnWlnPli+TrUm1RxMut7/sXHXda7Qn+wa+ueY061emP5cElhZJ4
WxX9il+FE+ujkt+6Ubqus4YGDXv3iGFUnWWpWq6b1+WL4S/09ChV8uDlzGDCacH3nSlX5lJOqaz/
wQ2JoUp2xJ5g2ZzIVG++MYx6+zEIdb1Rb+llSt9SGPIR6MGi9qAb1Aswl6ezsuU5LDKEiuAUNkGr
LNe/dVEdEpYlXM4hEZh3vvK0XD+Yat5lOKiM9DBgJ7e7fdnsbcj1FOUD6pFoVofeTcad6Gbi0WRR
xFlLvxhN7ypz87RWt9AQmbocmHeNxiYzuwuwBGn3VA0wTkQWyFYNHMf7IUS1873/hsbi9P7IkxtL
pOpFAhCYpY3MgcoZq6Hi2Srz5AzD1TFTM0ZQcOy3oIk6m42WY+b8wXy5wseqtlgDZAV+yO9WKzKm
1RsN3Odlo+2bV9MY354zhpZNeZmItbmWeIBmP649RFskIGKx7oW4Gct5in4+6d7lIbzpI5YNfqvy
J2c7UxFu/ADWuG4J624gzcSwn8CFvgOtwSxP97OLJiBxF39QiLzcUjq1e8/vPehN9bYUq7XhCJUX
BQy0GkhpQ6NsYDTgOYQrAQqcl2AvWQt80sLML1u4qyJnjXHmUEHLEGwG42yYJcfcU74DS7og8r2L
O+un3/o3dHrkWbQOr3s0UPi9+IwSC3gRmfqdfRQWk8F5Lihfe95Qv8SUbRPJn+akU7FaK5mzBmN+
VQFcQ9oPDvjjI20MHxaGjwAmZ6YNsstotkdAIdw3WvFZrs3SIpv2rnIzqdeJvXjGwM/QklagZdTW
Hye5ZT6EoxjpT+r0Pwi9bO6cGpxu206KzxNp7l2TsMWWJF0l3UBIhOCG4258FSMLd21jKJi04OS/
7Da2R5Im+f8KCnzKN+8JFGlO/QZkSGlSUjf2tJftjkpbFdf1pUa2HIx07ghDjifkgcjpLjj9B/Z2
0hh9osd6CYPjVXlLcpIojqQnwPXH/5D4hbNGq0sDST6ucfVE1Vz8PIjL+GXJ1nFcrLKji1ouWp0T
fiAakpC5sEUgl/dATqxwSAIVjaoG2tDlzC5NHquvcZryX+gwuhqFYkdpcOHF+fndSmHfJW6236fP
XuTe8+av/1hwezGqCDyzB7uOuLVB2apinAMP1Aiwxxvk5L/5EakQj9P3BoW4WrWmuZdLhTEoW3Yi
QLPOJsxJVQ/C4xFOvHuy5AdghOmTUk2tJ6uKtOCVTLtQ0U+dt5gmfhoF1NUuZxRf296fpr/erByK
mg9je+8Uh4COA58sSJnzxR9NmRBFX5drlVVAlmr/f3c5CM9LuPZ7WjPsJFgXkG2fNc5TZf4XiBcX
gF8gMyu7Iti/YNoTvWKEEftWTMg/waJPc26naYsDNC8PfpKa1CQu1+DoLmY2QCG3vfsSiweWv/yJ
FGLR6rkn9zDH1owPBJYnFHeXGvUutFDgw2nb+W2J3V7mZ6qf8NbSn2/jXfBMWwGEtOupmn2bxpzk
7ssfifbzbi20u2sLwsu/2eWqC/LYso7gUpw3o+vB5g+y0ctB0o1YaExm3s6/BIM1ma1ddGWKEGci
Tmp3dggesY/3Pe5pYSDuS4VBXJQgCnzyhLkdf066DZBWLajB7/zP9BrOQWs4sRHUTWYK4TegyODT
8yv0x/ThnvISWMhUW7nRHwHsgciUV/HOq87e7ez6+aGjKsRi9IXqSV7IYS7WtiDk9KyP3eYLluot
EussHxELU55pF17KrXVRo2LXVTKNy5kdbFAkUARMZKwzkm7+/7Q/ElcoF7hGQfFF3RTWbBQdEKh0
OSr+o41ex7pGCJ7Nfb6RNpy3aCHbaR1kaTGG9v34pVGvX/DW2OW2OsQN0aBx78jqw17v/iOEuv47
XWVp8dYidiEaiEiCmyN11uz1oEt46hgc+RgZnDLlbO3t7mFaBMIWrBdD1Z4rk1LG4tP2jscN6c6F
OwMib+1QYJmI5j+h38WuExrPIYtPG1gXIpKsLO9eJVnRZLAbqEqMNJBvMtk+LCGJEBDN5MP2M3+H
sJshvKHmm7MXLbpsNF5gKwY37JlTkwbTsAskLVyiebB01nb6GGehfb6Z7ns7CA/JckxxtUIFFoB+
Run3n4N1GqrLp8Sr4j1EJIUkqVWgnTW14Jhnf8YyTFhJmMGDl0KrcVOH4vVEFr20nb0RHBGH8/gK
WTQNMa599RpyxBJntLz/90yCox2hje/VBNEnwgBrdLe5jDG5f4HEEEodJBlsxx9kMpiNft0WxN7A
CvaMGjBtqHz1+tY5YGL39cxyYARU+tY4tcyk2dTj1uxYLy9MkBeX44IAj6LLcZKtEtjArW/yzGz7
q9xzd6TPaC32o5JuTTyiDG0BirwsBuFUrUxgqfNFA5aMnAH4GIaeh/E3hdsTpiDaLDAyi1z/8jOX
83Ip8DuxUbWzs/FiYfOOM8ewBXz3ETcX5m1PhN3PXlfGsnmHTaixRNZZQIkVzNSRmj/soND3hcJ0
CiN/Qsv9GSk063+P8zS94iMb856Qwt9xPVjgQUtqkAqhi0xp5+hpDDjvA9YzAiLoGZhbDVJJTUbQ
c6zL4QvfgljGso3yJ7COaSyxMTz9yy0nxmHe7qmEbXY88yHu07N0SFv9I6NYuW5zMlhtCeG7C3GH
9ObdWjDtIeS+5n5Uc8gm781/DtV7gQev118qTAS7hMj8ncbmqUMez0K5jVcRHeQO+ZEJam2tSvxW
VV622HKQUIlt0lUwA9xt5Vt9VViTjfz+InmTBlmJZPGIsK6ocxZotc9EmBdm0m+IyX+Ih6hjz3Is
CKMjcy5bDm07bvMF9HTlQs0wzIvOfmyEe3GSy09DKwpGPutvezIFe120KtISfh0QaliB/kap9qec
ymYpU2ARd+t/AzfUllltWJ5w6dN6SQ+wCmvzg3zgY57LfVdBHBvmVWDv4gbbwonuhyAfhsj5n0pe
VTXBJhJdfN+niaypCbhJRJIMRrbo+/eCivc9K015DmdpJeDVueRDxZuFlT5WNlddEYI7j4YZIiiL
cD9vNe8iCMPbGP6V3CELJFbCELhY2XpaYqEAVCkYIZ/0g0vhYKSwccZAA57BlFGUYac+0sXw36gp
VJuhrDFOq+feYLs/r9hUBRgBr5cOgKsCX6kqsEBFAL5FTnb+glpQ2xVl/ugWHd3IH+V6yZG0i9vf
tDexUGWdTDwKViouITdKZ0FiMDOr0zmVlcnSx36ShGSs+47UGLZB8Wgl/QEckOwX49zPaXloxhq4
U4b7fmOJPQSmC884xM2Z1ORFXr61wc3i5ujkRqAHBOIIi3Q1GqctH06FA/WvufMApxkW7IhyaIsh
7IdmC4KJcoXdQulc2CWIAdoaykXQIIb7RNB/dJoajpRBYKMzyNAGWa7TnH/STEuJqMpaVP46o2hA
Ah8YTftUQwsYmbN31lJCE3cN1dTjxsp+Gc9Zi8vnkBjNW0/lJ36QWOkvH0/6lPA4WbtADsBjzV0i
rEUAWwtXM/hjnlPB7ugnVrGbWqqwLKZRhftOuEoeSbjwFxFrEV/GoprUaODzP+nn+L1DpDkZYmJG
OKWDY8yD7lX+Xl9fsdZDqbSxVlFG3WiaUgFW2/hcnWTCuFlYML+hDbb7Qwv3yd6C/RbcfBuKlR5s
AFe7OQJ7liLk2oM4j7VIc8B5r7Esej+ecaWCo/qv6O19gW7ZybWS6FGcXtuwqTdtaMjEXO9y2CP3
2rUUyh6ZLsjx6Sz/t8R+8zDlc4Z5KIj4N2IoguefCzHYMCroMZ+f+TRIi86EBPO0a47cztdW1/H2
Y5b0JJ/s+7y9V1nU/earXwP9QEx/28K60A2vRUC2lmji20cJ1bRddbskzXq5/RPsbK8kCKDbwQMM
phvFiIX955uaPxdsA5oPiITs2AfZkdMVFNOAhQ8bV2wz02kHzK17Eal6gc+IPEkBXW9VKZxRVhil
4DZMpnahGE9S4bcSmySrYQ77bsDZ0Fzk4ofe32VYBgNKh95pFcTN1qt1uuOZOmQ8wZfTpoPzx8P7
2mwslZsjBzFmgTrCe3GGNbqGH1ch8iJ7J+O2sLqtrAbSI4UCFVXE4mSofrmLk9fBpUaUFNXlVHZu
L2Jv6KKhe7ax9BVBHVIxScLbvR0JnkL/u+d3NeOQCUp8yRcNnLOa880nsZhhC17qzh73jsD85vZ2
YX8FKxbDALAgzAwmyZ0sA6jGhC5IRDe8OKglt12UsrlxclIAsj6l/ah0lH7lPU/1s7D5U5/S4Uf6
5/UDypDkwRgKbXk+sdidLHNcp5YhTaxKSEYQzGqt0v6RDf0HV8fNswYmKqNLvy2ofmNBz1VNCoEm
q0cGNhEDBc87g4V5bDQbdfIHsYB8boQEYeU2mBc8KOqbyLazBXozutK4XGfhKPm5n1D0JUHA1ITK
WtO7pyAx4mmvU4DIZ1iVGBHolKM1BfpWDaK0W8CeCIDEvfydwgFA/xE3KXmcGgGJaJVITfLhNH0t
XT49N9hvKyRETi7SVBcn0fyovFgEjhuE1GgsThHep2K3St+ByT8A5xPWuMWr/wc2pq6/C6Pl/By+
fZGruy929JHsx/+UYJ1nkdcVO0HTjzMjoF82auKYfQ65pO39xJQykHqwVly3exML7H6CLsbAk9eI
xCP5Gqfzd8nqEDArK1UPedAxxKDRCMs26ie5QsK8FOKXOGvHQ+loD5Y/2FXaasFGdIlMYKvYA5Sk
e9cNKfqjmTe6DAFxqkmu2ND6OVD1YZMKNSwItbIJ8BGAUbEsUKXHV77rZG3Pnb4vbaepW9VOi/NT
JfpjDm6LiNnme0DyWTlinZis5bw9QILuAeV2m9hV43QLqen8f4wYxBgEYtTYEKV+km2t48OzJurH
o7nP+H2msHAY7Du4n5IQk820chb3TBnVk0ynRTlWmrcet/1pP5ydP4ELP/3exm4lZa1h81O1BhhL
+nynxpsPJtmmjZcGcGWawpGXbeNVYsOlO+9532LxPG4R7bf+ogYPbNn1fZGcET6SQPWPojZDWVNM
xj5JuLZWEMWHkwOK7SF4Bo4kspDXyOd2lhAlPI4j9fRxj++/Y2BiCsj4BR/D1GKeXI5H6E+iX1Ch
8F3TEV71IXTS0wIado6J+MLriUehohMa2XymM9sST+A1nG0tMMonbHqvJkdVIDznv0No8Akt4wjF
ZUMv0HwhF/gUFyEGuUWC1knvxr4uIl7Gzs1oTelRsWYRTehNP6VPhU4gLY+bih2Eujg5aFeOQihP
roT8PSny5vcdRlqxqPtcWIWeFppr8u5DulsQLfowhIfMKRIBLgO9hTFP4lOxb3zl7SVw/YoIpMhI
Zac7IpHJsL5aFh+/x2ZFkT0qHWQ0Q5uwNfLtPJm7A9JXpvnBmndGApTY7zjDSdBkB4/7GWWOP0WV
xHLd3Sdr+TMf65WNRWgN4fu1QYBakUa4Jjz/pXqyima4woR6RhYyoRZbwliqMtjilM2WXFybHVoU
VLeTLrrl/Vhh8B0748TZcrlZ/U2XTzISXqGuKSPXqH9adoNwJ2Qku7Vo29st+EWFUM8U+rgfZ2wq
RjdQt7wplidSecnLNIJQI0UWe2LrLqlTqE748y0Mrtz4yTBWjfxUxl1vNLEj1fn5E8EBTc8sdpBm
MUJVWdBOBscbjMHTa37PW/sF47fespKrXuea4arfdt2d3HuLPiXiRfuY0q3C0nvbsem+g3ltX5fV
pMVR1YcsglZnLrrNA30+WuHwuT8I7FFMVxta00aP9iZtvrqQQQEXTsFexsHIjL+Ee1U83D4LNfFI
dithvcptDkvk8agRXwIiFYeSapX9q4Xd2KhEp6b5D5rgWOSJbVVbXEShGGA4ew+vY5RfpfWVVHot
EVTl9UdFGzCBT1X3bn8dG1tljesjGYdgedXlox9mLe9YyoIA2SjCZq3rhuxdrkBg6BN2nqUr+55r
/dsSzuIZdctxNFzrY8kNGRLve1UeieFyayVp1Ay42ZHdXbVUdhJtl9YA8YKs++kknxN4aujkPmVE
HcN44x3FCbdqnR2fK7tNT+l7BKQM4Jz2m8c+lmSVwoYGkZZqAQdepwjN1Cx7qHglHjqiUzdeJk5E
ahNg/OP7/llaznReY+Qo0CvcR930VSdZUgDcIjlH01js0kJntPvDp7IC4ZPdkXXKhoqgHeKgA8x9
A7Ck/YA/DrU4bdhjfhe8iXL7P7CMzENC1EFd976klvxeurHxgVb+eIYtAZGhoMdt95HviRMKfi3z
sZ4G+FezL82/Y0EuH5I/9rbtheboYFV5/2mTCQ+kjGE6geqYXBWeuLtupq3vxKCxhn0DLxt2/ovy
zwXo5dSuo+vN2K4JlHBvU3eGtc4t52WeYW/lng0Vo9ZGNc2G+qvcaj6l4d3yblqz9yOXtLYTHUbk
x4423e689CH1iRuk3as24Ykm0tWg8wwAFFYkCG/DozhcG9Qv21hlVIahUp1DfA+00R4FNQmPibpS
dNpLkj5JulCZzgfDMwiJx7OGUQjctsL+95aNVv0cQ2Yyc9FpZ9jvcTMwbLvYzJ+L3Jc4PzcOcoat
ejmqv3SqHJHXwU65+8gOyWXpMCuNOKIxJgeSGiPr7khhMBpH4+Lnx7Bklv8J9tK8ZRgZohyzWXXD
CG2Pp88/nZs7ZkSd4Otn45KjONAd4p/Kv3gaoF61/dMY07H71woljuYjcE+aWw4XgwIH70nbg8KH
3ZvGiXVNQBqmqEiTfLNKrAb3nUzPPhBo6EjBmJmE2HiDnLEA1F+KymkzygJe6/QgtytVrVaqC4ym
RuipKyZeGvchqvTlZ/RTCwsQO4o78xmg816L47h+1fw2sEG3GtLNZhl5FwyJzyvmvmkYB4EyL0HN
eJUiCLYPN4EQNrou7mbaL3z6dqvVFNYlit06+CMpWUwRIivnDf6VIawH0whjODBV9tMDiE01NCwA
0BT0yVznr3NfKxZfyvk0QQA3BSDN1Oiq2jsqivyrpcXlnYivYHQgoOEu9xLrEOJKDyht7aronpqM
vfMOEG8F2n9yCVkYrmTTIf1r2FHt7rdsBSLFP4ThX83+KbF+pI+NGeCipVhnttf7yUF6sKJNmUo5
f9nif805fmJ3LQEKR4JIaWDZg/S7li5a+OyEtSGw/lvMyRE11oW8FypvSf14wxTMIMyooGKr1dV6
xJdxNFYJYkbNNA5ub/8GdR65VaKZy1XJBmfBARV7dO0e7EmJ9Q0zZORUzfnXNEFn7L6fbza//ZtD
cJpCPFFcX+rHessE0XMQ1b4zLzh2jO4jtUzXVIOSrrUq7VfA+JME5iLBvtL9dosasZZUXcGtF7dw
1yUimmKQJou4v62v5N8A4teNydoCp0UzIKMEXVmWyulBCLlX8KtOmMW+5KpiR+DfTACVsBHEDw4C
2KYeWg0NJKvKdWu3/b2z/kOKhBlNn9vVYv0Mwl2vwvSrY+cFrwfsYubcPtLRo/fN3esEZMRBAQPR
DGN6u1Dj7h+d6mrRxliJj9VwmfXqsLmsJwSewLAhn+IJDTRauEuotPh3rQvhx1AOHJurgL0/bPZr
m6RDeNieM3LZKnnN2Hgc1r6Q9N3LrbFJxZGP06Nviwk9KE92Q66yQXW7EuFHK0j3l7MK2xBAiEPK
46ESxnMmditJy8Xo207LyluiUniXSXPSg1EvKN2Hn0n/JfiTvkJMp5SJVyw9tE+4kty994J64jSN
q1M0vJPjDAeoi90HgiEfYI73SHwDxK/YjsuhwHGDtlD7RxZ3e09qElUboklXvOQpx3mzPsKjgSEd
tJluWkSemK7PDuq++ILViXa6yarsH05MC+1bWMXqu3N4HzOwxLhe/PqL5IDxTU1LSPDULFj9C/bl
hYkRBcx0MxT52YvqgaeAMwLVKdf0XOureoDam811uI9up+vOJZNFfKVahBMQdJXh//Eiuf0J6dPf
IU7P68SjK+cu7t1q+YBJC1i/QZUNV8ZjAHNyFWjUvVtN5apVKd2cLff4Q/Oy+hR6y29BrxX/sQxX
F6GMu2tz8aN+16uBwUaSU8CrRinYKl+Ks9j+puasoZ/QznOSDddhEffV+kMPvgQ5BZAbEVMUGaoc
jN8UDmYOY4GTF1qyO/HFo+jHBdthXviz4aHI8lmDC3D5stTkbr90WgV6O6tppdesxljvqBnrX/sW
QoilsfwXPoYMLqYOIeE5j55Y1lOkmNdNeQ5Ku9RlmJBzZkh6p2Knbn4KYebjS1UUVQD8GOuGMNNF
lvk9qP963aXidM/VX8FfJJCVH1ASMhY4R//Ctc6VXS97LKr3wPpeOMbxZNPjudNlr0mDr1RwNs5P
wh21aG7p9oNhwAvpsGbvMZ+JeSlD0qTUQNYNIR9/4U9NSR+MBImHpvOrlCYdSIKuimmGYu1si3hl
/8XEyhWMw2T5MeZJvbzrvrFLxtr4OvTgHMyW6iXJVNTUQJxhHWZGzw2BG1mevUFiYe+w2SDJ9zuM
GN1Rn97DGx1yO2vvSiVYm5fdSfbDxj46I6anADYKeMASSnLaZy/D7kHiMgA0m2VAIlOMyqiNrYJx
vZhwRHg0azHx6PEkrvnorGvAuiFdscZ5blYu4SB1MS6e62IBGI1Gv2OBmlYed6x/2INsaIIiChaZ
lp35yc/gQa+rRJDTA3a8tr1cC09szKZDqGX1vMZzHNSqEy00MPH5Q5DfMcozsH9Mkh4I2oRam42u
jc30ACvFdgJD1UpGlvzX/HkMSUxf6UIlA6Oa9nC3ifaOTOu4fhgsJM0bGFliiRD/yPammV+/7ARf
i/cSffMTJMS/eA6xqAs+ATxv0Dqtl5DVCzCJNCONmpTRwt26lhQ9Kvj0URtOc+TV5i71t+7iZGUS
YeVcweizcMwq0ZtsflrBJCdqr4zFMwEf5/oJKOGdkbK+ueZU57ws1P1P1mJ+N9OaDt5bewi36Lw2
hOBwcbleooYe2QkJFpwdFhEOOLG80Jfr/H8ajFUBjO1D8eo+b3GwJFOM3SC5ZdJuEcm9YQ0t5t/f
2XzMxLTZAXvPU7R9mQOXJZqSeQ9QpOuXIWvtcilWhCkPFxHrUUu5uSJPy6Vzfd2iz9DzDB7FXn4j
4GX2PdOSdhAGUeCHLK+1YPOgHhbJzDx6LJG7XvAUC3ce0SBQI2BYjYkjr2Pw2YqxGuZKd3v9W2vp
WjxG2+9qepiHlXFuHr2i65AGRJdYuQfnfOOwb5x1FEXc0jVecnRxeF8ZL9gmB5hQOBcV/T45+av2
KmaZhjV0mBLrq6wNv49uKyeOpaMCP/Xk4w+EM2NkomZO38qYkDX6ZbQjzYF67u1L9u7yaIAjs2Ve
2qFMFuOGC8r0kEuT+eTeGi8INkatzYcrHfLnCKx1RRdrvsl9X/wMDnBvKm8TMRXdoRUPwrTNfNby
6qHbL0hlgQ51+xTvZAnmAOnoMX6/+rU8BtBfG+nSDFPfTCJMN5hy1AnB2zH1S8lLP0zEbh4XGE0K
LNw1dgBvYhL29JyAFzcVtMU4XCGvPfoxVxcAVxtmnCYAv40QhiAYimWPHTGAE+Hd+lZe2dOgr5kP
gMRSmQntDIk9R7KZCWSnqsumbzmtw9PDrVmm25hKLqjEPhgddYVMhNtbKpHDXMm4CTF/LtZoXMog
r08c
`protect end_protected
