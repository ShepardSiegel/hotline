`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XtQEU8PjLyUVnjx8lnwRm7BudxbUHkRbtdyDkwM/XfmnMhb/36UdOuMdbmYW9kAXUr7WGRFlAmtD
5PHWHRrvmA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LrsNZtXhwPUW1cev22bMoK6YemGDDOd7znmLTzqpBE/HV9oOFuzF9I7xbFrzbCHFwlVSg+JzgYw0
G/aopx7rNfg/EVRDrYZoAT4tsK4CgeJMF1YB67WR9GzFmDvD9/OKCZMIw6chNj1RFedUxKnFp2LA
iOzlNyZJSy31ZFDjM38=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WG4nqLNm7AjB+a0MIgvZqWCKRYavAN/VmCf7nsW7FVikhGTH7XYq7VZrmkPJ9QBiqLBCWEVSJqKy
kf1B4TnGeM3umACaMJyaJ5hrMq9TjpHFLLnTZLYZiRo+7NCQafX8RErqyrYrt8BgQAupAn/PWV0z
3Wl0lcCC84T2DmHCWbREuUPKr34bCYxmRzsYfpwwRYx2undilqlaUQeCSRv7NPuPtUCXU9S77Uru
2skDfmzs62SwRS878pHvzLroh9n+gb1kcRV8eKU0Zc6EEUov7X5OGoo9WZD4Ehf7apj+b3jG5eha
U3TNWP4ywROiU+LuGJVo6mjzZTKlfbY3UnYWgQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PS2Ee12ZJIyoK3Eb/a5pSDJr0aOidFE9K3++lHVYnLRs6KhIl0kMVwiRvwHSRBWRKBvbfVIVqUvG
95V7tSzBaopnhvox+PJDivjx5RqXFmoeeewyGeKfDClPc0FpkNwxwlCdV4kcdcKa7lD6s4sgmgvX
wVZj5DyfpV9czMSB7mI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TUTYuMyiakjGYNege4i4MidKG4QQRWosmxTUy6Il4UhRs8g/cVSLDcKRCdXhaHOcoWdkdVnawWMm
NbkZzSJbW/LVI+yzl776Mcu1TOnzkodMcE3dXtNIXBe1CqRlIIxmZKdc7vWa7+v9A6l/pphRBORh
/PYKv/B7E9Y+Emqe3Obpxo/0ByouHbqmY93fKat0r0Zi+EXiHIKd6P3/yPV/CSRJpFYyMlqVuqQN
IqqHKNWMI4QeMsuysF7EoLTSrPljaaMdmBthX9BSUskSlYZ1/Ubgy8qgBaYIq2TBxMxrg/ns15x4
5Es4nAjr4LHuUEZRzh7xUe0QKFOdah5Q7Z58Mg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 72352)
`protect data_block
Qn+RwRrXZY0hxuIPbhju0Odj8znitrw6iD1x99peIaVP0llGtyEqLnmg70Yn9Xsh2acfU8VkeYjr
3xrK9Ysi53oUvlF676Y3pUtzweyFSGQJp+topABFDboyHiTA7Gm8jRRS3/zNUtGoTDhKyJzkFOdq
GMUOIPh+MZ1KoN5LOP8ooyQ8YQQBBRvB3AAEYNKQzyjW56TPfVKSU1eKIuiKd44yAWJ2gBk3Fwje
BgYoL2zmCBZxhvZcRSbIEABJsU69iuwHl2gXJxxoc5vPfwTaSqYKFr5EoXVYaQhLWgCbew1FMqAT
liTAKLMybP5uM18PBb1XQrckuOgOoUlYhOnuBPNN4HtkiR3sZXMUaTFVEgUFfynfN0g488GbQykH
Muv0LZ1sHCh3dH9NAU03o/oNNFK8Jt5bZuVyrF8HHxphRhzRFZgzGFpP53nhg1Lh4yKAh2x7CYno
AhfNA0e1YkzLvy66ORSb8Xs1Y2xhS3WlnSzFDn7CNYuyH8ctdeXyAkHF4h7pFhOtaTalQm5ZkQ7u
m4Rj996j0wtr+s9pDo//fZo5rlmNk7ipWYltLv5mroZ1amQKsd6dbjx6wZ120MrL5ZKrNRhsAfLw
GD4Ow0FYDHJNBUO8Pv58wPiP2/PAwAI5UyolEAw4cbJGgZ9ZM4JFogS2jDcuBtrkQg3k1o2SJEDQ
MR1bN978lm56yQRN3fCfXs1049CvlDfZ6di8r2g9RB5xDwj42j+F2XXCb5m8u5m2JjrFk7nXmfZQ
0TKAQhQxLaPZVumpAWv/PRLA3MikfB5f8TBofClNu/P13yF+u6xSTYf/TM8ZdkBwgsGEvJYXav7q
zmis5JcFwzgKvP+LP3rfVAK6yn7sKEV/RY/NHu+2sf+DzZg/9Qqr+UWop9qfGLMBAaIA10uvYnvT
m4z2+0Rxkcn+MSYnKppsPBQrKvhB/tekSiuiGOlWuY94Edupqz2EO+Ke2sf133+4TfNDqHAw5EOQ
enbbJ3A/YWsTURI9M5h5m1D5/IZuvqf+EaFj9xPU2uaH+4o/ta5uGpeIM2KDBo4EjpeYANJe9ymK
MVfItvu4KDjLPmBw33MDFUKJlruDY88m+uXhSonNo+Y5tY/tV0GODXk67Fyr9uZ0tKU6GnjeLYHz
3OdltxhnSN4ojVNqFDcaLpOSzEJCRLUpgMUJLtOZgDU809PLgx7a2PNYZpDHdBmMEp/1rTcgz1nS
n2LiI0S9SrNoZeU483pCvaoyj8f+46qZUG6QBrSfNlifrcxKjR/nUPMGXaq4UDNRSd/5vY8CRBN2
XB0zoqSRVuFbQ0aStPngF9Zf2sTW5/FdG+AR51YIO1/XduKbht7CwrWs/QBMVLEEUHEMK72me4TI
+JK1q3PGyVS/e7Z56S38skdleRyue8aL/We1VWVt4j8btzzBZ3d74Za3R9Jjkesc4ai+3pMw0nqE
zerKvC1EcgbGexrpqzv/j3Do4WVX/kBscP8BPYV3PddtrYKiIYG6K/vqvk7nogvpTnM+JCJlc7Nj
CLorUl3xl9AGYa+QSN9cky0NdB+RO2z6utKQJ5dZvI6dVxkcMoSJ2kzEXzHidFKNhwRvgPnNouu8
V6//SoK1KvLLqk1LeXHtmL4a3U2TKziaILdPthrqIMW1qQJn7zL7gSixFrIJKCkDKe0J3ATEvsJw
0CvwEPd1GBPhRRoWcAH3j3w9n6K6IAIvIDw8V9zcz9PW3aDT+wNlAU6zWzgT77NGc2O77qXhZtte
ZIOIvaIniMpu1KjYC2OmXrXYQ33Lxb9e9tIQCV36ia+RHFBvHWTaSYbPZg08akE6Lf7aSl8prpbI
bLgqGvhSWDvbBJxvLna37QXVze5zrsumNxsK0+hb6hRtL3ld4Z6lkcdH24VXk6jEB+RjpJrbQVja
vX38/cONnR4YlUqXOsonFVjY8ye44unkMF2YvID/uKNHp79MOEp9WE4cxndF0ceaVZdDEZgP85Tn
oXUBzjOUSd1FJ0lug7pSXnr1YsqrPwq4OBCkv0VEMTj9wvjGUTSRXbdmNqIesp6u0dmOq2Xwk3la
cynl9CTaxZrp1BQJzBtyhPca9whYk87izhyk1f+DmH6vqcTSh8wqTHSQalRvK030mUI0pxuWt5tD
HcbW+54sNq7Ww996VSxFKLlluDXry2RN4WBcNM6hdhHvprA+CIJyJ9pnjCNA0Mh6aoNCEaRyOMsn
BcM+KWp5hC2jM2u2EKMDtr59p+sAFkkvt2zywLD7HgRC2rSJtVIKvk9EppnMyGMi/MCr44x89Iuo
L2SfavSabMbBgqdv9rjvNHT0YUQyHfiEf5YaTW7UAwpdx6ih2xyihAlQILtdR4hj+mo4QH3AEdJW
Zxh+b488xS/LwCQCxM5ugmUtoUg/dgTgzvtE/Cy8uGmCTwBfxce4EeJskf9zWVmJBq3u2c13QteL
W/2WvBj4WZxlMNUaxCfDe/d6eBBHP/JoKdi/53hLASFK8AGDKNCI/WTCu8G9dt3daZFgmmnXvmw7
6im9FE3nZsD7GA+0xpo3QSRbNqRyVebFHQ2F3iiPM4V12ACYcYnQmKLgsakjlE3f4GXOUjGNYvvc
gMmTAMeSMHIlo7vSERgLaA9GLxPvEiTI6+XZJ72DXXLXXbZawGlePOcox9xHPiq9V5mKnSrxhGSI
Fy5WV6JjR1y+yfsYY66+Xqe3LVFhx9w4Tdpr3E0KUprjwYZH5/gtDxacnXrefZF1vYEFmKJ1YO78
WOmDZTbyoKhfasi9wET4xnwgmt4XlE1XIccluBVHZWLdJAWBb36G/6g9kdU9q8O3ufEniWBdMUTR
vAfFzQt3sQxQOeMjm2Ts/Dl03eKNheovySQWwHoDZCBKWYpfEc/S/EsC8XuOFiGkXgNLaTceL2Gh
TA/ee/gGNYz/6lhFJEbOWwBXxDO2sAIWLJufkO5LYqK84goc8iDtJupnyTNBvPukkKmqNZL3lJkC
sPwSHV99g/Gy/hrMdcxWUoyJRL0+EGSphH6O7UhlmOE5tygKbpCVexxTT3A562IbWELnZ5MU0j/b
epEjilgfrG9DFyskGUax/rAVvfWXQSY+xWy1TOXqJeBx9Mn/XyA/z+JF6QX8JFfI1Y0246pz23S7
2JSdso3gDvsjg2EpPXXK8m+0fGo+Z/vTRuP091MkZRS6d4D2TPPem4Y5SiKn50N3U5qfZMBduuX4
NTp+ZnzExz6hORaBNiuDo0ZlwxV1W4BxEG6Y5BMfE3GqDz4wdKoZZd8hi/YJrJdLeCa6EefumHFV
/Q5narwz0AIfnr3TPx5PkiwGCWrS83mqjyUpgaVGmj+bQ9TlOfLiE+qSAkaLTvH9tXerw62hyrXZ
dadJPJgMZd6gTTXdbbvllVhw002sZ4IttoF2Q2lTdxeTeSd1COdMm6LhWilN6i1ZLZ1lbABgXYY2
TSUoiRQW1VN5TvlwvyGFTle6FdHbyy3IvkpcDroZ9T5DxyX0MsTPLuTA81mFW5sE3CCE/OushS5B
jHPJLDIjrSHNOfatbhw0xnRRJHQD4SfCIc5oeTVHI0RmfZyq0imeAFCWErtm9oYowwWCzRWVgctu
SR91/wLFFEKx270MEKidLHepZCz6eDbm1LgbAyzWa+WlKgLtghUkKv5tlG5ACI26kxZgHh+TCtFM
Cg4tKmSlYTauXKchlPmH8a7clBbB4rFewx6mqWsrYTFPDCGNBmNL7NheXwhm9Ck/SdjY+oPlonol
pbP+4ytPsdz3E4elaobc8ZHGb57eohc6c9JzK0nulrrZ30vfxKVI3KmyFKEHlE/04w+PlEpAQEMa
oH7Y122WrrvzGWjvUa+TW50DbLKap51t57QmI97NCRdmwC66hbtJBueY6rWdddnhzRK1i67lKTbX
nsBwJ2L/zPWIcBJF2Yex+pn+C6L5lauKuiL8NwX6fjT4klJDM1cbqeWb/NmOwcR2dpqQM/YQBNia
FllN+4zfLVSDp8ZMY9+2iku/nWT6dHJUs5xbUZ2x8s6H2a+EWj+ermXPJptLFGzNpWupNTnYQeHL
NO8lv4AxP+GJISkfqZ77E4dgyFycpDu8Q5OkP0sZCh0LCI6dV4kT7EiqOl4OMqy57H+9wO1b6m9W
Kkvaa8iH+nHD1GXsL8M9wmScMnGfXjacfNq5Imlr/9sLOY2P/ewre7qMVGulZDAere6wpyRvJqzM
0ZPbdRHnFfPaKGeJaeZq1+BplONjsKrHuwNuxHFGlFTvjPUiC+m3Iy59WZ2HglgLRoCsTpof1uSs
iwJLLDIjswCK5/6KWxOEnoEOMLoRI2kwseEcErk0VgSrryGR2iTDNAXXanf+ggExSJ3ICJsDa9Sp
971Y1/I4H0oyaC1q9++/nGCxsdvepbu5GBg2H2vw5vh8QlpJYFt1uvnCDGN3zpdRO1hRJJ6e+iXU
PK4l2087dNigYb4QA+Jn74hGP5zT4oLkYxAujE/NIDItACR4uEtmuw1YpcBXirghsOeXpXuvD0sm
z0iHVM8O4RBHF0am3DMBOed5OzZJqYLGTicXvo0Yv1hBqWwWrfwxkp5HRzLH/3TQEfX2cR9+mYvb
pZ9m/2CGQPE+cRnELq4xyHrx6Tcl5+2rmzq01Rl0t3KqZQpIi/r7tziWRF92QnMIFxqvFx0wJ2wA
zPMmXUf2eZeEa1zHbc+Chi46W5clyJDQRE7Q1aZY2zh9HJLuXRWXFHAe3sWtV8IeNjb1bn0wVLFk
uuurWhY/kXS7/yKG5ASw8pWx/tOnrDlv+3OZkCInE5ReZZXAlYmXw9/O4ExnEliV703IMWy2jIZY
V57T+VFY0PHCbOfOOmNPzGEPDUHL+GBw1hMNiQSgKuP55n/1APgzxSJgawG/xGVxtGS+dK1KwTRh
Xrwwcun1wVs44HLinzgqRCfuL0/m71nIdHTMM/FX8GsBFapT0G0K/SdLz9QxdVbjN3OdAxkEW7qt
KU588N6YfrKaB4p6z/1lNtQ4mHnNNqZWKpfLGpkwzHfyokFA44RDUMveT4WB/yFpc2xgGd6T/VCK
RHToyZEP5z2Ik6IJZE3r7p0Fc1T+kBOdcgkxtLlcrICkbF6YQUnSe1Zg6KlS2EPszqw9vF93/fs/
fjOmRRdIdiHCy40mu4jPthmYKlVk0aGvGZDY8gtOVaMhwjfJY2xgRCfb4/W7pJe1p443R7vMj9ac
axAYFpXOoCS8xRUQ5FTi1Wznr8Qtt+pXuc3SkYuQcH8mqDZCQvHF0mRCh0HIq6i5c21Q7IFX66Tm
1fHqLHd5zf7/+suzNFP+nAc+BAsxQIA+szAPTKpR9baFv3wZdy1IUXZaFntkUOYdhwKoipAoeR1+
uLx5JU/Mwe0d8mVuUG9HrO5PlmJ2flf7taDyWpu3YXA+Ed1HKVrSu8GKIHa3NfW7+W8mEdIr+GuO
zlIPyzYVKKjhzduQuNawIY5E2Ud6zo6MGUtQjXLttQG2T5B3AWBkyIykL9N6Vq3EXc0sjgikMKhV
WyBRCixBB28aJP0Yhb78jFSIMOclMAp1SzQKAuoZvyOVrhFtLa7fKyduBZGXul7Hj18eUve1vI/z
sycw+nQpjFqR/kJlIulgA6Of/v7y8JvzDI4JCAOeIPigznwSU1BDZFWNzhuMCXRn7lYd+OuRCbA+
BzUjlmV+/j04xyFHu7WdynZ5ON6ectd3CuYZL18vNxiCa813gsj3a9P+huO8AFlzXIuTonK023cH
STqkOeNtMjX7ZQfCs1c7EmC9N1d52Zo5VkjEOUU/wtlt42WU+7LJEDFXqhysFmw65b2zmS9/0K2W
f1vpXdtB23T3+7fwoNLuImI9yOrm+tcJ2t8ljGnDbo1vOxXPw7A48uusvcnSzzfKumI7rNH2273c
RBf4HuvVM6o/0gNLcvqUHa1iZJKtthwO+u0Q6bgP24kGrjyijy68lHW+nGNje90YibGk5xy8Olbi
DUPjp91duU/PVSw1Y8SWwqKOHLRKWt5hAl+yUN/IK8BT0tYR8yPbSclHJ4d2jIQJz4WwQB4POpzi
fxEVzHS1sMTgBQPJy9kdHHwvsCOO8VE1aQtGOma0Rhl5NZc7VTHceFnxBc2bq4R/WZQlA0Irq9R5
l5uDV4CKs6Cayn6quw7vcNQHtCa58Ly+cgrRhIknHVWgY6a81DE0inHzaHy63aNYXtfLxGDt7lw/
z4Cl23w9pisKnr2Z68+WgAKtkFwE+8hR1SY/jQtmKTdf2Hu1+Z42HZqmEDp7Ea8G0m/aXDajfNL+
nPr5vpsbJ4JgN3jxhhyrggy6u2PmH+zKBzITmMPdqaLnv78t2eNbkjDxIGs49RERuMg2Rzylz1xO
vYp7UDvPbNHVpBoH1Elrjc//HvpjPxLraSXWJfc7IwLO57/aq5Sg+rmLkPwmpe9xsK1OJqxPlZcP
elz9Tea0yg6T02UFBWtJ7MnYarYzZ2jjLD5X9yN+qKWS4EgVgVHvd+iTaJqxEaocjEeC1ibZtB0q
IbAjeAJWO/ujIQRZFMqnAy0l5PKTAenO409W6/FnoiO2RiVmeLw3wNNA9UD0eSquOGGzBp+PuX1y
4i6JQdiBmmR+1BXxKo0SjBmcW9cFrXjhm4i58sQ+1fYiQ/32OGd46BQ6Ns2u6FeW3i0Xk69XCe7p
qEWmdyN2+i0GpVotunYWK2umUKPWbEf8vpg2u4DFkLB03aStuCAh/B0NXRfd3JUzyUhk3eT9K+sB
rJjIXULxhmR2IZ5aIxAzzbLI82Z/pTQMnkMNYLKCvxpqYDQmXJEnggFeaEihnT7aLtWlSlsfuJX6
FVTDuixbZ2ifpOawkzRAWz3+yWeqgfutyeTWMI31kwB8OhLJSibEvCrmJFUM53wIsK7hJpQwgsvB
xPLCNX1Ws7qR+IM9gyV6D14P0RQ2n+diXyuw7vlUtF7ntuXS5BG/k5pkEew35xscwmZIg5w3V0JX
MC90HQojV/mB3yQKaHBIOfnihymBmT9Y3ONRq0kA1ES+BshCL0pyp8h6ZcuYeNQ6fufjpC00Ht+A
XGjGHcMcmDd1xRf7R70VRejfhv5ccx1EG+KzCRalF5wk0f3doS7wcHntMDE8CagO6EzXSH8KGzVz
7h2/Jof7FmnvHPrabPoRLzQauTuG85ipgoISZzqMsrBv75ckz7RaJGCswAn/uzIi9lknB6/cypTm
NyCd4DY0v7lZ9VSSA8FJTXAuNzef+mPrAVBIlrlS/E5BgG9mUm9Q4DmkglVuybHSm1FIjq36uM+T
oXezOVOPr6dISnDUVcBI3MkBB2QeWdxXPLmKknX4GbYmLpu6kwnxE24d23Xn2gwq/znTKaxyH0Wd
D3nSNeU6B/UzQOuvvgEzVnsW/EILkB77MjPyAKQK2tAidZQtfhMFjiEsyPRCiAebQicdUNq3bO0X
YxybG7LpozH1R11oy/jJbl8uQNI4lmLhlu4y7ZXXEKSFNmXOLV+vxULyA5Z4fkN50BQdWJtW4Ckv
f22Y6+cYKyc5GkGpUHPwqEHhhOkd1HJ8g/2vCqCEdrsPBWe4QmSLHuxiQrK9LTkhiWq8T/LNPu7v
5I0MJY3eEePdzZl6ZIbQEn4huOijOYKYfgU6UuhBqz0zSBr36jC8pnqc1megmLMgot8MUxz56UHm
GUnr6IoHqJE9F4EGY+74lPM0QFiuzZ57L5R8aHuRQMYIJFFal4LS6XtkKNpP0EqHOi3m8j7os8DV
ZdKyvTL1b5WCFLVzSJ1SemxlT2fFilJ1cSAZOKqCAwL0sLYLurAmmE0Z7ab8RL8Kd2Ad56Zd5S/W
aPsUBusA+xz8unn1Z3Fhg+QcJgJ1iE2nahrWdCItePq92duhCZHVepXjlpUIwp3a7jzTrHivqpHP
WmTwq5q1cGi8B5KC9w/2z/B4jgDDufA6yFJQtVrxLm6uDXYQovOSoG4LWJ2zovNmuScV5g3nra3u
f+oMJcF1Th4EVT7U5S1a5Ct4eyOh8TLADO0lZdvb3+7vAuQzjQsQIGqQuUf9EhOX8SDXLJfklyEj
1wfkBfMXoQ9e/40znhQ6F31DSSrSwHXwfhyAbQbk8O7XWjiUPxHeOuG2CjSgb5jJlKa8lShOXCL8
rZczcwqeUTtOzKK02ZSI0STSfdmya64ZZCpzOZ72nTpIt8osN2sLSyf2GP33BA+iHyXfD4AerYIu
2w+QFDRlefzVCjjQi6jPcI4EwHwqyTNUotsSqhzP5xYVE6wgXbrgQI3pg4PYZnnk1X0OxxqtCu50
BwFsym+4qgX20CqXoAxQq1rvb5lsqfvfkwoFvncOqI9yOWN1G7Tc+qpB1wTo7S56UhszPdjgnv7g
iGfbf6mcN1D004kgmgAXydKCXLmtfBsHd6VHw+217rH9C7y3gJOfRC3RsWj3d9s9OdEU49hyg9Qq
Zs5DBhkgNrs0GY7ift95py6w83dw00r4Z902M27bh7vHL1zHe0ch9k6SucWtjVZ9Ke0qL/D9k7xc
AzLhXtqqLE8O0HfurqemK/UDQS4deIFV2UZLUpuNj1oxJ7Xmf3UTZx3Zze0gNtrPLZZ0mXUegHNi
BKGMIp3t20dm5BK3RmlVPygW5VqwFKPB5M+gTSH6lDAmQFvg+Cyc9Xrhv1IPqlfOqoQ0TxgeqVf3
ezAhT8HJ1oHBqL7yCs7llAl0/6yE2nul2Aly0sqYozhIkMl0o7D4GHPi9PWUfa3F3hhId07OYT/7
s0298bgbQLU7B8m0Qd+nwCVXOq4O6L5MrRKHeR2qHzue2ghNIrRUdOIF4r6jU2GutOQderkzPb8C
BL8wNzgk5pFyb7EM6TZ3lB5NGoSFZVHUbZwW/UB/MSn202ezWjuyNwVlJxiSQbWau6H2MuGfAXz/
iQo/PgLcGnyBDNLx/ufVgXvWNHqjYgZvY4ozk3VMOfvvZCfyHf95KPOOr9F3+MWX6TAjN2V1uBDm
Rm1itN52yD4FhLIVQEY2/PvnSbTKEnDZ867DmLANWi4PBohTSI06r4ZQy0yOgIkK3G7Amj0I3iR+
FS5j1+gf/EgSzuJRzpcEn1uD1ubIaWnFr1SpXPWGi0a2IOBNrZtV3iKZwIrp2DrBYkDbGLIsZ+Cx
TKNepvh/T71hQXTe8egXmejBiWFsgcCQyA2DMlJ4q3z+qG7hvmmk7aTdJiyzhQ+NauZF9nmppdsh
I6OPSuPG5lGXNHETjFU5+ZX2jPMzz+HIpHUEAzogPbRPElm4kOwuLwvEmDbbQqyCiYoWGA6mCX8Y
nce2rJFvTQU0EIh3WVJ8ekDL14BKuECi14oWXNi2Gs4cRMgwuLlFrDg6Ua0314NWnyeP64aJ8Li9
tMakej4xwtnilozRaKD9yffgK1HhfX84mTbB6D0UQRkv25kf9RB5dEeeSKXZfFvNV+doOeIDyiWT
AbF6kPWjaN9D7QxBD6bsxwOAwjQ9nImqtcDT64lnXeIQa+MQ242Q4SOFL9a/qSVoqYeXsOWGQtPy
MFEPIMm2ikB0K08y+kXi+sgDHbHRHgodkcIP6YsFk6k4iG+fjrMA0b4Z5uSmuUmP1Lt2XHPv5zwK
r82fZR6sZmGOCPp3pJwUYkiERXn1tYWKEk1M/o1h4BAG42v0CRPUxQlZuEVHNKo09WVB9hDNkziS
DcGpy29/UNdArqQwsRPw6nbaMBJC3QkPHRT0TP7ygP/HV3IphId+WlIFuf8Zbl8He6LXwS8HKKWv
pwFt3h7nyTm/ZW9H5ZdHYdwDXmzxuj+sDA/qCbaY8ObBI9TFAkaKv899iKgwKVEl6EbxRQ9SynPm
dApfLHqk1ygSAC3ap7uptUzgdw9daQHYA6C9edPPQPv8QPUPiGCE/+yl57qAYnRWorxpF+v2J68W
+VOjkvh4A5d0atruE4iP4+r3fjGF/q1k82aH4mCPXEjADL51/NcF42Oiao+oj0H2RKWOGBKIDmrG
UjyftBgVhNVTE2KHu0GXL0RqZAA8qVYuHvcgQZ+XJVi/IfVPrbaUfz/uaNUxLiJL85D+Ol01yz1C
TFX+v3KjukQrjBMFEnbhSpDh1jXcmblj2UaWcqml/lRuclB/Xczl15DlxZ4wjvNoO36Y6Vgs6MwL
lu00/RF0rxzoTMmO6alx0CuYsMgeELoLpLdIfx5NaAicScQkZP/IMLwqUm1zplujSYTUHX1xzqI8
2kpGrSg1SuQiGVbNTf68DMGwn/J7/PaKdsDT19eX0T1Ya0CAUk2Pb7uVTDk4Lwi2rHPDR1Wdvp9D
tTIqINKULbAqMDp1KlUEUHa6tL62jMrniwu0R66/mpfgK1Pq+vRtqqVBn/OjEstZ6Mq7cBasyWgv
mKuWc8Np2sbk3iOJ86MN8CFTnJXPKP3bN2lgJY2OVwz8M075lSH2YZaUqfkaX2p2/SuqE0KrxR16
RQDBatR8DHeGFV+3iZd49HS4KXMFSrzdfIixryRA0orqB/PapjNqw2gwievjR6LTqDbs1eJz0/FM
xudthOBH5yRoq0eMF+Rsbf+/5TczXBlNmSTDlsjJlYVoOruWBW0Sdap9KsSSvsiAjFDlbrQWQeQh
f7+1F15DqdgTIrqldcVrWzGXHLpnRWs3ZBAM+F355mEBpGNkaSrR1ALDJ2NsJMYL4FcWEvW+qsS+
0vzlz8FnD7u2lVdZy5Qt+e1SPJwCDaSTbJUocO1MurKKHQI4gu/NfKz+NrIuJJD1AKd/Wx+wrK6C
o9s9+ixvLWS/qsuP2qm2Z7Urp5bhbez3BSkQ8HlzDv5i4L10dy3Db+osoP+wxrEPY8f3sskYNPGe
kl/v61t7vkudOBE67hhnpxRHJKmetu8OwppvQrLjwn42Kkb1k+ccQEFJbXInrw1U6goWwxdrwcx+
n4i12L5tLJUzt11ErV0erlaW1Qi+IBqgYOzqBzSCwOl4NfSbeDcMijvpSsXuDGqY1C1nVXIAcNAV
wGyIuXefNZXsfjf1UtGOTAiR4BeIuJ9kof3VvWW/m1z5RhLrhqvzigLxhw2dYL8meuvj/SwxDZe9
GFIX/oOroHE+uhdwZbuhrVhbZVdT+qDtAGxJ8gfiqGkl1L33EgoY66LmX3B6VzMK/qBwCA1QZ4k/
Zf59ozggx2JqbGUrpBPvaA0S3kwk79altrB1U2OWWL5brf034RKiurBmrHMHtIda+GpMTpFyRaBO
qb3sl+DMQKAAnM3DXwqaxexXuMOspqAfLNmpV76agy3//+tHpc9MklXCiEz9IIHMWnF+ZzqSutCu
sbK8au/clYiN9RKvHFuv3wWnJFKHCJWskQ0HNGxq1F74C5JCdoFpzqE6bdGxAsbvszuK/Oi5ZRJj
AwZBhRFZ2gW1kr/ry7cN0Au95o4pVjffmcfpdOqI8wts+bNFlYc7hH2ILx3KrspUCpfewdNteNGr
JFxBJOu+ueZlVX+9qyECpYGR8FqGTnaV0JLSCMBhomv53A1C8wQZmnZ7Czo2q/A1iwWTG9xb2Lpj
xWtoV2f/CQRj4p+uxQVJl783S7E10n17lXZ4bAxvKpMDtZS5b0dPkVyWUA3N0ZkJAAGl/If2bDu5
VkNdMKXmPE4VOqn77lq+kw3BZQzCKk73H0bGamkw6KWdDn/HCCiQNUJp9NYDKct+Y+zU+kZcPRlP
8SywyRUNyVpAapY8t9rxjlqPbKmAho6K7Gu75n1GTuRuigXiFirNMMu/BQR2RxnIy6NfRrnCdm1j
TUPTlBgvqk45n0kA2b9/LVe7UH+2h1e293eThArADPJdIhgfAZmADOPeBvbbCOsatwrOhi8yeiWj
eL/podIWHPS9t/b6F+yN7h0IrSa5qKwrazHXAQM9Vhif1a60k3uZgnf4DIdEfPxVjwxmGLq7Rqn0
PIt+1rH9MWjqj6+CT9tu5CXWgz/QpWlUt9lpu4klbVU54oWGrx7JcVOuMjly8PrjMc3jXHdouGyT
9yqjYmz1JUPA6hghlKGXWF+Co94qNEaPHSUNjWdepnobspT57UqOi9LCGahWc8JAtpGSm1NogUnR
gEDrowJLxXzC2528J4jjq24w/CGtMUjrf0lXQQewiJde6JINkIcQhui4ksVSPq96Ns6QoSM3fm0l
+Da+24jp9NcbvH8B5qowhZg4lSXhM0LRUiXcXBGTwCyWbePo8dr8+WrmPgQp9XVabr0gDpVla8Km
ydmbE3wXfY4cfGUme2sw0chQp0UGPMBuvDmv1GuwLa6dnZcoqHBDvIxM/javC9IByIKzw3JDVDDd
l6pqsqqVoKLqneZxOh8iq2eLI91XKdv6z/5s3UjA4AJ62qBjGFAEAvYxoH0m6hCC21EZQ4t85ep/
dGyzKGZ36b+TBelKqnt4CLmQBLPiyPWH6pgsAr3cAko0us8LR173EcJEEbm2XmKvfMIZ6Wge305K
AdRW7XTGkgVfXs6uJ+vE+JQKK/D0mK+a1+0plztPB67rbfl1W1xWw+v1S2zCJbVvuimFPhUZnzIa
o8sfbHu5/V/wWhytTb4TVkGKEdmpy7tG0wxrofJ+6t5qKIrqeZj24wE3T56V5yo3+rWWZxtg5FUe
ADNsIJVEqreXgGFaSGddKgTcPT2JdZP3gDqo4OAmmTD3in7pPrelI8XacSmPDtilyhH45sIQx1zS
Fw1fEGVVBkDW92oxKjp9zEL4GSWbGQ4nlhew7hGgEjxOJERZ3+jUCbuCKaH4c5/a6PcGWEkLBcGf
5EIUk2z6EWfGMvjP6VB/60a92sHdIl+iOrneWpa4SaSek6jrDYdMLpvpkMrr0ZB0DGSEH8wYUx10
iruRszgPkAfGQbmwPwp4DTXx4SmiZ+KQjIdgWGSwrHFca1K1pbsHSz8if322vmx7wRqrleoypIOD
4mnoypXjmEpytIzU3GvX8OARS3u1KEZjYDGE6V531EcpBudKzn5sVdtUjxe1wWTGSllkwicdzpsf
QEjM9JlLCCZyFf1NqT1zSIBOFVlAul49WaXLyEkYX7fuxWa9y303cPZHAbrfDvdJsIF+Z5f6SSix
rIa2jTMGbTQ9pSJSEyFTgeUGo1nTTwLaSTE2O51xUJAGsUBCgQDxHwLla0tCfY4APwumsJO18lO6
KrkmQ5gkdMJ5jPO3Sp6k4mV+7zUn9igphbLHv5qSx8AA4LZkgTXJ4fT/nOH1qkxGFU3SIbNcHHBk
ag2JuNel4n+jwRZM1X18Kln8TCZCTqIIdm6AktqOLIHGDs4weiSOU52hhvLNdRz9vddmAlfh6RyO
EDYbq47cF0MFYujX4a3VGA3RhUVmmgqepWSbqI3ZWuFQFKpT5MlMj9uDpGB5k8TAdULrqoxBVBhE
yI6sLTT1aY9srpmf+QtzvhqJEgfgcz7moPi0Pb45voomjML12f4oCutFQ4t7SIczQ7S2axK63cxj
QAPyO5PGXmbPFKI14jniK34owgzcjcWq7c50ymLESieifT2RkB3Wh2UGc8zWc0mEHDEuQx9yKuf8
ONJ/Z4hlRCjO9zXbDPlXQPISe8JDSqYF3/lXNcsP4c6QkZPNc0pJ1jwQW0xE0lc0caTT4+3+8yyo
b6hwWETT0YY+a8DxSs0PiLl76/uQn+6xo3j+a6zvcWu/RrFFyC3t8NQpjoAQStmnGx50VaXasBFG
M1PMh8xersI2s3sc2OMVAaMDWxywZeHmEPtlla4oOJnGyL7w+1ywSQYNGapxc0bkOakC4TneoCDw
lOZ/2HSODyChPSUAzhcd3TLBhxWs0HBO6ip98ofWrnqi6vYizWyiJesnyQ1xF4yecvEdMvXyLCIk
vjiMN1+WOvrFCzEnt+aE9QR2RsITkWLvYCO7b5/qN2b10spu8E6qOE3RJDvh003pMcpKIu4Pt8qt
BGxXAH543d0zV2uH23LwkSmj20px7YSK/hicgr+ca7PKR9Y0mgCuBT7THI4POekP5dCQETKeRcES
NuqQKEe/a5/xmYfAOQOUi8DiOBD2FDtdX0a35JYHtO9oH8FFpRJxmEOAricjdxqANRkLDmR7AG+s
A8ZxvxpvqncVugt2/maB9XPxoaw1sEyJWGhmDYskVgEGesvCClhJbYoD9t6DgOUJgP8NygaKUC4G
uRs+CPe2XHCBcNsCX2pd0ntdd1DXCeBhqUmUQ/37sbN4zJ4D1GXuWLskQSLTB5Awak1PVVkkIQyB
/+3M2k+hURuu62QeurdqMDW4tmMkadURdeSmXyb5MvFmBSbOMEvHj7Zz7B+2+pvaKtnCHgY0fsTt
ucypqIg206gxWfzFJyJJ+mQ6R0H4KnbKQkfsQRXhxvQ1mzD26V8ATFMIWECgBhuLdErkOigJabzs
RR3C2BXVP6v5MQOcejwns69oz3GWbyfVagOtDqirQ5ReVKgJDe2EdrEIUoyaGjYz/5Re1lzIM+mB
VvGov8c4uCSDxAiidOWRqqY/QE0eNCo60u7Q6MoPxDltSUa7dHkAlbHCKC5BLYzbMg/Xy0v3vTyd
T9LHCimw2vLwOf+lhOKkJfy9RHLXODdKr+GLGODWlZOxC0RwzMyrQY43rpCUD7nQn65fjd7N2EvM
4A61PwxjANZ9c2EPjfhWyJdlHf3yV58L+UmWHFhf+vTmOXKJHaoXO1i9B2PmTLKmOloKjWe7jlCl
mwpElQglqeyDp/MSU5i7oI1i/C64iSdnGQ+aKIvp6/+uGNRfB88mB5s3D1godjg40T0/JlZehfG3
tflUJXhcrFvxMYfKytklRLlDD2iMojD19JyQePYEDw6oLHkLnPom1lReOt8B/GCCZheO/YKR8WEc
xzeICZhesLnSI3AdE1l3agiX4snL/s1Ju4W3Q+Js/ppVQANEkl9JH7h7bSxaavvIuFciYuPjvFLl
rdrjOe+i2nVW6VO+qNnRyVJzDGZ+XRZTqc/vi4I9Kwr9OV1dETsjbDYb3KC3OiIzo6j9VHPVbRMZ
JafIfais2PGm9sQSyC3aTqYILf83GSTynK52uHwLNRXmCFkBmh88vlcElvaaIpYuhjJeJTNAmdgk
58LMRudh9HVDSgdoIhIOd4unGTmPOtc0CiXDzSwhE5eV/yUJWpa0XhHvgcGg64aU1mEH9DArjNZR
HXtXATiNrEqeZJ0QEmanRAqCxAYodwJN+XX9l3cEpu/daKwPX3o4CgCHqD5zTau/ojcCACym4Fs5
TKF+N3tdyZY9eT4sWOzRcyizmhT8TKNM+n44nPtfA4HaUSADyd4KXqS4y0zq1gbPly0p90Rgb41W
5HGdwpic1NSR/zFL4Kv0k/n645iXnHUIqEoCnI7bqTukvk7E28VqLWGZCO+D2shdraN0UlGBQWL/
ttnD1Qs1ddAyqBI3Bw+gDGubCAyADUlpPGsD1+qSHZujOObhDoPaOtuB/QtEn2pdd7MWvDEw0zws
4+avZx/fzQcRPLtac3EW3thWkcaAxv4utOeAoLEp6k3bZ1+NoEO4TSQGFmH1HmsPwSTP2XArybHs
+Mb0AN4fpp8jYIW0473CcwjLpqUQdDQTFvLX+34a5jPeaGqDDp5afrBm5eaX6s6xD9FUBPQQaPzB
JHzuKCu/mKUrLdXHk5jdtHQrlPUrtHXzHyphWluLmw3ZDYrqBo/8TzUe51w7JUFNtynEQRYonrGY
3vsAWGa7xlrst4iWuWz09jC3bOyBfu5aDPEuq4VbkRgj5TraHcYbJ/Ha7mKvap4Gx4G0ttCFqVRR
T4Z4NTSmU5ITkSW2WBSEuA+MsQHwIWepYnC1640fbGgf8RTTygQvlHPU/xabOSCH1mkWJ6gun3TO
9DZlVUQJnaE+mZQT3aSBho3kTR7+U1ShiVPfCG+9wOYpg4M6GnZDYo/qQpeMIk/RKkUdRXaEvzJZ
8pAgLiS7RL6KNH9TFkoGeNM7a2vKD1/4KuUcIam2U89GqG5+Jj5/wVNW+ujyr0hMeC3i0+KyMYTB
VOzvObz4nfz5b+s28ODReZZghk33Rd5QHSSk7rlKAFz37ITnMyI14Zq1nozVXnz0iWuMgNd7AaRV
DH3ibmm34MVDd5iP3OEZ789w8cJJmJ6QY6V69XONfOIMM9nlpoZr+FjGj0/0ieoMHd4td/S9S5k5
dHhlbSJQAsPK6iphmVl5RTF+9PH9oc9vtznhlOnnfj9+AZwL+LbXlm5FTfa5j/VpsRoZpZ/+3DCf
AfF9ervLXfqEYHFu6IxLRsGT4ZCYj1xU5xMm3rJQ6LsEJNZgNnvg/dVb59fMWOqDTvnlyBghb2Kj
mplplMIqRUBMcioSBdf2GjimawHsWlL6utT2lvGH8J20axxs1yxUaLOV5HzgR+OiKyCG0xZsnHrU
4jZDxW0V+7Th2p74HLproh9utYRfOzf+LYFoHZQ1wUjmJxOxHQZkIR7E9JP7+/LTJn+t2Y1zl18t
+ILEWl5Uf838UzCUjpuNwuM3VujXk/I2SmSHR8ZHhlmZu6ORxpsofNoA+NGifV6Ci2ZwvRMOB4Y8
qs9xN3q5gkPG/h6UpSxZ+1sFqTXXKh77oyFPIhrA/UuyTEfQvPJmKjA/0zS9PXY/EYctALEif4NK
oM4heMPtWQ9XQiNlxAxk5WAzCKGf0i/QkZlqITss4WteIiA7jEScjeM0c5fFIutk02mukl4NNR9s
tImcltjRqIz7ohqfwKi8+vvkFvjBLOyjlKtit2ARm8TLwu86Q0CZgpImxNCeDeLygLwX3yWCFCDY
m8RKfwinMK0fxWPjE56/cO3Zw1i9YTeGHTB8Q9KqP12eD1K+9E16Ye+eQHGS+KJS7pEFLynEK7Pp
frVpUHDKLlWnzl+cWG2cGdmxFd/dCc02vtqdKHNLclxw0FLgJHkwFebd6ebtYJzFhfrg+r/3RNXa
DQAjgS0MxdoDNK2U6oouR3I3fTnpEa86A/0TqhUPlS/taDDCBxy8lGrefaPc3CJRjBRuml/mX1k8
6/tNRmLODrsHki2UsB1uEFo8/YPuo+z5C0i9rt+hMqPzMiopcFo7chWf1Bg7ac9RuI926T5VnJsy
1KkubRN4HsopGhZElMvDnWpEBOXs4b4+kRrtvjftgkugiYVp1aFHnbJ2ZdlCvoKD1fP5XlK3SnOf
oahaSi1wpVcvns2M5zwgWDySVMWGihUOcQ0pmcTS7UDv9UtKPiXFU38Iib9aTJ7goSkOP/jKGa3g
7l6jGDi9jvi0Cm5R2G1gTVhCUIa8dKFZjcHuENjJyX+2L8PLgJxbjv8wY2dF3bsk3JAEAdLpbkZM
mFfuhvQHpQAA4F7FDNqhZp5pmAf8NX2q3ZtAz4FjC1KnlluJJaQsn315YzhXIyUeGFDUdO1NFsW9
YB+t2kbrqBAeOF/9gIa0ctS5C2+Cj3uHCt9I1IXycZqg+qStFgwSKiWX0N9KNSWTXlP++ad9ph+O
voQZZN5zsq5+p8UyGHuAHhETytQxOmZH72Bfp71VJAwgwBfsotS/auIB+ypI4y2uS15ul9ulV+5N
3BBATiUayzCmpuUiaw2LnCNQXmkkcivrH+lfDB4oRkK5oy6uXCC24VggOpH42fNXa/iHFiyxLDNZ
H8ib9ZhkfevaLn5a/fXCf+aPchYgOz5QKYD2SoWbf7Psn6CWvgJIuIj+ZinFlBDO3VTvoFjUeIoG
5DXzpNjj6eKA9G8blkZKcHyvMP2vGuo53AtAzAc6Df8AYkoptOoEyX2UZPIHHF2Bz3z0Ju1fT/yq
z5xQo9HY6S2lVllbF8F40sY/VSGJTiKAO8rPW4SwcCfv0frYOXfmP8nuOvbuMzeV31sh6upfYyBm
8dfzgANmp2FBckI49VbbGst6MrvoBKMnyD+ebwi2znbCX1AmSxPttQfJbOWiDoHBFYmjvnlm6Yu2
CunH0FO8XKbX5g+ExR08oHCATKhCECLl8ULD2Q7b5sb5kpNiPel5nm163hQ8K6BQbal10nK0k9b2
nNRrtp/w8HMgOYpOKeOB41FqnR6+xDxDjcjc+8YOzNrOT9VYjC//i6457ceBC/9mMMZoy5dwC2db
4Sq3RE7Pizi97dPXke4NyNua+hWEhpwwJ137/f8BS6WmKldYUgRMSxBqNa8Qi9Wa+MAI9lnlXVxy
M5eEWM3aNHX2FefATYX3xEFYEYnMpi7ftKeiIr5u2jsa6j3I3zyno693DNnAqF74YigEa9J30aZX
MGe8WAtMVpm4I7KHXBZzGMwITHJNU/MaKdbRehLfO2wsXpWhYWSfW/7e9fgt7vHEEJLZupTl3dvN
Mb1pwFDS7Y8vK+gPT76P17ZT5Gx41pF3ozkAwPq591alqGWlTjPjo7tA0JCFoZI/1IzQWFnuyyu1
l0meOWfodNGkkM67sTvSMe00XK69Y5T3sTj858cWVaYwYY9x+ntRqDZIIdd8rgkO7/TSGB9xD47k
nyfM1H1/M22iB8ucWBJTQpYONtv/dQwmx+QburWe4u6I6G+OFsddxHkBGLeGPdo55q9B1pdEYAPP
xxwxOXdJprtKOe/Mkv05Yh7zmPu+bKDe6WRmWPSSxyNG1XYuZmpHbANRtmeH3PHDm6zY6rcfrFh0
FcnNQGvGqN5qTXPWZg/J1uVinaUY+gzROxjmNMNiXCkHLEBsnZ/+4n5oFZg0aHXaAsOveeCQjKGl
APLPZI3Seh2a162F80cdM9VKiwZij7SS5hoOOLiaTj0/JEpM+XpqUlkqtfhblqC/aYMbhu9hSKV0
Rxr86PVvKdaotrEgUptnLD3RC7ux7WYrMCn+OEO6TfD9VW1ZZx5h/bjp9wEEFX2KB+AiOkwEw/cU
6Si1Kt/jSVfodMEsSaXStxaNp5lGOGREG8GRXM3rbGuKWh0oVBgHf+NOl+HHMPjXJAsj2HG7LNtz
BzrGfQJWm4tuV6jWuRGujlJs+IImXctTQQTTEu6CH0depNewWQ4f5eIj6K6tWH+pbcwq58xL+N13
oMSMp1SIt6WsgPG6Mxq9+hbBUN9/FzXyP7IEJz13qMJ+Ytl7UERFytj+waf1mWOE0KrkTZddcMAt
HtD7s1hSJ/o6Hntfc/o9u6fRp2Ohkc03r5wN2JvEYtlDttl8vKIqFJLVu417T4abCeP/z4ofnxPt
tw9UpOCt18uYc1qKEW9XmUphNVs4mLCWBvG98sNJFLMjwg1PBiRQIgFOg/Hk3MZiXAugUl/Uy/pv
Ya89w0OXChKav+jsGHuw1vlK9AC2gLj9DzZ7upYvv7IVrUuKZxEXOpt7H36J0Fyl12IV4H5O4//W
8lFKYxW8mrwdlf6ECuBvLsM9TsyfSFbp5ogBTrceXIwqHwJe3CzQNQzRAu7pRx7tIByNxHmkx682
QhtiiXEVyV0fIJIUoh+bMKbLrv8BMRSE8SGnqSsezJ8kwBjmqslo07JpVhR55XOXMJfx6I6ZwxeM
GxcVFRBl7YWaxO2F4v4fdXu9eB5C6Lxjlmj9xvaDlQtFVPJKXIdeF3luG2ytMTqtXL9Z9SB+knXU
weCexPHyR3e7c1tX+bbMGd3CIEZ4OUbNa9TSwgf1via1xmSUCGrpvHLaOnmTkxHZ5W/gbaqQEOKM
ZWsotmDmIFznT9lmIZzRu1VAcJ1RpZXtMzXbMopffXPL3eaE4fnTo28pGsh6j6s28b0Gj9jeWZ7u
dN08lqiJ//g14+0/0riRcfh+V4Orzi8+gpK/rnHBUOpb4iBES7Y4gTJh2PMK7bkwD0M58lEY4HuF
4UimIX0TCM85vLb4v4/l2WDQ93kT+NmsGWuyGjYV1TnLeB+zJi0U75rksW7bseR2aWpCr3OLi7jm
0QyrMEkPXeCqw+QUrjb7D9LdY101hE76e5Z9xtwAVZq2szYtOgcW6bWrpBJwKjMydJYiyzH+gvpr
VX6qCRVZchYy/f+w6EBdTZiQhKrgtgP6Oz+IrYKfSjwC5qduBFofU0jS1oS8OjC9Rnk70HGRP+wm
iLmNqxJvB5sUxBKFEOReupNWrhGwfoeyHh9y5vbH2d6lMiVilf0vnMhQhioqemMR/U+DyM8k9f04
sitl+K48IjZBEkvviJVo/Prt1t6MOZ2Ki3ofSm8O7U79G/g6fwqC6iPRcQMnCjawabi78X5Ycxpu
9xum16O/qHLoMiJCcdT5cODTnZz7M3DMOARQdvb+Si6tmqN3mhmcqeXVQ1FGJLDkCslUv/CIqrHf
l0XP1ioJpZZJhXmPK1XkbpmcTyeThV7zoua8P/NgJA3x+27LY0+gF4Z5NT2MfH0uu0e15hCzRsyh
c4lJQ13+93CVZkvlERFpkS4Ch5Q7Rhwu4ExTrgXJ59Q7p4Otku8u/F0nkJAEJ88I7/A0ioCtvICR
/XOnV9V/NyqqW/n0cVHWyBK8l2WUxMLL4xzCg6Bd4D72ef5MITHm7Tlxz0FeSmGSWuMRS2XCq/8H
pAIchkH20ainVgmhJkCIbX7dfUbozsAJlto14yz1uGRicmmqbM/c83gM5h54D+Jv+nbiQCcuHhL7
/jxZj1Sxw+yZzhfU7NTauYq740IUdthca0P9MK96kKbMHx9ZQxoumlFLlkxsDllg10GuNYMtFXzI
L5fWaFhxW6qySkxrLm6gyPIaXj3mMbZRpNvruGOpxU1m/h64egv/TOhoqcDZhKVuJH02T60r2mq6
z8OPLHeJsEnfzoHtEBSBGq5fzFJfrrxeEcf11etm97qVkfni6OlkrzsMM1EJb79yTIickM9WHI7I
ZCLaluUFJ3ZqnhOfAzX+0qd7zLc5nbfcQhnNvZi+NbEaFSsYxSe0rlFRudPBO2rwAHVFwGbTAGbs
z7AS4EIW7LuaEU58vNH/Ug9caPQJvXmpLd0tKdiBme0695/AyS5uayTlMBdXwY7qCZ+cl3NnWBKN
oZ7GpB8+dAFPke3N0ZQrwaq7CPwretjbxXLNpvZyLkof51kTrWjjfOypGVzbjb/Fjzs47l6egOTX
9JzktyafNtX28dtZQtFa6CJQVFCNMIy8dEHuwTAdTD9R41RgZu+kHU2wt09djQqAgNJ/MsxQBRwb
BH8AnHjbxY5S2KsLmijP90PLgnVnR4zozkIz6GG44NulF9foo0HPKOL5/zGBBUCcX7cBax0SGzmb
T3zYph/k2oJZ4xdvumtCx4fYMV35wAxo9Sx5Aza70QcJuUwdoERBxxsmW6G3qbM5hjdzzYmytK32
EKd7cskIAzzkiMFvg4j6UG9elJ1UYSrDj1PjDeHtQPu7qH64ZLGx2OBy6Y4//SoghbkytgtzXUsl
AcwN8xoZ68rwXNZm68MbmhS6TFnxyCWoYPBIF0/qAZ+J2GftOcIUF3nrf/0XFWVvdXHsu0t8oQ2V
8qb4foyZKrQsPIE4WYVKiqyh6FS6esvJyv0gX9qMvlDGiBGeksLwGMZfq50drcxc2BY8P49KVtpY
cUyd4pN/HxxNjphMNzrH5VS2E+vMBmlQP6q9JiD50bxARE2a28llS6YDdeTuH+57fqVOgmJCDzEf
untmHzmmW435+AFAkGztRK0WcB5SuzfZ4VriA63AtNcpXP+rHaNVjzfspBJeVjRCzYtCSsN0Obsb
+4GHEbFAc+xTli38sn3A/HEm3vFlpGBwM52jK4FPPo0t8uw5ZWQ+/GcOm2uaZESs2rs4Vrf8/+Nd
3p1SifJE/sxCc6HRaMghLJbcJyDqIxhyxTpNrqX09yj4Ej1fMiKw3IYpWx5eAIcsVJ6tBVyyRKRM
R5IwqOTQ1tyQ0uQ/fkOTRZnJyRMqvQiwda63MZM6M1tvswfC1LCsxA87hdRnH6KOxTj2WgKpbInK
4otrNSn2VNgqrGlh3m88gm1uUKCikKbZ7kbsegC8awx3IRZptp5PKrhuT00LaxR5Cdj6u0ZBRi1p
voFRHqH1HR7RLtyRFQSdOgiV3NWO4mvwXVyE7fIuqS28/ZIAhvvIRESsYzsojYJgX+yeox0KT0SF
BVFtUxwioAMJyxtnj9H5fidM9Ei1t9T4fAk4uDtCpiVRQLPl9i6rm6yNoKbESghQb+BbB4c14BKB
SxbELhm2e7jGTtU14sI8hyTvZ5S1tJ8r+nbDEt8Plb5ZVK/1XOth/pbjmimHnxRUZpR/n1ne4hmj
CCUQmsKnACiag+PKj0C1DELrmVr1r2UfsXtWby2SXxStRna6wRHs0l/iUIzicRHeOLJNOiB6+0U4
KDVaytBuqnsuRWgc/hCAAPFghmNooFYr5czcmYCx2rAMeMk/xmSN4gUBaKTeaM2mMhvBl70GBtT5
aLWWN8Lq8NHENGp99kzA0XbfT3Wr0YFym6hzJDeT58WKvG6sVSRkS+SUn01q4JT0x0oocKAMFGCR
CfJtVwqNk8+1FAzEmHUWuPWI6wfUXd7k1Er7+6X97In6xdgJum2O70c/YAskSmxLCU6x0hJ9lKzK
Av/LpQkVvrXnvbMwBAz63cKZHI0KH/5ikO6Md2cdWDzNLZjGFu737VL895kGTRe7US3kfy4SEYS8
Fc/8nfKEmA7tNWo3kIACYPdUVognRwkxeSi45ISGF2R3tStnTUSz6PHCRL1qrGCHbSCGRqseh+Ey
uspGhWm/P/AhWr5Rip5FBHcOJUBlpL6uq9SE4Oglgk3IbLGJ9JzqE5Le1ECt98QaHPKVUnTS3LsT
dlrpeHvM95VtjhMC2g+/w4Gk7oG1R4zsbuoY8EssSE6XKztvgO8IXXQxq+zRpEkQABMxLV0S8xbV
vCoiSFb6gbo9lncawbpMKIYCBMrIUdsPA75SarDzNDx+N6Q8NdjHHUIF9MGZi96F+L82yFUxVTa6
YE8VkuA14IKTAJeG0TcnpIFdHezOaX3HZJWM8/5jkuruw+FKdUmqRvv64ML62JdbEgmiRyHR/hzE
gh6ISNMiK61iuuab+1RKH3flCU04pwcsKujfKzLLsUKiQEURICxIvSMKZRKV4HHVCbjPAfkwETAP
MUT8nc36M4eFsO0MeBbTczTuNvOg3wTuRUkMtxEQhQSoUx5HPm16azZc/L/FdeapNSlggfGNKt6/
LznV61bAvnsz1GQ9OrE4ROooqIA120eaF/3H6PbUR3473BtwUWx10D3+CfSW7+CzVvx8AdXf5LAl
wnkJhL8SfpiU6T4riQwh1HqD6d8YBMsYHi8kxZFgWhjyixA8xXlRYAYyBBlX+/zZf7J3vUEcYK3R
mCx4Voeg1qxU02nw9zNOWGeIl+0piclO+eC7Yk5CpwR0BqqgCLa4uQ9Sabx/SFSzOZC8hZOofBpp
VAFDLp2O6LIw9Tg7e9uwEoliEK8fSInj4BOUmq7Xlh3/LA93fbu6pSFgD6EQ7Z2hfhFhdl8xxWdN
8vJ2/IVejfEauY0xIqo2DnKRTN83nFTVn8Ejz2kOZ2/SHcbe+FAzNjcL4K7KUMaoRUWmC/V0XwU3
+7mYvNDDh+Rwu79lTZyiHnNx+o468p1c/ygNgWxCGvScaM3aX6cgJygnNHicyzI+Il4ChXYOgeXg
mEKLbPGkqpGsC4ZCD6dLKy5OOKqULsEBOsqtrRTUfzJKhgRAROvDIw93cIaftkxEtDjBRv0N2D4R
GOETw9qVPspwGYfHpGT0D8jJVdjhXcESl2qUn7lKo7NhMgze1FJc+22NJ8Fo9/xjhAlwNU/DXafw
sSPTZYkm0jwOjMQ4jgmLIV1QdQtKX6/wQaPdWnCWN5X820w+ackorhxmOByfbaasIS094uiCJZ9D
Mc4Hhh+taVmHGk8535G/DtNRZKaLo7feCE4W0omdYgsWY1MfCmzFuUHe2lDufva203t+wYlea8tD
DQZIv1sV/uKReqXnRhXaMoLvucSMCVwVem0sxh35PSODdAFEljTAr+/aA3RQyyvMm+3KNKNRXzwz
3CnP4xtSkDOnovM5FdGXNJ0m18Q1pYA1Flqh3wH+sgledifWJcUoy3w64kJ8SkwvMOfmLsmFnNy0
w/m0sG5A7c9splqE6MlFl2+JxN8g5YjG+piQrsslVNVBLsJ9eOJD5r+H55GUNJDpksWUx1pGU8+4
iOTIWvkX2la3O2igNW/sgI4iIDiMRrdc1Aj33heXPXSH5KPn8WGohQKz0voH49EwoJOMmdp7YjwO
eL0V9yWZ0/34aXv5EKjmx5YC3Pczra7h8sHUEYYtheNs7srA85WZlVWTcIWn7P/fy/i39oMHaVtK
OpxyQdKuXCmAeSN/BAKcuT5Y1/B7BPaLlR9NmDN1aq5NX1IfTUPB5xyytUXA78+hNKC4v5aSVkoR
Kj+J6HJRLRNaLiQ6Sy0FhnW/BYl+0goL9ds8sIU2Hy68Ya2T04CwUSHOoYMfYzneF1eJiYDGH3gQ
/NDhiFi4AeSSFDwOYiagPcgo/81mwcGeLQwWtAKqgeRncC3VnKHGlMnQ9Hlr9jSws7hAEiWJs9nm
1mUsSd5cBG8UefnhGNcploWYz7kb1D2uJCXrN4x+hnkkIdB2pYOlBFYbWvvzgIX7e46GcKiY60mv
6l6QT8Uh4Jqmz7FXauj9Xac6HZ055uLmiwz7+x0Y/kf6yRWXTDNnZWkrtTRaB7UFrxCZxy463Uyi
AWXpuO31+iBY4GjbcAlKwsLfDdhxCkEOi65rec2PMEGfmsKkbGeUXTTtDqQPkBpUXBJqsLEMcR/f
isN2O1UpBnAS9KIapExfFzCE5XLcF9P/MWiJNe/x04ad0rFFIw4dhXpTSNZ8s+kYisyUmYO9S0wg
okhOTC/8GKSyQrcFBuWGHhDbSgowmPlgp+WY2zVafuZ7uN4tkURTU1A8IGc+IQ5EFsijgd9s1VFo
qTULfVKGZYvJdqa4ioEearT1ohQV/mM/ZZw67Gp6mSuThlHq+suLGKvCYE5Hu5z5jCuSfGkU+9X8
0H5/9nO/o+zmr1aro158mOZ8ZNtxBSqlAceK524NEgufRtyzrb0w93NN4FX0Och3oYWdcnqRD+Se
LlTzvhAQDZRNN/CxGejxkai/sAXbCQpjr5oGGXOelDL6thdK24khZ3JRcpnsWj89Pg6tRn+1V0Lg
EeHuazTY0JSC2K51tNOUsTL22kjPKgesQvwRtvy1h/fO1upeaiC4hswYaLnBU872lbPlqhxSAytQ
Pr2XrbcUCRSl4rlCAwh4Dz3Y3ttpaTlWToxs8H0qlYZKShAbLG7qLFtSExZ86vUBBft+np/foV0o
G1xiMU49BxCQKtH/g9hmnK4VSI5Yo5z7ULgxZL5dcVLZgTpeTJ6QT9sFqoqtrw5YmQ7TfKzuDa/1
x7lI060XxV0Oh4yuxxQ0xPilLjuaCivkjnzppAXDGtTXXbpPjj2VdreErM6JYIfX+mu9xQpE7zKn
Op/sYm55dFsJoM6nCaSDATd2YXsWss4ycmi43c3tA2fqyBu6l9qZgEpSdvzi4lhEKRGw5uM44/Rw
4FnziCXna0HWy7JHNx/mtSJ7QsaekduJvVq4eAsgng1C4RRWYDVNDoRKpHR3TTR77ypsCoJgBXCx
dgKzoePPOisaoAgKEE7U2/wTzM1RralMh1k2wJ8BWrgBP5/nzX3G2EoOGDjpK+mFTMmrqlE7ofR4
zlNBnaLwtw3BazTfj+2QAhiGZsYqmMGKXbn2mNpB2a20QVwzt44+9MfjgOoAUYDFzfrvd3T3IhIz
rDTEFq+JB0MUTlpe7SWPlY5oI6Jkvygoq8Z8DRWW/b8+lQ2puzmKf5DQk5RBi2WibbhEw6GufXE5
Cshg1djsTF9PI8Q+sPdvSmHNEKh+cdY/b65bs5qLq1tqvy4XoE2yYF805F1zHPWi+7+7b7SoVw/5
Ux/pPgokWLnhlYZs5mwmVeMmSB+QBDEkKANQlHXQKbevFTOfJCBTj4ABY3ch6+84XkabWvLbwRxq
TOvCOoBBHB/+o8pkmHnXFEFIVlqac4giPnl32Gf4zRlfzTazBFxk5BAEFdAHijO6vpN4hnNiZd+0
ovEkZGPR8ZcGXFht/e+5w/OZT++v6COJitZVv7jstqxUUPOWWSrqp+mVy7BXu652YU6fCNHNGdUR
hPwlfDewMgXG1Kzdvdfl8tXHVJJ8iKsGrjOm6sRx/cfXMyQd/JZ8JhCBNN/8F1rxCfgGsF3slwmk
+c5gJ6IlG4A2buJw2f8BABTDfLs8GJAYKKZFN9niJ7tbJqGOiW+QVOua3qiWEIQzQpbaAb6M4D93
WOykfUhSzxjfcEazo7jf6yMoXHGEPDdcYf5rmjryHHaNvaNL54nifYeMbVCtSwn/bQADxQhGc7SN
AK8fjohgK0xnEY8Mujs+Z46l4L1qp2NQAsjqEs1PZQEl485LgnDiaffDZnfAz7j5a3dF+io4W1sY
jrtJC2nSlFIg8WDYpVrOJnfesNCWkZfl7O1Gf26dI44dUy57Jf+8V24FpJYD6Rq1oGDYRynU1Cv7
M6QN4C3OyETvV1HYVDYcoC9TaJoDq1NsoKu7iBTsTyCWh1b8IyhfnuqqNQdlkJSPYXpva+Dd4zoz
GlaW90TjxHPnMuNEeRO2pFUlZe1Hd8U878Mc8gjCgptt/Kg2YstrB2wgnQowivsuEA545wU5kuls
HNHpaWtRsL7zIh7G2ClnZAF/vuhVcQLeWps94F3KiFk+aUMIf8srzmnVnt+N+23zdygw4ocJB13B
xfnTEfutxnj9JbJQp5zOmxYRXpD7FzWqEdkRce3guZ98xTIxPGp3439ux3ugZR5YpreDpcqknNwG
IIht8A/oaUbc88XXGn6GhJGr4GQncAYIoyiHN4q+DPhRCf+6q57XbztdzAa1I6l9QcrtPfq812Wx
e5zX/moIFhpg00UF2AvtbWfTCxnPNDOyE9x7ASLyj1N0HVknq2e6vfJLPtWMPs3bd6Mn81sEUaHJ
NwQfuZEMSICEJEME5OVcYHzRAaKs7v8pw/EsojMsdRbicVBRtYkrtB47CnziSiuU0GeDIthHRKCv
PpVjRUxxj3TGdWceQ22eNKwZofTPahfMRkV4npW0AMfGJjeVLpZ0Czh2n5RYy4+gW0PJPIABM2k/
3c/f+jYtGXhqManyRiynEZaaHBz5MAZLXt3IoumvLeY5aBK5RKTz281VVpysp8JkbJ8BRa9GTZ6O
toz/bazPAN5QkVpK9SXeo6e7tWklEeDfLo0V2T70eEEFlhsbxZgvCArNgMnnHn8E1g7Is3Trzimn
3AAema+x+R6Cn58Mmu1nH/Jv+6KKhahgtd7MSM97kq86ESII+N8fTIqOqE1E77H4GftDPtXdSR30
2kxazlsuQpwMRVEmwOE6KAa3+4tA5RohLkn+C/3HziaKOgqUt5UOnrtDSRoV/Tdp+7xTivK8Komj
i9/ENYvECRNJoJ46Xm7eqbrOX8R0/lZ0La88QvMu2cYC1yDrxNxzQEahcn/CHA8qUz1az1xSAxA2
/YtvJRuuZ4F/8ss7APweBnULZ+Xi8qiiSgClg6WbRjG6gbs4Ti3L8dhaDdg/d+bWfs6cMWyl3lWA
+TeSuLG45Zt7FCrRzNnmkqrlcyZJLCKdcq0RUa0F7fjwAU1jC5R/gn8K0ldHAQ3Ac3mux3upBjhz
tHy/ZIWAHTiKb2ILyH0BJ5gPRgVlyrb0bCB5xO811bJ1Ie9edtmy3D3lQqTsrCad8/zHayCAZ37H
3sH+pSNbWGw2qeRSzLe2diMwMPLN2dJU+piUzF5Nz/DwspzgV8J8bdYrMBv5JJ4NJS0LjaNDpRJ+
NZ/hE3lZnvIILNpKVhdHD9k7WsUWvqBU/R4qta4ofWN/9Oc22XGidu7WfvuYIyStUfDPbnG1XNgH
l8M5D+aCYn2x5Y1asZUXL3GXLcJFPpEGZzJNk/tnL4oSlO3xYGFIFrAuJXL5CQHfFcYuszhlPSsL
766Gx03cTBE1OaD6UFA7GdtyVN2qrL9id98zXs+Fi68KHzx/W3PlpUo9oc7WO3H9BcRGGp4LY9h7
n+9ilex3N6Zr1ekBQBGlSTmPgh1LPduAcTBAmPeFcT9GncY5dQs5p9a4p/FOvcbmyTVj6utBEx6C
BAwDqFfN87X8uAHvXN3TplsNIpFy5md0yq7z08QdqSMrJVAmTHSqC0ZCErnb3j1jWYRrkutrWNKb
PVnK7afCEr8hGf09n8qYQNcvdyMA++HClInCGsk3qGiUyjouH/31Kj1ph46RfxL3T5FbEdUVgbfa
ysVZkxONMmSzwXEMzqjd8dL1lcoYWgQiFjP31hup1zmte7wSJ/jXT9bE9Ot+grJhSWH2uPdIQ9cj
tPmWM0e/17JdL0j0HoERuJ8CiyotBZdJsavRM4s+qtGrlaUGIR/e4orBqDCnCnD6OJBKy2XwRyFp
PLZtdcREDTMFfyV0RZPePPG6MX2hzokqphNHsc0cPVEQsU3zOTnsvHq7kbfNikrakBOrHITHDqib
NsySY0HqVyDDxrY+gFZnFYNWhtNlTsDU2v9QqmVismbXx4zlgq6Sx6H6omnXz1+IJCE5l/rN6FCN
ocYttwmbTIDO0eWTA5pYBqb8j2SYHJ46WHXqGHfDN7R+s6u9sOt2rzyN1duymaRIEISIrhvHFGyZ
ZN3UgLzv0HaIkMW6pKkQrGUDLRFfKubgzIqiAiNmjh2ufOFdNqvJ9djmXxjpaMS4eYLc9uckB+ml
o4ApD86bgkBEcZ3w+PdGjcj+OJ6WBpZeoFbdOR3PkHCsyhnFS0OThpjdP0vUUixNV6J1BIEseMj3
cZYmoNgs8x8X7iE/efNiQp4eDsOa4CbrnN9pKySMJTPb608HQ5iJOpNAR7MlLrKdbbbD+w1lg1Ww
SgzszBkPA3arBCh7hPHSDMUKoI/b/rRBTXezhDa/KGo6Slnfnuop4cb2LLS9CSulvsFygF9NFwN0
BqkT/eBXYPrRx4Ev1qCfXlS+cIu0sXp0xd7+lr9/oBGXRxsYWCdIveTQDOg4t2O631PB9GO6b5dr
9+c5sQ8X1s9a1VWuIsNY9RAQJe6wEgGIXFhwbs1nEMqwd25Tk/qsR8woXFU7rdWgAFg6PTTZY0YS
Ch/8vQ3rK38YQ4mQrrdkFwMyKM1+Uevff6y0xjyfk/y1foivwUyNunoYXLYxgjY3xfEcwtkuK19Q
katzjhXD5csThfcO7qGJ12fJHuPv+JUAyymP5ov7gt5e3k5pwt9AYW7QMwxGbpiRq7wD2tQmRG/A
5ZEY4dyHY5ha8Qsd2oJv9iPbk1W1dK3eIBUBc4GJANvkfVUYOXRE4BGcXcNRrqoSmKxEY28CCS1W
c6q7J9Lm0bCDm96VoItYydoAiDVYi8blwFH4oj1cqoHozOiJBNuLmfUaVScyRB0VeiQPy9aIumt3
iflumes1s7J6wymv+gxS44gT9cIcICKBD3/aQpp+WcwwZBeRq+/qd6fdwfBAY2yn4uwg3cOb7Goa
sXAUn52bJBbGEoF3a/TOh0F7EnkYmjYPXOe2GSeAGRqQfwzIovyVxMKE/VQ0iSxn/aSvvxo2EKyx
8kJqT4anuK3YlHJyRud6KY0/tD27/3VFc07yQL45858D6E1468xMWMlwxahbd+DX8E9r05ne+tsS
VZRGs8urkWI55yha5ePR40XQ7Pe7ABA6Kl8EwS/DVYa3Z4X9gS5hf6TPblQ3XZn/MB2CFd8pmToZ
Gm+AU2aosufRjxu3c3HCP3IvY1LIK13VWGCfB8/CiKs0sYpuwuVO2oj/2HWPBpCUsbmLQCnY7eZL
twDBlIX6KTnMQFFIBwM/4oOpgzi4cvR3E70qzs7CpeaPnJ0Db+/U1lvEUzp5liFSHJwiCRlmZpeM
bysrAT3XE/mNpDV4qsgk3Y3JpR3iWyYX38vkW2hufXfIxDmzz6hsiaGrL+HQioVB5KxBzGQt1YwY
gIaNEdK5gFTOHbMkmzvReiYlHsebvNyYn9NOHHWLGjogZoSV1d6VlAtiwoYw9eoKA4yE7CnC9/Fe
2HLVUIBHm2xXMT2auujXaWQvljH8Ov/LMn/EbbUJhSyF8shIGTwLEHzU35JCpuv0spNAzNGO6Kgb
blt6LZttUB0ozZd8UGZoWgOxHw6CNalR2dqSlw6Z6DybAr/IXM1GiqgQ11wjpFxkOqpDvH80SzIY
j6ft590asY0Rgk8b2jWlARq8hDzUokfSpE6fkUa1ov6eRM6LY3nCGZKRJNZWt3k4Jb+d88Z+CxED
S4Z4p3jAh8327EHoH5R6fD/q4ow/WZO0sbw1e0TIrj6dAWl1HEIWlv5OMslRi4vN56Kr49Uzcj11
sr7bvIi/0KnwNZsGSolLbybt5qgXQcGEp1cHytruZ6vB5nIWekVSQOj8MdcMjbn86PO1qCrlJzvJ
/oz6aooYrN46K5lKUo2I49tnnAkcw5ZUkJuqt4oTfrLJrW9gwM25OMbGchffw44ZOKgYQHfyG4Ev
yVirTAI15aAPOuKUEn0AXBRp1DEWWpGnLd0hZ2QLQJlXXR5SPd2hfERtIfPbQBg9Twkp0jk9IM3Y
dwQCY6Kt+XXDIDO9XwU42HOn2JUyHc2Vt8d9wUywP98+npBxBdWzXzx5U/RH7eUg/GW6hqjqcljQ
mD9cDZhLuvVUpmJ11s589Vbj3K9ZGXCzxsnKjxxYNLoXxApEiD5iOszQGMZgGzqm8R6Gqb44rFQ4
e27oOWCd3TpBzlxFpyFEnL2yJ7sMoqIB++fYpHSsfwuTpuB5sJTuZR4VP/r/t3QMSmzxLTDmztUg
Xz4HqqNPYqSOiF+5HRukP/2/Ikf3607aXiXFMaO2dHuzCt4PvGKhm5y3j5F6pNbgo94QQFym6XUA
uYC0QC8NdtoFwAVjq5ODPxPJoxafZS9OXemipk+HPoArW7x9INy1qXW0LkXrcXUiL70IVsms4wqv
0tzWB88IwtSEGgcwqvd/UPimaSjWWyUV7l3tCiX9dPqCpZnlzSg+fHnDUPqYOLqRCwvkVr5TxOZk
E+nieBUcdmxQ9v7BlsdCttSKaG0fO4U70qRxV+ZXY5pn3ds7OhvbojSXEvpqC26sU6YcmgClqnI3
0MSQgbddf2T9BC1z7wh10ANkbkc2I0xfDY+5qOGW//1Qif9i9tlQeKgOQJQbY/D8hd8xJu59kTLG
gKT0tribOKRNgex3sKwoLPQLL3T/A+mExRzKmcCObFqC+8XVx/7PltW1HElZZuB3nxjx0ZMtYL/s
KcU2EJwazERkLk3G3q0BpDZQeL/q/uA6XfPrRFxlqIXyf1kLwwIf2q0kqSJJPowBsNYajSGEJtAf
jDIKyhopi5Z9BM3vp/9HAAPNpZ4gQMFlHWy1UDjbIszvbzPtmAXZUpLry/BCutuH5oQXsNw8qnNT
w9fQnakhUqUAIlcEJCYt7uO1eY7WIQoJB3dSQwGkgScCuPOk8QpIkriFed0aKzXkWUACCgkSlpEs
cITlX1mfsZYi2MnX929eTkaX7jAF8b9y43xVOHWzGQw3w6kWuUz45s73bwb13S1xIHVXKp+k4U5b
Pmr+MMsVafZIu1N5jQD2abIdduYZ4ZoQbkrbRoHClyN3SHG6LsrIQeJ5g4FoF4jDdLAYeKXlQEEh
3XK5IpCcVPp0oV9vEfTnIV6by1QGiHl9Z/WGHyAcE1nNi3vQjTjfAMwlN5cjRJqslnTwBgw99D6X
Fh1tX4v5RmHpyD944snQSVM2R66CNNYY15ws6g7J3F8nl/mlX49GKorjQ58VrO7+nEq3RoHjJtCA
Y4le5XVwuLeXppV+Z4bj43MxEXFbYISzdvlqWk7d6KxcjYQCmwdnwr2Xd9KVKLKI2YdSd1ptDluo
Tj1FbOluKILa67ab9a7WLDvwshiO1F9jnOCup3kb0uXMGPChtQ85r7TRxwaqZ8EhetqpkNAQ89XI
JE1hCyXxR4xTLL0GsB2I17wTjMiTI0ugPpL9g9Big2eAqMD+5u6sn5MTk80gZEILLqigW7wfgx6t
V+YRhySk9/kIFmmrefx6e92KYBoEjvtDkTff6f7HqaQhTLXYHytyfZJPO1vCSn81R/u0FZ7/nt5q
FoXudOOqMEh9FjFzSl/bfucmrqQa/3riGh+YfaKtWMk5bgpyHeQw5Z0nKGTrAsEDvupUpAITX5YZ
4SUfiSsQIu6WiWbaeuqx96SM2q3Ad9XEA1zhSWXv+Jzev6FnIhzzdnACk3hNHaH+6C1xTK3p2FH5
jID4Ogj7xwLj2GYq05JwwZaGzpLVNtL7aY0QQLaCGnbEYeTgQwPkSf4DVNkt6yC/YW4sDz1J88hK
pgZTciooimZbtLDV4Ry/TDfcKir5u84r+qVCVROyZbNMthCU+4sF6gxm5dglcM4fsqYYax6jxpkY
q0awhO+xIr9W5gJhiwwLRfJgZwgSkMyvpA6iBvPu+8O2rtFnQk2cA4Z5T0hwuGfODYjr2VQTpPac
S7ZMMjCbNdsHX8Gi1p7edXq5orvlHu3BvCEixHJk5dmAXbtig5gGBBuRO7K19VRF9zxur1Ndx2Dp
6s6OlR+YL0Zho87bv4GvpXOd58v6weACfDnrWknzwnqjnL8pdh+jkbP0aDvOlvBBPHAPxARHzaMF
IjrwS/UQdEbTnqGvAGTxp1YbjNlxz3ueoF66nkpTh+lqDwGO0NT0ZtNN9ARQsKGS0rrZJyp4jm/r
1pIB9TuhU1mKnrrkjKbbzj3KXQV+7QNF0YfuRrAzcNY4iKiKGakQ4aAsM4ebT5EzLgFDaHaUObKA
hc5IHM5lkx2fXychWs+KqcTBHppsMrlHsS6uPulF64jZMUzBJQYLl8cSOEOxtPCnYryjx+QOLr6x
jZUUP7TLgC6iCsPkgsyYBvi58vpfsJdZS4F2IgNnT9hLVMTmdqGebnntHgzNdMDzjtheuNbhIzkx
4569H4pI0D4lr2KXVhOz8Eq2OzTmbSJRP7GYeogslBFDs1yvJgFG/ae42uHvUwuaEkVeEuMgBtE/
hz9Dso9VI/+gUE40mCIdml6JeJzhR0R1ZuLtqUUkvJqYy2AupNY0zJLQQGtDbNBYXBQoJnt0PiAE
xioFuRRTuAQu5+fZ14RE6dfwcxWQIG2rrAm3+I5zzuLCNFV++2tQpV3ywja60yABYBgvnA2/axAy
438Lpdy5hNyx/wPnso6g28+iaP46ZRbScajoC3M0Kacs4rmo8L7Q4b5LW3jWILP8pUwxFNT715cw
ad+J5UWo8YkyURBO33MgmwvqNBd+/m25c1F4/b1vQbG3Qt6osWMqiuy0IDgKFORfogrcFoqKfnpe
KMvLvaevVGZCVYfSXmus40pFRr8NoQlB0Q+PNY75njOPpERhTxomhkkN4zlmmEKyT9AFs52moVdf
8BcjU+mcUvWlD1Q/CRie/lXhiAeZ1s7Ueiotkm2ntIflopOO1ns0wIb9mped1vYT83Ui9Nfmmi6B
yg0/S7FsauyjskT4Xju22Zk04e+/jUe0/rB/WvGV0a9XlXz3ptf03QxdMCsmzmoY6VvV0xIsAY3n
LbwGGNABb2CFMkjPqX7T1cUEIlpgQNhrxiLtipT1a0+hFxwWTV9hOIcEZRKJwkLSTPgsnI2BrpQc
ReBQCoUgNZt28ENLjcKPokGFXqpmfjmV/FvOfRZ5lTGn6nrJS8+hR03siLF288tXQFogI3JkeJkI
0uIw19JmwLHOfGu5AmfZmZkhmJNEVQqnLeWgkPHYMWS4YK+DsOD3qtCqUR7jGu0PSUkDe8tXQi8o
ghhxBPLG4VOKDbVKcbK58BTzej0JO1dY6FQGszCLDX/0FwKIlYVjUOzo2Xv/fiEihIL2HlcpwZ4b
u76r6AWWqu2yfl+O+OMPCmQT7VCIs4az/OuBAVPOinw1psFnyBl2KeXZls2uAalwmOOZgfQl9pk8
xMdUlXr7I9oqR6zAtiZU6PIoUWuKc70WkIf2Ii3u/zC5FqrNPgCAfxdS/srLNB2LXwME1wpMtxH0
JWbwVmKkwNUozNdAOWiwct7zVEx8lkgdvodYuPPmpDTiolzO1yQ9dArvm/zqgU3cOEYSoWvzpN07
M596jmMnxzgt8dKOMsGCR87ovfi0YGQbbuGVgW8EvQzvjTQ7XyYglG/yuWhTejAJYd1eKBt4lblY
Xe4Uy5CXIl4+xBwqc2C2lFTph7DeOjAWEy8KKWE0lVJy5ScAeR7FiDkFOjz7RYN/x/1qmsaac2sO
+ITX5mof0OflQzPPZPc6I/aBo2VTp1uoMEYDqCP88oY55KWLvrmuleKAHmQuUErJfERoU3gdOex/
ism+tQB+/8uZ7SvE/WR7aqML1cT3isAnjZZgjMLH/WTuEHwnuN92IaZfpAae5zvZABnqxeMSQuET
chVhLoJPtBqmvL8Y3bphl0VY0BmfIsSdbZa2lvgFVF7e+FeSKI98tMMgsUykyTC/uqztZj9gUzkB
jXtoTR2GTLaFnpVzakTYDfwF0JNQJS+W5d0P4mG/Kx3ToTyIoDW9PfqxOGcQCf6QgwRu5qQQhYsF
O/w4enHv2ygEUklGFGrc3ec77QzqNhYjUaN9nm0nfSWtIbpdJEsXgUvORcY9x5Yy8biNySejQe9Y
UER1zhJ/jXyg7RSpv4b4CZgZhPAw/8NYJk5Q8tDowxSaInxyc4BTX6mx+dDpbEAXPoEmCdc8YIH/
G5qTl/Bj5zuHdxfGexMl5P4bFbpyLeZw4wWCbV5+B4LJYReQXxUKXrYReFp4u4tWRtQR0BiFHWj/
f4JqomfnIlh87815IOa9nVItVAQe2Zc2qfaViG812qv+TkE9a4nkAQ2DdvM+d/IJkH/I0O8Vfoqs
tFcPaT2FWwGif3OIVxQmhNlV2xtmWfn0KEbXIgFXUUc2Th+JtIJAuB5KCiCnX5rh58AnDkckslO3
ahErr6aqlMdINL1w6mgR/INJvJJ4pxhMg3Xu+MQrDW8dFGxZclTUCVDnDy31jSDgkhLln2KYgh4b
h4AhwMdAoeyveea/yGy5mXxLm7PsBIytpr17Y8wCVduEHHLlCOaSHmrNjJhp2ftuIYctPyVQh2Xp
xyNxC6QN8du2dfzIbB/MPy1l86hxc7D1S+m1UE/jvfZqxkdDrJaFbzF1noVV6hAZ1tO5gA9Jju1v
/QsuRed407auU0uHQDR7MbW4DMpgFKZw6cMnSXHn4csd1c+dWKz7yjgN2d40/hoHwfy4PXAPUoA+
6tmX/AHTJCw6wHQdlm7t5OMnQudQmLR+/7vsLhUtVP7CfYprz123p3baBYbOnT6+z5UzPH8ppgFt
fJEAzO9iNSRLtaFgLc29Cd+hY/H5veOYyelgkBmQ3f/1hs8jii88zyq8RfUJex7G3Giz8fjfTV+s
tk5pg4BMviBqiM0IKxIyqpomQYAH0dUxO/pNoJWa2QUiVvXWzdFOyO7RDgsRFj09ZxqwlQ2mGKDs
u2qO62oswYZf8RZqc+bgx2vfXOjidiRAwaWh+yy3YRweorMikxd/34LS2Hvk/R0qmapAk1sjXO7Y
bcTWOISVzhFlXIqqnxwQd5s+jw7CnNQRbgzUjwwCaUItYuNUT47fgMXT8HNg5/neDFvtXuwdZaRP
AkBhTRb9jQ3KD2X85uOts1QcxXoFiI7IAgobbQSDPFhVF2MCkWFVs3TL1O7v6b4C5BnsSAoOjH09
8CmfngVmZNgUdAMoHPYNvv8X+mR1dTKeqlhcuCUmyWSqIZKiNeu1tL4kWnpVmdtUnj5FCHzUqrqZ
HT+S2cuqyAhOriM2K3EMn6ooKMUzhGUFkSjqWnWJVWrh6ZTd6sxdcnvHwQLblePYVTttjzLH87cD
FTBO2aulQHuY94zZyX501NWCi5+wea3tXooIUAhnWb5gxHENCl/yp/n1irjhkvkOFsu1TW1ZN+LQ
M6smuoXrGkzx5CN+XypRt62c2RK88ZGLwWYPYvx6jORO/7jPJcZz3N5CVEWIb66pJVZsPtD7tjPj
oYiKv3WN2azOrzsbDx9Ejsn7jZRWimeAmT8K3dJpXD/zDzrFoxOVrXw0AJiMc6bxVSkxy7wTO8KD
8UbaqOjAWinFQlwwS/OHEldnx6BnWeThR04FUOJdRJMpAY/PV81jTsT6z68WgeyzriDeO/Z47HWj
XW/E+yZFs212KEL8dwFPJxgZdIfo6Y4OSiU+OBWw8nD5KHtSdbClKSD2TG6myXGaYsbVBukJczhj
WOGhxCJP/l50Ybcj1zxV4CGKdCEBMjMtWj4M2GKnaJhomzwtWr/oRznilliPt1xBZuWKZ9KgvJEz
Yn/JJYA1IhPoBfsInNt46U4ciDXjCkniQvpJIeTZH8lKnuJbPo2iVnSPW7YVpSE3QtKe5+89pepq
4pRPmGCqJo/50lI7Bb9JRMH+ihdSiN8Y9fKzODbx5uPzv0gy7V3unJ8J/NdduMvVP9IGlfSkuKqn
mbNv6Umb1ZavS6sGh8U9QCkKq4tBda58PryQJl9EZHUiGmlVgLKPCTrTQjAg/n/JX68RwDh79W0u
azNMekTpijNJ5qbnAtB5JtgWJ2cI88hjomfb1uV/wH7i+16o6EPOh5Xno/Z9N4/vkNdP/vjCGWl8
TOTSryAptj6mBaTYknQ79+5p4JQpZB5+MzkZEPIg0WjQl98Usfh/h1JcDYFCFW9HF1jVPYLnejzI
jn0D79cjAT+vEBpzarokUM0EK5j53H3jm7gSI/cVy0urxY3C0eQDwmQfXfso0z6iYv1d2lRcRWBe
lUE+fQV1U+dLj0csY6jKM3ybPOz5mqq1YxdHcwiLFWLXZYnTnqi8nOxdUpHN4Y+h69nQ2ARN8P3T
fmIts4wY561zAjnki4YcPQSsibL31zPIyqin87wEihqVQ2YwSK50Y4kRGM6mwPKC+Kw8JVCsHrg6
P2Nkj3NwDGvLRUxwXV2LW/dhvqgHXuMpqqnfSh/g+gPrOkHg1tXwuh7ovOdpVQ6mZXz9GQmQDOGL
r4OBdlezSbwRYta+saGqmLbZw2g3bUN/jMwiv62BK+k5ezyf8g2FYmcwTTGhrK7XwKbXIBo1m1wR
b0meF5ZW171+qasE6pA1nBynY2vpbKQF6da/meCEMLXe2O0j1F/zeS5g/ne3DFKDJ0IYfeoTc1IS
F02B6OLAH8A0PyiqaNCb19GgBGsTIHN3YqdBPzCaq8Ejg+sm+Uwb8srzoAp6S/D9F5c8JVLUcIn7
37ADDmveaJ8T/6DLb9Fc6sqUlWZN0Y8EybkT05fGlAGE3sNDMnV4mAQmK3G9FpaxfPpcnh5TLLBJ
MLOOhlGRqmBOwACWDDXskVRpLYrMj0g6JnC/ucJRpLGHupPuQ6Okb3P9P5mXQ9sEcDt1YbcqboDv
pvtARjPSsYmYkU1Q7zUlSCETFMpoM2iWKb3WRzogOm66KhD2sOXkMqNDEVjKkyHIlTznLFwifvpg
uwtbexjvzIA/5iaUjCkMifgtch810S1bNWNZRkKs1n2ZyPJqXtkywfCxL1+wcziRlvNvujHJXQ8L
KRXB61C3bUSkDw2/oAj/hcK0CH1UjCUhPLmrYKb7QDzre4zo+MX3T7nkhZhC+mzWGb/e012ABXGC
3RZmDvW2AkQ8kfr77zYNTdcDWSzIoPIZf8QeFmnfJlB0zERqQWEfZw+EE7dx9spFn07K9YvjHdNH
k0jCHvvmJH7lejsvbltM9t2PIgkkvcYSCFJV/MFoMYdUCi25bQGqYT4ZQJcIDLofZdnzZfPlxnJs
gNQm6em+4AAWIIafFKtse4rrCp2uo1qUM1hPfL6c00C7J9J2gD2CT3a0YMSCqhjLEtxDlcnO8Nu6
8jcbI1GHtzLJziEL0RoNs8qm9AdfLDQZbCcxXD1KnvbbxdSlBV/qg6OzJwh54p0S45E2O9yTaOoi
MnLUQI8lIITzKRjvgZMHCeVsl5oUrvMXezKABTp8uJYoqYzhpiMlSqeL11pGHl+LOcYClQ/oCqws
pcDVcx2EZXfJ9doSlwmYdYJdZ6WaeHD+FZCijLsoPjKmGcjLWZ/wa4QeQVpyJuxdGFEG869TAky+
y/rpWzdeFhJzzjR+EcKS/Z7jouDxE2EpyijjLySnRcOQPeTtmArdiq2L4eAcEpfsKwFtIq9fnxDq
PIeTCD28z+9ZSqzmyjtJvd/Bgq/BSuRf8vZ0drYtkFajj4qIVOOeSu4EFjEGCdcm4TpIALL3iFQb
plilkdoz86h3vi3wsTQcDVxLv7Ig3Gc4K8IFvz7jL+6vr6KCoaoJWVrHQHFvnG/xhNOGLduje9jc
Uerev8zdC5La2y6mPyILPNlW4sGhRXB/ul0N+bKADjmxUtUZo9pUrLe547duVaa47d5W5VFIEBFX
BhviCmJoUqyg57dnraD/hpwkjGFIMTp+1Y1boqdOp3kPTtpRYn3ZnzMGjLnzrRoVh4yqLe4lwPlb
QoFsOO9iLrAqTcXUZGZvDdwDcjmZ+9kLHXw18wKkKpqT+3OW0V1rB31gWDqYmo3mF5yc5kQv9DOA
kFt27gYc3STvpCHUc6pciIGJev8FbadpkabzdHcDsTlJnuqDinSP6Id6dA+11Z3LzEUrcduaijC5
Ok0xQjdsQSRD2TrtWzfLkLj4XCrqJt8itWpzlNPRLkChgpfRnWAuWoDlv5lflsrdai/8jBnkiaLK
AVP5yPKLDBYX7m70VD01hB/CtCOw0bokFl6ZpzSoNHFuOxf4oN08+jnsOxBFSRlu4FDdU9LI8c1C
fiWkEYplRvnO0DP36OpqaKZB+2p3XGsZOsTlYyxH1PT9oX0fE+7hZ/v86ToAwRV19h1t7UpRE5ng
ZgK7bsPiv+hMvqNHFUJm72rcRBXu/NkfcBAdZqnVKsfowbEveA/1kUriaLSX3vgDEg6rzWXs4prs
jekFiYpkCsvNoR2k/Wz4tZDbhC/YdnZXKIA3vQabEa9TaX/OT+ZXXnqDWpbTonhEmTGVqSibrkhz
gjLVPZtrYvyQc0/7aWSVESMbMDRDPyHg/lJZNAoHv682jPh0Y7T1UUCdOa065O9UpL82sh3YVXQJ
VjCI1fgfUeU2kleuZM1ibLBMNKm/xd6fF4AXoic8X+POj6UBnm8RCTQaqc3X2AZIqgowRZ8mZlwB
ZsQYSciTVucGnAF/oVDxItpNNbVuCvhwLP5U8jE01jrpJKGy1EZlyfWM16ve5KySCPrLLUEg0HKV
VD3e7s7afgwJNjDOOeV+lr9L8EZHhfgcsSfajiUboerJAWkbZmOmSzIErzU0GeXkGk7w0BMiixBn
HGQaFK5U7whdE/k5BjDdN0TCdbhFfcHiBlWTIXAVfDhIFCQUS5kgVR4Sjl+i+iAZFadTo6jhrzbV
8mbK2wm+Bcb7jZIIGrwah3Y+c7LwtRZeQBs+Yjf/llCam9M0U8+9WjoD/cF/66rjMivZiiWqV2Hd
ogBjWfd+uid/yUeddxLob3/gQuGZSgWNXTbWmU9NJHhnTJijRE7g7OIzvMMl0+BYM0IB4vh2Crvk
24jFGZg5wgwWsiNhfgIXwhZqLSwscbxoKYwaaWleYYwPcG9fg3BxrMzghOICi/A/G/AqBrCOVZtP
aZgC4E3ZJDcD7XINCQIH8p7/TgpGkG6WrdJgJ0Kns5o3BpBNjtD0KcMdZNtyrB8JTZDYnhY/1LME
fUFaPHvYW4lLVD6bLQ8M5alGMz0qpdxZFVDH+nED7C5udEE4cZJFDSGpem7VpaE9AYRud45aKtfz
m0DajpLut2VmC3Z/4IGJjcYx5kYnXlnd8Gta3JgrY1+wf2VCJ/s25OJ/0gMqXPg408Fl6N686EEt
rZtv3SiC8dt9QkIEQrR8P7XuDsL+JJQn5pz+ddHUrLXHoGXN3HhUWSH04dFDEXYmHq6QEYxUQB+q
lQoyijgm878SbNGCiWo35S5EfYkX3i9QtQ0EnH41huGFMrVKoQtAz/fRpLEXXLN93e38bAVjC+YO
sDmIKgmCK1F+9Gu5H70eimKX86qxGEJK+H1jTFptzTdr084/dtxKQhqYqi4ONfPQpUa5e43RMU1G
12glwE8hK6LCPyWk95Tmkj9nQyaDbtWMbRSxgE9SUSzlH9qkZUWY38ohBOkPhU5tznj591cRYS0q
3YlqSmUOtSrOVSOpkn8uLCcU2IKoAqDj+6gD3gInF88yN6ni93EsKXS1ByAnUcbFTvlVW+wD1qR8
jMXstv9B+BEjikxZXNvQWo+JGOFKkH3z5+tDbxGR9w9vifT/intNtZ8mb5z07WzbPB8C6Z3qZ+s3
p6WKaWEKkXpJbMFZBDUhn5kIq43t8IPaqkcx+IJgDxfiEkmpzXYKwQHUxY8EqtoindWUKcMJgObp
8au5EooMYfl89PJBg3ByXUysYhsXSWmRFqlTMVvg3GFZjTGWNtTMx0wZ7Sf6XKG2ZpFRtCb6OC6D
aRKVn6qa0BnGOpM2GAbW1na5zjfoLJ/cLOwTM6wjOGKrlNHfkjjnLJ7P5YmCkM0prCoKlJL9ASoc
9gajRiOzSwWdTxpvEVMSie/mPJw/lQacHDrW7SZGBYrE6qGM8OxuPoFxHoheheS/snCEIKYUzXci
cwOtlPdq8rhkbK/Tz1GG+FvsOZ1IbCCOdktBGuxdpF85lHDv6KJTtOzdp+9a6wLJh4nl3mn6uVFv
5HYS18LgbI0XXiXeBxoD8x4RL9e87505kxpdpPUm9f6D/yFV8C1zzHalJZR9wofWPEGEil9ltVoS
XwLRj06a8J8HVTARn7itrIW5MXyQifakc7a8CU272mdACQIvpMdjllOt7OHtS9QlFSGF7Rq7Lcdt
KX5Zu2EuPdDl9TIlEITY5nww+DUJYvTtX63gj1ikcNjdhJjF1NWBeH+W5XMPkiD5SkHx8uv2AKVh
Yd/FfpJtKfAHc3Bjs9IMAwLEgD3VQ2uig7yzMdWFKUPkcwYTHPcQ3RJY4PmMvlawclmdfmZNOZq5
3LtsZnvY55UsoSU+0ddUuqXWnPKSKXqx20aLKMQm34UZNkU8WDuIqYnrNHM66WcpxQnG1OebAlR6
I+8VSp3cEcs0Wm9PnD/KEla6XdnXo53PYfH9Bnq/lx7YClaH6TXiqBkbs7GbzbbeFIGaw/0emX8/
mAyjvO3U/AbD5jgK7qxoLu7YL5BfbzYEfmJr6dtsgX0H2MhJXZsZOpc/QBwt5FYvtqBxhozA+s7o
Ny9zZM3TtE8r6PJlQJ2qVlqDTFwZapTtzb6qyEdQ0SbXnXl4OkR/T6WYFDCCXwddDQQ7BkcZ0MFQ
XmDMFPf7HmAa/RbyL6IOT+XA2efReZuvDe0w+xS3UVlRnaeh2Akjf+e2qrs0Cvc7y8l2CyrZQZ00
VZxaOP0x9jGNfkwOzKvyjzHtRbRSTFJwpdGnLsu/H2PiggsP2Z+od3m80lBASmXxvQ21JHkiqM7d
1fhbL2LOS6/fGKq1geTOJB+98luaAA33qnvy/Eo/BkK+TzgUxGI8+aQv+nK8IUa5piZKHnbzUfiD
FvIP9bJ+QSLAUVImf1F4RtUO6pui5Z1jl6pumDNKH1GZq+nfLoADr2+vWRzGLLkIw99eNCqUU2r/
xkQGEudbRiKB2Q2Lgu80Mc9sqIuet6p4SeCHpsINuyMVcB9qSsHT6QbfolqawLLXVh5mJio8aG+k
A7OaUgbEnsZBWf1ec5rOsOJucnO33xUJXuL0N4WCWENb8214b7SVhsHAFH0xZf9PisgdGBiPqluS
ZQ1LCcTXxR4pdOkafnuHduQsnQLN102WoIH5yvicYFBb1nZTLk3pdmMqmrnEy9ZJV0SqznADe0Bb
ZLlXreinhh2W3rJAqFsT/TScOjQV2cFkFEeX9MUVePSCdKLUhVbBDG8INtSXhBMxqAcDH+xZtet4
3rjGU5ARoN38iSr+4pjFmxGpXPr55NiewN7XuS5B+7U1fYZ9qTa49fFQhUKhiIMiZb6eNXoV0Xjl
Rigv88oC1ESPdbKjxuh+tAAkFNc5MVxUV7ERJehOpeLlkuflbhy0K0fIPRpcVgLI2BtCt1PUOzXl
IeNARQlkj4y7CxQAc31BxzVrY+D/0lRmEdgP8slpJjZ2WCxJ7LgLsvIxeuRkvas/MI1cfAIcdOFr
rSdVmiMDe8q2hTn1FcYZl7q0bju/HCFA16hbRcXSQya8CKrmnhvPsMk7FEH4xNYV3FFxZGoNe3ot
1Z+CHw/joJSYj2nF0McSwuLjrylABrJl5L/bwz3unNA3j+pswPPgFOa1RfUqIuDlYtf44GzEu3XX
cd4p/4WQ29JJ5qgfgR1Hw/1iPQNb3Uc8mh/17cX/PmcrjMvyJpOaTwETD/WjeswIPDBgbCOrrAcQ
pXN4F0W5CSDxT2lX3u6vo6YqvcJRZ4LRVCpumXhVLYERDTUOzVBrXIVx76PBiO9BUngWbW0o82mT
vmBHDEqWqkXt5XHxaP0VgmI/k3IzVz6Jx8NRdNfHk3zgtgKTuNpdAJX8YJkk+bZJn4LLHuxoxswr
Czb6x6V7tkJGr2cIZ5+kd0Yx2fszDan/Mmk6f1Dg3dD2fgTRdkksgm6CVLEEHqd/ZVDt5jMgbDKE
FWFYyhwTsiK7n7FioUod83oNpmZtNCGyBFO4ccSWJDj1vf3FNtMQGspRNhYmgfTWZPDzPZunIj5E
9rAjz+O3SFdME4TzVhBYMD8J0Y+bjuPtv9aBYU6z64wR73LihfeFAy+2YI2xcglrrXQfpd8mZi0G
EbumRmgJQDY5RUUnS/God1f931b9UJZ0tWzSEby4ucxpJNc9DGa0r5Fj2uUJFGavmOrAvaPab625
HC6w+geqmJ5Ji9rfThA8LXHGuvNo7Hk4Y6nFXsvUbfn+/SW12pjaolnOKc6ukoi2ltLrdAxybU3U
LnSMVkXDMUWF6WmQISF5ItwFkv2AeMy+xA4xQZcLpCGhaib5WgS0h/cyYlsLtg9Gyoqb+BA9r7GA
UqcwC7knI8Rl19OSvZl/38dgZW5EilnjBb74ZuI8YLqLYokL9BIwEgi1dIeb04W65kf+Q834Cr/1
sXAfGRFgOoPkiyh9tbMc9flDzBtXs1vj3+TW3uwr67CkBVy1XxtRk5+bmFzGJcOmUKKQ43pBJ5DL
YqV37/gQmwUUyAyg9LWifsCZ4Ie1mr9wYcgDOKwrDEVRUrmZdr4fEwcZYoBBMcShp+P9IhrhEics
vgcBZr14p85tKPPf10xfGy8t4pPg/mutI/UtQTLqRGVOGn+6dIu7ykLgJV399zG1XSlceUBHOIks
nyw7ppsP4cEdEaUPuJ+OBjzZfO0choTEo6LXAfaVr1ZTn7hHJkcu5ni9Y5vnZcVWMB/6kyNWaYyM
TNQB04ZXEpgsq+db2PBBiolvAf8D6N4B6XRJtUmt4+k/y6tdMWVoYSpUPrdkY87p1+CUTfxq0xsz
+okrFaGBZ0kznbDOjX48VtZZlJxV5nWFesVIMixxi7FnKM02y8Nnbi8IIHxjgDHIbes0CLb87ao+
kmBEWCDoh/XO8n5HZmuwMi80tEvSgjSwHeUAoD41Rkb6fZTsiCGsw8N+fciq1wWb6lvSjr6HjlKR
HvuseMwnyXXS2kaH+yweZePxRlF9DsWtGZZ4dkjRMPxMh6xFGNFLjWIfNKkXZG/Q2ofl7Drv1J8n
pUDf6s5CkHIpLynL57F1j1fid2lSUoxL87qzo9HemFQZIIkRK4/rTWz607DcST/64rn5a9ig6Mzb
cBlmMNWwoJb+KX9+He5MAHSvZ1L7YVumFpV94jKrc3WubyrnwTE6TCjR/35jq63yaAiJFg8hyuH/
jTxEw6YStiXGfiszGcmxZmUYJbNpcU91Skz9FYn5JjecslhnlKlHcrfAiCVErEHXcxSlwsYcpTTv
g7mbukjHiwIW+rMi+RIDuq/ENwqRWQWtRUsqIEn8oKK5d2hQPTK4iDbn5Sbvfouyg/CvQ71sSLlC
98oE4ZzOtaziUVQp3Wdck+KPWOmtbKMXVIgjKU+ah9lIEenkia4WalR1r01SLFksEbdK9/G9cojL
HS+ye+zVu+ZnvpZQRRlw3fgxeun9HcV2pUw5ZdGw57ojoszS4ccnaPgT2XmMGCyyc53FYovcTGx9
TD2vU7vYQw92ya9SMg9XcVmnD663t3RnmUQIOgEn3lKACzIUbnHwLWWLkWEWOYxlBSSq8r2ACcTg
MFZfiiu9+osIdka3nHA/OOvoIIMHZwZIyi7G/VX4RrkuUFPvUyv3zAZ4OA5CXqqSEAP/E8T4uxv4
P/x1ppIS3TlYPn+FgqYbGLE8ahfUq3bTIDCdIzkfZ45GJNOBAwIEZ70OgFInAFGLMp24x8D1o/NK
znQnpykQv+ccofxTCVucjdE52U3DjRqnIvBIVyULqen2nJ3FSjKJsaDm2BmEig4vp9rxk5exS4bm
2gYZBaIjInkbCSZH+DeySH66bvWkDq/GEoU+1RkvqVysUn/oP1z/ySykChLfriNl2oYq815zALVX
/c/NHDDKIW3uynpT4+Lg00/Y17CLn0RVnYbHZrmzoCmd/RGX1M0cGjqgifUsx0h+QeQG55vf6/Ph
lS/WN3Qci4gVo74R+4cSbjTffyRw7L85ZQX5UZ0otCdaJRiJTyiTre5C1to91o4y+hiEpTsYf0mw
0VdvRm/cIIBrvoa+SrkoJqZbNFKC1q3r9KylJk0s2ItMC+SsFa92tqD0ybjEaXFujFiDk/ZUMJYW
eGNbhzK9YhF07MKWZtYYl2HIpF2eQn9abYynHDMwrDVTMPsVMdNbsAfeWA7CzJmS+MKIFTKLawSe
v5pUXeWCNeE7AffhoQITvS+fkYbLAcgqdy2mtDnQZ84hPL/JHJQGgaTVj0aWpZ3WhPWwwCn4NZNN
B6u0d+V57vf8S019Tlg7PeALhjpgGOoKs8E2kpc0jNf4tnXXmmQVD+kIX5oiFVepMr7sBal6dXI5
49nGKNoYrnHLthH4LOaX4jzqTWldH8n+v0eFdbf3fLpLJ61HBOuvjeLok5oLnbXfIDv2ypWbW1ld
/iSfdrMwKrMfBD8FiWWgvv83XrNsf5FWK5qIudafs17XYDa8jNxWjz1/HCy4KDoZlfD866jwLPZK
w+r/JtveqRFgbHYjftIqJnmQMemV0nuX/0c7pf4s4J1wwjvHPvlePnHZ1tMfQ9/rcbPo07r1xIww
OhEambLFK9okqafDy3FasdZwGQmKeReUgpyGCn/46O7v74DhMrktt7B/BH3+ygJbtVmqEv9QBgCv
GkfxG0h4ATuSNT3sPv9/ajtCSaQ2Okg8upTPkM3/ftKFCkJi5MVATclJIlPGgTXLH3aqxiMLqJWQ
H6psRL2lG7FwpC45KlQTgj6/T8FE5DT2o4vTc675R0bNJSZfWtaffaasVmKoQr7Ln3oZXJNmOPOD
vH8WSOeooEq4njFR0gqG1RH1j9UHuteHhNALwHtq8lTI4t4sVOMTRXI9DoR1Ih0JGKXifeiECnrY
Vec3EDBOsRSoCc1uW646Wb9sQw17CRQ06bRt94g0Hcqnifq8RTA1OxmLS8PFB8WFQTi++eVTSsl5
Tdd99mW8GPYY8oBJqPQ2ZSIJSIUUruwF+zOKLeiCOgCJICtNvnia7suRT/nHgbcZr6tr1KjgTMZx
B1LPEklTR0Krv7g9GBfCCgZylCF3h+qt3DPclzHI7HCeLtcBlGtoezal0dsmCzk4hGWRmxmXUFIh
KwK0gOUBRC45MXFupvMshoIUVnPVzAoDJ3PqOfVK/GCD03yTZWH0p2e7ikiyj4s0P4WN3TST8pwd
y0a+28CBVRK9ZC0rCUMucsrd4Hf3kRXGbzWwtUak4ySg9yDD6Y2nfj1cCiyLDDcvdbRzG7qv/18z
IpxMmP6q8FkTA1tUEoKrLjyEwShCzXauYtO9YRGzL3cOjZj/bolupjJJBVivcKPuwhhW4RmU9Udy
VcUzCVJ6aQIMw4m8cx7ko7np0N9NETlNCXacrc3Sv+ISwmvNmVoyXFquHceWhjZEpikVZ0XmyXXa
/7t/3zZy3+JjWapFLOpv0MfcELPLqJEz0LtY/glKzsQup6kr9tNYgkCYYXXH1TSiqIVMpo9pP4Lz
J7L0CZh2IxJqpT54Gkn1RWLP9KKlcpLLu6I1cUBH9887+UNO6gNHag/a3rDBE4OdQQHpAT0Trq0f
nmt5cPn0jFbQ13B0mMURcbZzDGy49c8SWg7cCe/UEVYUpJb3My5UB69umqXu3zEdAfSXIWWxzKvJ
7D3YO89pJpzZuqY5K82CjAyH+BHW7Mh3I6pIyQjEIwF97A7dVCA5JPizCfT3jaLES0+pr4EQPOil
Hyw5n4J1nVLfjLpB+mw/trT6m+m2rGj7aNtrYAT6z06iYxNikICV3cQsnXScz++4KRn4dqL8bMZN
D+jAzkfzGYdy4D4tI3FtIda4ZxCFEpzWN84fq9tX/I+OcPFckB84CDOzWYSoUrVp4Zbez/Zea5tq
b779JNr1baQtGIHF6ax7nR4G9W7YzkRcRaoXeDDWzgKgum1Ujctic1bkZ20o+2Hd169abiYLoNJR
rswZfhHU6m2ByUO+u29lOmYnnPQAUU9EY9hMkTyH5ftjD6soEjLMGq1x/nK/4eEXC7eZmxvfjsS/
AxmJhwZTlL++oUcL2H9MIu+CYyrfCNqMo21caIwyU5WmFRNbXYazHKBPEiwc57ITBGND+6KXv4tv
4LuO8TTSOFTDpSHj5S7rprDoKGHhm9X44rzbqt1yhkhwxt/kg0ZdZ/DJDU+HtdjxIsmCHUiAcgNd
DMDITE2H7oFTZyEb9lM7Ui7l3xHXHjb4Lk8OCAlBgrt65zzKHDyxdddm3iY7TU1Z/2CjzIC6v73w
avAGBSuVI6VoBt+omkY6L0AyH2P+fit17a9i/k+Fp9mwB9Pm4Hm8mq3WqyvT1TcZbC1ECih/iNUW
Ng0cIb0Fb98vNKqgelcX7lBRNCOoti/RDNZxjColrJ3eK3FiJ3qxziHI3ic99vCbjmoP1tOahpWe
6XNz+BubWKrfIsyM5BJ1R1m/hGBKxXGC5FLa6b+YysftgZRWSgNVH/Vwk6Kk3MRe5tohCh8EoYMU
b2Rxc0SO2T1jyB4wLGri/3hOVt3QKPDcJ7GZQgGB3LMH7MAeUXMv3yM2RR6JiMpExjy0K9dRQJMr
wQiG+PDIQe3A3Qp+AKvXm2Olm/xzHQ1JMTHeeXOFzCcMkiS8VhhdgprxDswnc9uHplku3aBxm0GC
MHfSR2p3j2IvODFig2vRd1FUZ5MMD0WdrCs/fY4SP8Cce/GwfKKUpXFcL6VVNp0zyBEhjnHQSUeE
atZMg7RlC4hvUWVMA4nXPLp0o5YUhRn3cIgO8QxYyZ22QpK0q1VIZqpR6vxxGedCL/0PUje6oT0Y
m096vhDjuvLo6Pysf+hvrKKYYjBaRzYFB3IavEjaUMofO/VENSdrpDxUAaLqpChCUxmxJldDTTPZ
P6YaWs7yMZaII1y2EP1pLepn1O01fDyCn044vt5R9tGGe9i+CqBqbcZH0MP6MnGlt3iEOKUjteWP
z76Lf+9jqG2MKUkmd7tMLbvjTUsWSp1GykkTPcsHL5miAMwNlYoEO/9FcVt5iYxcN8RPvfGr0uGM
8jH4WXpbxgACI7Hga/hvJ35B9ihIHYeueD4Dyu0ciS/Cb1+D1fxPFit3gXPHssZoRrMWfyDIvpXg
s1Gv0nvsoy6EP9sXzL6DhbalTKoy5D0oFktZcLXJTFPagApGIBObLelwiLGFzBYccHPfdBNk+X7c
FF1b0tIlltU5Qki6eJCr7tfvnukBUX7/uEVMlv044YehNAfhOQ23weJ2mPw2YQmnKNHy85K6r3Xl
aSiCfIOqM1fXox4LWASLgx2maZQddMssvxTTiCbgBqtTbGoluVJWl5wL8mXzo2SbHh/aRXkGpVM9
1VMxtArbg3JxMtxpVCdCFi/u5FYXE85tmutr54V4v3kUwVgwNh4sa3Ev7MD1gFBqNyFQDXqd8fXA
UIdL66jLxRaiIEKqnKDSUj0FzkLR69FEExFkIW7YTDjFCI3732kXur+4KKCgrNf2mYANPikAOICo
nE6fR19Maaq/NB8YkgsoCV6Mi6ze6Y8o3wYQyo1fkRB7ImlVeZnceZUNvUPctKL0KKj460hpgCjT
nFrotooL+gC81E/mz40Y+zMpjs8mnX72MqcS4j6geMnpAiZNxZPXKvKPJTvwWF6+MECynPGvdd7Y
A1eDEOPMCvigXmnikC69oYK0P0arLEVBNAnVg575GC3KI18R1xn+vuwABb6aaPzxjdFVhjS4zRmM
ZyjetdtGzu6+sCM53otCVvV2r7nYHlw8IuaJByDrUPgP3c5xNUcB/Cp1bjselESCN+C/CFmt92pS
FmWlPLWGOnaqYiOb1pMsPq0GaoAYgyAKuqODgt4WigxJOQEL4sp0P+6nv1tM3lIT3dTMrQsFvbhE
5F6+sY0Vj2heVjtv2Rp5VDwGBmXJZJTlBIHYtAoYQ6MJNP1BbMoXPTOUar5YEh+97NUZtp24UYFK
eR0uLT7M1TW9XCRhd/pc3pesyjzcSNr5a9cRnFUOBgmfhRIB9e9lG91V38g8YcFzOh8dS3eYFd92
Nbe7U+plo6FKAcFdAZdPz91IPTgjoiJwE3vNGMa639guv+jX94kIWB38tX0n01+aaNg/Zo+riz6F
LJpUL2sLyQbtxfvr8h6mk4LG8nc4QneouNPE0tmBWJhdpFNjgvNo1NhI6XCYg7BMWV8QHV9elTRU
uILwOn8+j/vhO7p34cRijufTD+m/I1rHXUc6FWS3wZbaBR1fOiAUv+qOt00zJr3Re6hZ+4YBoxt3
ppj/zcTIBMnqfbwHWiOz0tefuf+Dtt4n32TYF3xujFdI0mRIH3ZQ2mBs5X83a/S5UrQNoGYPaqv0
dJSQN7/s/1B+ZCMewvfhCYjcbcAALWGq0nxdgsGZkW4RruLIFh5plMiYB8e3jW4lzAzAtjv/91lV
MjWoIKY96mlWF62HTATwj/W5etPLBckhBIOYeg+IvDSGQJ0lqCShvWD0CaeCnixy0QTfOhgpZrn5
AaDKoR2ngc+3ff/XOvSs+xFL/zzsWAMuFFLg/1WLK41SpeEGYmrunaBsui+8a780lcsSOUpAERGc
KUqgeNzPl3i4+/WJ/G4j+8Fzrs1fnpig6Y/fqGBVHHvrqNbtj7IghlfHJDuNp6CvN3oGnq+O0GeP
9FRD+8l+OC4CPTCUE+0Fa2rXubaxAjHoJl91QupvvE3aCWJ5ZWpRXLooEBNVBMKrVGlEpPQC/zMy
s75LUoZ3ZwGM505tCWXGhoKC9WoOfz33OmRsdtsAi6hv5Yz9GHOpXiGY9yq0qSu7Sg9EEXEH70Ww
CfVL6rzHUMzThvkPq4NNNWDooVXbOb79tWcAx7wqp9uE9FL9FOxwB+e/Rvj2+PtyEMKXVfdeD/4I
o3tyE8uThY+pTpPXukW5SiOF052G7GowtLP7qBpNvwZOXwwWZxDRrOl82Trpoh2oF3wC/jWedRE2
7LWWOXP2jvL5kgrmcuPaFIQnyxpqVGBCFV6RLARJu/HAa5jZf47t+xN/b8cCTKA3MNoGCN5abmAw
0sMG7cpGJ5hEY6h9RR4c6YPAdFOTav9i9cncAA/ZAkx4l00w9WAVER3NaqnAcPcLt1PwP2kBJrHj
7wqyygWSY9xvFksuuyImrpdjgVfpolLuJezwmYT3Xxrua9abQP3BH+72zLh3/85MwFMNTIRfS6tf
YOXbg0vWsfLxK4a0K+0mpzuftKVEhoV6plOGQO3RHzySKUXAAJ5ZVuZJY4ihZoPlA/HuIQx3xwcm
T19nwwc4Di9XvF2Wt1kxrUnMp1XoUd33hfQ2TmucTumJzucBbSQIbcZVHjf2ojHVGJH4gsDH9IDz
G0x2ZpOroRdvPB+ISdy/0ih7Q0Yt9C+D2qpaPFN6bRmqUfu5EKscuu9XUbVMaG571tKQDoaWJ0le
iZKN500/UViQQRtdQfPTVv9bL/O3LIMNU6qNk+zwpN1wuVbl10cO2relQgm66v+e2ciiqYRmk1DT
LvM41g6BlF4lo8u4fRKVEz5ZNKO+m2W1eVN5sgCTQr/aTIZ4Pu4LHEWFdMmW9ecWkXt2F4EBHsHD
xk5cDr+f7SjTkK/ZPGR/X82XTS27awE87WeFZV36LiDm7+e0/89mXNJdNtZ4fKUUwsMylAQQ/FeX
mrR3MJB6/Iir3WHEb6+NZhwl6sN9e7UWFgLnnXrV9HV34E8SinIisKNxHYTSE2wmds2Wvk77sZtB
iwZGd7JwN3NbuI/OLmB397POVQf1iD+OBgZZEO0TphyDKauXYphZqVxtZ3aROnLUYRkL4sTzX785
ti6bzKMpjY7ekSeQ2QGw/GjrJDwIIrMmbYv9mxiYcXD17DGdfOA+Z0sbOibwtFTg6DIi96n42moF
Zss0RlJwtvoNyRWPxPhLE75lfBIkiMCbGwIhkcNu+k10GMSxOXFGiX9YwPYLgLrOJqNMeK92jsbl
FmKo813mPAsJVCoDuX+pPDiIr73eD0Oh1txHqJOkLdt7new44nLGeiHKA60shBhQ+FD0s5JSKHCd
0Vf8Ly8jpINmEZfkMuej4UZOrw+BMRrwOMLscatvj5REi+TUZmPqUYYvu5bRNNLPXQ3H3nGc/5bg
NH9kQXePUt325cXRHtxcqn7kPCVJhcitIgTw20bQxs+owxyGiZkR9jqxrJG3/jRJ12AmIm8Jepfa
DVGfa9OweGZ9GPeaKC/7mo71SJvULg+odfEMb16FwW92zWMBkGakrTDamoOIDl6iTy6bNBmgu9JA
PunzsDJWya0iiGf1luzdaWvoDhUUrht2fNq6k0IF0x0RLtbyRPikJk4FIWdtIQdG8Tl1zZn+W2gx
FC/B6UDM5zzpY5w3diENx1vK+vivpYYCfGxoxLATjoBb3hxaz0/9T/ERCT7lUnxmAUG3CPh2YP+V
PcIZlVvJFJSkA/oyVaDujztc+vnbetYSrPmOyS6zaS1BNVH2lcoJvwY0zLAvAWd+tAeHlGJn0Iio
ZTv9Ok5zEThVRg8FdN9sNn3dgwqeHZmITBUIWcVrodiG2igwLpPt9Nqyj9wjimwvqWXNXanu/Fhr
R3rTzb4wCRlSn0uMZxjImRJdDn4VXWcSqb+61mHs75j9mvR71o7yzpmOw2Y3fLqrHmrgVqTqlcOW
8PTA+u+1XXZ/nixH9J0zERuHeVJwgUcjtz1i2xjma65uGrqu8AQ7IwwwkE/vI99tdrEQahvMZ4hR
d16Uf1jbrU0DsN+jwOJ80J6Ou97fnNuTCZhsBzsD75AZql4nAmqRb9/8TDPubXAmHdYnC7Rx57IA
ERojxyaujv2bknx0zwwxUVcqZL1+UUtO7ztAlNe7lB6MY7IikP45Vrni5CMmEuoTgF3L89yUTDKv
9tKkHDOrhhrhTWOjDTSGiungi9dn+pTy3OMa0UqTwtJSnRrRjSg3pAUYHLWZ5EP/fzcjvPv3N5o2
RWHNl9unOWFXWDXS1mAIpJlM2ewnNAgMD6ZWANg5yrILajVLDSD4tfzWVS/3ZZ1ASqAqZTa2+C5j
kmyfZcIWIsI7Y/68QkgBb3VfLHHef1Xnm4TJ5r1dVeD/QM2vOpZt1+qSoHBNwTneFBIyI2MWMI7R
MwjpqwKgRlQfRsttjGHT99e9eIH7Yw9ip7Jk56vfQi+S179oCKN7vdwHrO+HJrXZkpz0Kdqe/6JR
DJmYSmG2J0LzrPfMfTLe3Yilu3PRyv3+n56d+XqFcnmXLNuLoMgIEPYmgmx5VFtB+A5Y6BTkkAMo
FHmWTZAHuuqNxcIIw8RMvSyw2P8e6KdqzJErtQQMOTClIFJUOAet18ThO8Q+YrjDbPbncUsqLSxu
NU4hzi0NgEMM4Iky20oWG8tNopTxUVYoW0IpuJbhcXzLlp54L+xD1y4Zyg2TKSLqLzpc3HhptRQs
o6ZhXfHiE8qrtB9T3wwKUtVZSMpjUGHa2P72GJ2Rg6XEXvoacM9HLRELEAadhzkJQbBmbUJxa5Ey
g/6K/Yu+FHEsvRq3jzNh1AzGGC7fmc1XCeE9pI2r+p82AvBpC/YSjYmyo1aqHBDzGiGGPaDodsWm
PAHE6YrO9M6e39GH3K6RFQlCU2Fah67uVHuO1yyIFrH+AuLtA6tJ6C9q/nos+HS81REC+X3ZvGuP
SccS8k3Xtu/aF63Y6woltz1L0o23ZJGBmMeoYt+njHjSpEHCyQDZoq4GlfaJpDqOdNcmQibP5SJ4
kmq9hYaE03+Sc/Nei4rKdogLV3zg9Mr7QXOIpRQ5CwtEINRHFO2p3CyofxIFxtJtQHzYU1pxs1FH
AxWchOC4GDTHVPbSqH1PQ55crGA7YwcvHZy7CxKHG23tq4yVv+tPqdcwCoZcYNLLQNS6KPWYkMlN
Ryrug+yoN8qqIpIymgMcoWpr+jsJ+Ezo9ZXW5LA2MnyzIH69/njH4Y053PTIAHOfnRgL8W+POWbX
6XCaY1t3S+84LcXs07yU8meZTo0YwR2EeeIuCH0pFE8qws7RKdvsmgdNpsJF0cREz6Pfvy0m6nLW
PSuegc+SqHT4I3g4QCRcaqosGhPHCYV0xpt3LcK6z3PB1UYYV9S1fo1pPznpn2w0EeqDfRGyV8sw
QmbmTN2tFErZ57Oc5DbKWbyqiE3+3Q/5MnddTdxPMWISK/V8dwt5fl82N/q5hvXhXk0yRxls8LyN
ucPI8j663pHjKSkunrMNvSQVQIexAk3+eWlAV+K1AZ+edIm61sRbWkCFDRYlM8vWhUPqxxV6Bfz+
U76QeoM57lKLAHZ170+owiLQLZ7OiOQUsIj2raiBWJvkx0CVqZPv/LG01JiAAg9O1OH17OwZQUDO
0nk7xzxIgnJvyEtZGwVPnUonUbNtlSv9HweeBZ/gaOxnNTUSAJ7VYiZKEa8FRR5wHJmwQ9dUjjL/
8a/tYtIhRuNjmOzVVzzQeSzo6c2rgDVVl9OWLN4hMglj6obEQwUGsw+VH4o3xKAvj5tz1SF9RgYh
1LCTXDowk9/N7sQTn84V5PhaZ8PpfAdmRQKC1j0PtgUYIBgQ9IYqA6+MM3PY91oM4IdH/qx5Qf+M
y7GQF9IqUvxQqLYvYCckT7Mc7uRu4xN0jgOt8TP1NKPP34OVmkdyK/tHQLVpfNOlnBEl7ZRCgx5W
CNiMr2zy+LU4jeVYQY6UzISP8TEEu/xKLB0fFF5uMVnVg7ClGCg4RRasHPVi3cCH/2ytIPSAn5UY
bbY2kzodh1WWiTOu0wZAZ9ndlloU60l6cuN8+Gw/uR9iM4h5e6NTuBXv9WqYnlETuAMt9vY93fj8
ByJJg4Yk7Bg80aRx1r1mCR0rtPyFzQ2ije7UXSw6AC+hDTXk9dai6Opcly+sKzO9Ke/7GUEWFyG3
ayfU+MYrmoUnb8HBdbtIQ5v4ySHtRxLGKx+iR2WAvktLqY6HZaOQcLXjR+ruQbtg5K+057vHLztq
MNlVWqmuYWwtasru1cObCe6DmyvNJIGzStgbYzzGGQpE1rnQv8z8qweSOz/rbuUx0qgTu5maYvDf
8qe9gkNGerNE4OC8Vno+A6yeHYEAVy4B7vETYlNiGNYDypEI0BFDVdmqPO+ozNbwp5aWA49XanoK
aY0qxtyXmQf3MXykvO0YkzbhKfnd+yNvvFIwFbIj62rrfNBOteJxy+57/gcOzGujfedEMbwF5Sc3
9L8liMR9Tye8lkqolV48GuAju4shNf8p4eFiyr3y5F6G0J6gjNoigXRO4+MeYS/KD7D2a8VEoOhg
d4TQFy2Rc/jU9kAGrLJIxyP21A/HvIUc+YwpDX/0siGEj7jtPMEWDsVpkIHGGivkTPgW27MJlZHC
u10iv6nztBWHH97MkiM5olZHQA5X36i2eNxd7bdxRsO7uOxf5GqHefbSkp2Zng4vSDkrv0bx36UN
NM1IRdExCQuWjWJEuhM5qhmHybYdwMIt9iEcWn4RYLRJXje+P4NLLYUgi512x7ZZ2VDopnC28QsG
/DI0RPXJ9YbGCc9qy2ZODwgj0TTkgqTuv5mS9E0ZypSgjqFrGeT9xG5x4B/pPuXCEXSLb/kTJTWu
Gibcch2EuVO+LUMQfgC0hkA8JJVmI91KxhiHx4OW8LZAnfnS4zVM9akldt22FMlYvneQctyxcypf
pg7QHLIUXKW09t1thyfs5zfbgxo8mR6cLxPWT8fi08ZOdYCmNVeYqz5KdhpTufiNAGxaHLU6Ub0+
xB5ecEGcPf4QmCNn3c7gQUIhuM3f1layG3RnhkBW8zgUhc+bHfwuit8F5cK6Pd/APZHme0Z4QPOv
I0fDJkaa9oBOdtSZIcjFCUcbcrzTyQVG2i5fvp2SJqT+yUaLnE/HEhs90f97XFp23FQyD+8M3O7E
vxWAr6HxKbGA/OrpWSxlhYUlPMgmnAnFV/nnvWxABElxfSzTmLmmBG7AthsTMYnI5ptQiz5pXkyv
u/G1ugVMROPiW6CLVO8fZTcfz8p8siVt8mwIl5M9veiS1aOOOk2kGYfB8vLrHEyIUn0PsCrK91hu
aiVgx8jB0gSqi3rDHn5ni/e+P+aOD3dbU+76DxKneqx/XCh1zuZZnGhlqq+h0u5tAsQwt6XbWV+p
bUOcmi4c2iU+yB11ejMViOx4qHru7cQsYloAyCFmdpUCyuxiC7CjjfbgWsEx3xRb0n9U+r/2j7MS
LS02LYMl3edb/3+rKe7HPcFxWDdm19FLwL9KQffFvvupcqszljQUMCQ+taxvsOTp0ga/DNc8bPc1
QbwxTTe/rdtLyUj29A5cIb9/s4pB6RrRz7gHlHBtTbw5DBe3YKaXbenIilZnNLdxKo4+maM3JUH5
gzBpV/pVJGJFb0TX8C9VGvRS+F+QNWZeTBL75JqTd7JSsPSvB0fGQHpHRz+s5wzyl9LsnihlRISV
EJFofIhz5l3M5lymvwUgkbWXf99Mu/CgP/X6mqtC31byc9Sv2/OZCT75ncaQv3csFgjx+vA1Q1xc
kUnXO2QxfHu38xzU+GjJEcGzg+9+2wNpeMbi2rvoq9Yc72BYNy1yfQVsZNWyTrvr+sc0fVSCFg5I
CyVHfGPEY0G/vqRMzAdmP2filjHKQlmckrW4jIhHTRDf4h+O48C5EQPh3i8fXJu5N2IVYwyIF241
uPKHHHdRJpFYONLuHlK9zm8bjofeIPQ4cHnoM19SDH5nreIZ9jHzwfkjy09awEBhBdiXkQD2pTiY
w0Z+YuDOu7Q5r/SqlCAsRdVuRSnFSkD4lul7ARSAB+4J1X4Zm6bsmW14QI8dJgYLmlzpMv8fCyj7
ng+csxu7EA+nWkOVxB+PdAvdCs5oYERHhu6mo10xmQljyhgejxOkZVAwyzZoLcOrTyTM6aHTxGnG
rFQQ7Mi2SZTKA8+GcI8/kobCzUAYDZ8zEMBDSk30wtC2IP8CCyPNMWP/zLRWw8wQgaF8O2Acgz1g
JqzAvNgrQFuoGTkOxPzHC4i7NFp38IMAZbsQIhj/WdR7RTDbcgAeYlvjWzQKOWUaYrVC92KZxRBO
IxZZI0FpJEv1tmec2ckvjGt6EdNRl4tORwgAQD962RSSaj+AeDRpRLDizdjxVEWtaPZuCwRP+D4U
obBbRkSrijS+O11FVPQg2VV77Dfal2ccsYSG2gC6PM5RXEOvO7bQ6lh4lrmP/MRg4xqQxd0nG+fo
HfrusaRaRqATc5g8nNZb90yQLZkxAgzY8HDZTWCWBqlK4VRHPnRKib2QMuAfi9JVkI40aYeIwu2S
BqaUmPTA7l8bCF1ZffQLN0nBFG15m0/jH0iqTT4mpEBiqtrr85Ayl90DdCt8qoOVevFRSzg4BkKQ
a/Tg1l7badHnWhdGXLhCVomKcZzBgkfkw8MESuoWS6zDvKo+kajumJsHzU9FwGqV3bhxJ7ABnYxW
Ku+vLGoKVFEjYoEOk0r8olksw7+aycyOs3z8FZ7+r9m8YAZgKbHXIQIgSjkELQUhu2zL4yqw6f/5
SyJoTMJcL59H2Myn7R2xdrWC9ujP+odxBkmtR8AdHmDJNVHrfMoW0wrWca+QK47eNpYE1Jspcz/c
EYbfpVh4hxhXlz0fwsKBkqNGYHQk7VBVsZpoBGtw4UBcxYi+EmHsYHZonjowI5axPJcmnEmNeWGX
at0Rt35w3MGx2VrrjwpKy8lY7GhGJeAvIespfXB+P5BSLPmFNF5zHBwCuKNTq8jlRCge5nzjZKrq
C2XgYVPB4j45fzvF0op4MnDooqtLYXNDWJEcFuZyOOaIzTSIxXArmsb/RUb3YRgfdl8f0k1Xmzxc
H301V6avi0rxHpUsOfOuvLJf9HhjQKo7R51AcI4IYYgSIKwADC9zKZKQfWzUSVLOS6DGYlsLhB/Y
FmJGmT/q7UyVyQS9x33tTgqgWwIHfXYI/sFFkmy1NzQPNaQKyEhPHlKkYUgtxqbx06ISJY+iDx5d
n3bDfujm7slniv2kdQx/8COsM4EU+oOK0n+3PKwa3d4/OaYoUGq7Lg6SGuBDn+zMaHbogOrhYe7B
Q+suzg7EJN7jcMGeBt39jHeAuvRT0Yzs7vgNUn7A2GDvOBbVbiQDMlyIZaGNTg0uv0Fb4FapTqZR
Ce7aHr6H0KUdWrWoShpuZPJEIvV0tbZoCSo7LWTulCiNr38fu4xJ+zjCjqey8SmoTLzmyQoW2zqc
gpgIdTKtcGbjlt2ZLv8rYhNHpPHQDT4fLjb3tnJNdvn6SbH/nXJhqA0+QS2B9E3tTHD/kb5f0kfZ
VTH1TT6kD1QjoPoVE5vY6BlBJ9fs869uplo+gLHovZ8ZSsK26Uhl+6hci2X3Y8DQEWQLiAW9lq/z
8Mfvh9aJrHPqIqNgOaRQyxRLB+eLANsAYMgEeOMUCy+TyqwLSFm1YZiBmIlSw6y4OQc2Xy61WrEr
63VLkuEbDFo2UGwjcWPWEkCBNBcCPgzk9gMhOxwbINd8WLEwHE7+YFRwGbZZmQQUTdZXOoZ10JU3
hvTcZ/Ann9gxQJ3DveAzLhzBP+MQ0mEHcnJd6JG0+e3tIN75HYa7q9CXHXZkPgRjWI3DAuPWqJ04
iBTa2aSH5/jnwGGml/kGCwvVLYztHvLILkotS2yut76SuXIgp1yLeXmT9LyXCZeK7OrGqUERgkMj
Qcjd/CDM9z1B2FM6LfuiqQbL3msAwqiZIp1Y/tVzCpMWw+THJ4fGs/DBiyi8z/QJnk9Z2gCxCqGD
qgnGJ/WohtSSRO4lOSBe8JJQ8buOljyAc+7eTrcZZrGapj+u/jJ/o6feRlE6pyAUHBZ/NQM0HlP9
1ORyT73nzGaaG5BhHFvFQIIWX1aVYK4sfw5Ud+KUVOKytkkKXfObL4h1sOTUT2//5CZoqhufrRGs
feP4Z8rqW+GbksdyeHCkadf93cVBHICDmnA2lwHCWuYfjhOect2QFxOFo3muh97jHyaN7vvR44qe
aFhRkFHZiM/7W33qFHLNb501QK4B9LX9foZf1r3HrtUSLk2ylGkHkcgCHwDSc1cGw1L5t2iJ29yt
hxkY1Ra29z3q+QfgAF1xVYkYYLbhHGz8hCIVJJVzG51lRqq10iDRCsSSWtHbdcWwfpMYBP4mCsnz
cm0AjAeXLNebOtgLYIv6bwNZ5KnZdPBQ97RsPYPYsYYGV/hPKqGdsAowrkoOsTMk21/AB61ivu5s
J+Lksb773d6iuAeDARFJF9WhkFseaxm+ugu6Y4oLqdp97li4SfaQLMmTiXTFWRKne6sJku9xAVHn
d7ZY9NSSQrC5bGvfK9kzGNMjRo9B5CiNROocB/+3EQZe2CepPWBPGlLfXyZ2k8sCoXQW4JyepStI
q7+q5xXzs7I3Cy8vrh53WPCx546S+yp1ZYCTnuF54FcNx7iRBoK0U5OrtOuRaX6n0jgBOusD3pXu
fXqVdLSwL49oNKgenii6U3W7/QsuwbWNlp7S1UeLjE7e8aFfttZYdk74wyZgAh2eIwOhVDYbtLQH
9KaR9caBYAdPfflvoH13dt9YJ2EucSIL5QG+6S1qZijaMvAUBG5K/d4s5+i+J9/Gu+xhCgX+dJa5
wIrG14UeYPjkG6a5ktuZeMbww886e3kiqYq11WrT4JeyNLxWAg8KosoBF/7PrAR3675AREDnLazb
GP8X/gVfv92pgiYH9NVpT5rKPQjD1u3Dp0idMxKxjZBUWaHdJXdPffJsDA9LrOYXIREuHWvDdxWZ
edMq/7tsgI8Yy2J/JdFJ7aTOk1DsesgRgdm7YfreTuBtbnZpQCIDCImggnX7WDRXfuUvTRcRn/of
rnm7O50IP9dBt1OPbM/fmVrho85RVyG+3IliIZ3Hm7GCthxsSYYZVcJjqD3jarJrXX3pSkq8EzeG
Sfeqhr3oyIvTGGXl21lfh3lWkvKDgqq46BIOXVixN2TfICetfF0GcdkoC5Y+Ry34V+l8svpIgnRx
LCUoDihrEMVLa3f20SLoH4mCll5YCeCxovd8RC7qGsUXxh5JQYkzOSQj9uhKNCMbfbbXerNDvPAa
1nZ6EjI+cV312+TZCR6SInrneDnxUVYMMzZ81L8fUTDxof/s7XXT0yP62sZrQEnc/I7KbghLRPw+
8ruyysy0AvUhJVokZ+ETLXpwOcfoBI+N4NPyl4kikVIwJqXgj3d42CXDwAtCw9pIunm+K9LnTtYK
vAbpOY4G3jORXKeopyEHfSqgDAYA72bUILofRSuUo2/pRxBZ8eTnp2sbO/4115IFP6M9N/LmAPYr
51CKB0Vbo6hi06l1jg3fDrdTnoWr4vJrdTz+tFjT1aGTwch3M7nsO7ZGaREV/3xiDldXhDZuT0z8
76oJ/rOLfGuTgJe53f0lfdZAOaZBLz7vym3vDHvMfMEqmEjwLF1AIP6ouuOQAueekrpD2utvmHVX
Qx32XfZ5xr93rYRPL/bZaMYkKTzOqNpyzBPbIWXKmHPDM1AC2vFGVvYi3tWIiSXQQ62gYvMyNYVt
Myf/xHLUgqVBiF12m7pekKZVh9FDaqXEpIQxKz69LNfKEtGY43Flle98MBG9Kd39toppuEtokk5C
i8lhLk5k8Jn1gJgOL/RlXy7LGr5K0suj5CagmKcHt5yNdk8Wyqm11gP94EVKXq5ytoTYfX0lEglB
OCt8NoQGuwHkuGW6hd6B3Sh/592w8y22DBT/EpBz+EpXSSAn5UjVX7I1NEuqtD8VUloaLCdgrSvl
1HHb3yY0mvc+FSBGrX0Q8i/mit44ACZUSw3f4+re5WtezMc2x3YwWbowKZcsBO547ashZth5a4Ef
NQAwTWAOuoNzCmD2E4QF6NynzgyTT+hW0CnUVxJkhOZBHjByC3JT8eQnXqPjQ6GwEUgMD7hDkCKX
FlqM7h+6uDqblreIwL31J1tbApmjTlWEE39i5zaiAI8dsU5FKP3ywkMdWNfjhjRxTsgPSBfrrHXo
h73IGbkxI7OqyDrY0XMVwA6PzoDXTyxh7GHwzJChOJixrxFGldFbeVuBE2LTXyKtAk5bXscEa4j1
zOnW/blxbaHHWGTiNgQvvM7F3/amFGZDvDI+eyTFJLSwWsiEhbnRpU0jRtAhO6rJhEVSseuLudQ7
FGSDyzDz0Jo9BztoudltPSqzrg0w8Ihpru8ympiJeb/uqvWJl6utiWxYLqqQPgSY62Qz7PgbDQdE
ay/MRVM+pIzQs4OA4a1gOnaQ0XeigwyLEkdq0ltpUSinsY7sChKDkw+6jewkEUVZ8X4VuVYPfAKt
55H4EtW426cbSUXHte9i3pztggtLNfcSP0VjZCdlCDpKFvowouQhU2ZkxNyt+T6l2HYU2oyynRRa
2UmM4n1AcytH98LBAktXfHepv5kExnsqGE3iBuxusq8byc8zGT7DXhrTsk6/G8y9XxYpfcFfTIsH
U4n51H2i8Na1FcLXvFL5u4a7TtXJuc/fmjc8VbZC80mNdQjvwNiYlzp/HhB+noKr1h4+QbAC2GYp
rSmcQRc2KQF2gSgPe5TVzbvb+CIj6TCm9IxiJa8hpsEYXkNdnVFQgq62DEeBWGNoBjCGqCNHdPqr
OwUf9PSdD1cxbMw6Yz07TPxkeWROXgzxwmlR3+LneO/XLPtYbJdNJxbe7sVQogyrBEJ/CC0MTRI7
S0+mgd7h5uXa6zghuaZ4SMw97yx/Ve4vw2rSDOcH/W8o353TJkRe38EYyarQdJBtx1/s2WYG3N+k
jFi81H+C83VDTdN8gkR3pXuhub7+h0X8Hlogt8b9NRv1hmF3eWckm6GeD58yw2g1YQIZYoB8nIqw
T+HoAJenpKoWsC/iEte8DwAB7KIX/krj5MQ5Pc7361RGqFNTbaekcCiPPFeabFTtKkck06UdpQie
J/HO1r7vONS3Lxkpj/jDVCOKFiI/mnPwcHluHpgzOXDV5dyiWN+cqv6YvXuRavIycdsqh5Gwemn2
iozFEmgfpawD2xnu5AbkGG6JZfjPhLK1frA7AAN2fVQhAIjHqofgIwqBeKMkR+ODy/78mbwdCLXd
z5dSAqLYytcKcny91i/x9NryUrUcel6Yk3P84HzjS6dDeEvOYzDOgh3VpaYkLWbwc1CxJuHQpReM
CM9YCqBdrDYterKIjoubj2QDY26xcauNAmKTgZWQWzAXe5XLhZQOwm63ByRPW7AeLlRyrEaoq6aO
Q8ebjNQHrA1aPK86sLPT7Yfk9JjIQyiyG25CD1xi1ADJWLFdJ8iclkEjq6PLzZtKtbx0vLCMG8vy
FxWHdg2FsQ3oLXYW9f16UN76rOyFqpVGjCbZBIXQXFLXb+a2cXXkScSG6GKtMsEm2/liljN/sSID
Z92PIrE0++zrUKeMh0Nckez0SDg55Q2M/0k2Ajv/AqIBE+PQETwc0L2Un9B/ya1s11HF7lnON3Bx
gWuLJO68gMdf+wMvXSuCbRCONVvjBbMDB8goYhh/6s+l7+6ck1oOGjgtdoaeNoBhFgH9YoPBkZrh
MBveRmi/1rSvo4RsaaK8sT2OLRGstMGlWZ56shR0WyC1tSLTOanvgSvbCENNbKS279PEN21qpsTN
sL94cfDtQ3Q5dMTLJHI2d4DEP4BBdchKTmTy+tdDa1vdXCBhTB+/lfJQAsAd3OZFN1C2H6K6AsQB
OfPgqgieanKbvTYs7XyECTEhbUVfWBgfJUuSSUuUX22TB8TbHUlJejn+xSl3gfXAt6TJXkuDinFK
/LiKVsj+lHKlZVKNgPqSUazaeWG3uz/ZJ56b00Bih27rrPEOSF082opJN5M9yIzz2/A8WSA4w3CV
D4cz/78I/gEFdzmDj+kLNWNtMhXTWaK56JlkwVxOYJTssBtKOAou1lN4e+OglYf3GsvH29Z9V4Ce
N+W5JU4fGWl1i+RIIO8kypFDUjSzYkCCX6IvlRbnwrtMBBLmHIRtU1rH6P84qkoL58QshioPsbHX
XLfFmBFhLpX+v1IUQPVCpYyd/TOfDI4JeJyEuMBRxMu2iRA8nV8HQSwGFKDKdxxenyYO/xhhz/Y1
YIDz9MGigO/1xC8NVc7mkNXmWDg7TfqcMpT4miMP9lLQICIM9DYASjmkv4mUDsaSRhjqHUaoGXsZ
PKgDc6L3aNv8UCJAWVJkBOCmSgenGaZV6yyVrKHmNcZKoN+14BS24GlkAOc+/xFID879OYSRnXAI
Lz8lwAKHgsPD0AmVFR1lTSi6Ta2MHDRXy7iNvHAKqf8xlEayxh6jkEY3F/Ta6ALes+kkEwxtmXH1
bxlaXDFVHrWBPXelKboKIvA+dvIGIoaHtOcaT23VOPQvSjWcJ5RdSGGwBmg4DlDbXRnHziVHDlHq
PpXkkLPUUSGgi1iqc7QVQyC6Ovn3Rttzuy6rVIvYkRGD5jmDGxhrL7tjn1IaQ9Zflpd8lxfXchst
rv6LNBMgywiAgBwMV15zhEc+TkToVDa2dZwF7B4u7qj4VGy3dtwWaSkBd1sKgWZ8h0wSSQYwt0zJ
axlF4q05DKzaSsXclrI7v6Cg1msEUEdQxo7x0zx00nT55qEidjWhzthVrL8yxER5BTVh6wtLPi0J
aGizTD5VEFIKmlCnW/P8j3kUSZrNEpqWF5loiupuyu/PagQn7MxAWbio0NAsFAnfn1tlXaF5xdKw
3cqiltU21LDQB5glFD5eNQzSvI3/o1m1cOX3IvhwhN0gt0TM+cK+Ae8KN1QpYa5sMbPniDfQejw+
FBt31Q7D6CdxeVrWrtkeeGeFNhiuqgNqBuX2GKN9KJfImGqOmmYCfK4uOpoXs5+y97NLdTdDp/WV
CT5D6qOdU0mF/cfLPwEjVgc8atCDl84aZLRBq3AbsO2CAyM26bgJkOgV9H7v89pM3tBcVQlRSZZg
aK53ZImTb5LRIrOVizzzTMg/PWJHa/qx1dasrMnlCSP6UyBOsYIN7pILvkZGGgreyVOxVwTGts9I
u5r6bkQfKOmiX60nvhzkyolFuAmsc6+7Om/RqV81ulf+WMbVsmXy8aiCtU0bfZprHkUaIgzFD/dS
k4PylO4v41y2uSlrDiHr1ljl/Ek51+D04bmKwOVELKdAoqvzu4hQzj+wQQfnHyXG7c2hTnavRTht
Ju4IZaQH4/9EbhVIPRq8ZdsOjac++mFDgCx8Cuj7lXwGf1pHYFFcEkGTog2ZoErS7zH8PV7AvzvO
LbMVll8duyaL1uQylECV9eZIv/fi/MBREHj5FmhX1iUHx6L78AK6uxqDYYXzUYwkG1YYnfJA7jnx
M+Xn9ARtlDT1p4ASAYS1Anhyqued7nBw6z0Jadb3r4T4Xc8qXn3bwszP1I0daigCNM2/yY4FfF71
v29p/vKgdvFtk3PlrxB+GnfqNPwo655yas7mhuBNbk4abLhZFr9VpXE3HbviUBlilmAoaP0kSMUJ
0uWL6JfSO3Do/2mCo2Hytl0yDGV8zPFZ8ZaC6ZWZPFQA/TUbmtYbVEGFHHQw6XiT6qqAjNntfel7
pwsRY2melO40fJWRICEmDovxnvQ2IROgZbvcVRTjHXQYzdF7npVqMj87t9iqw6jhiQdbNsh3dm6o
AqlzobT4xqfzxQdBk2i7LtrDZtH3ZOcPcrAWYv6Bg+ot2yC47Z2iNCiwBj0s5Q3eHiQUxUmmB9AG
LZV6MHkBSJgIpYgEPnF1EX83C7Erc9/dzgUWIZb9GQmLPyIt/AUK5DG2avfVWBNxst1Vl80z3IH9
wB7SIZlkK3ws8Ev6nn/pbKZ108v3V5A7wcg1xbyG3vxcjLdQdjqGgaY47VduA/VFv5xBS/8xJtaj
4Ji7/UNPNzf1k9Y3QY2MDpKI6wgzHOqBoAB8kBF5a1AcNAPFh+0T25fuyqlL+NoqWtYq4ekFphO6
hEMRP16iA0M5K8MwzJe0tMKVF7o7saUyIlitCXRypZr6Im777rZfcZ7dUTde1IBV5+Tjh4CNWE0A
0KsTEhabIHsO4uuvdFe8zkQUO/pyUfYJAG9HWZsgThp0dbtNdgttZI78xIEblXmE4PBfchKT3/fZ
2AzwlV1aDz+ItYf/Z/tbtzMG98jjprqp/i1swtnc+N3n4m5sRw6G4BF/keWAUzb2E6CX8tM4W8M5
9Ai2fVksQmiBI8FPgctMD6GhgpF/8l1nCvN7/XOi0Cq1n+sGZceqqCmt1ihjcWwNDCJQPJJjY6xn
cT8UGNiQQb6v/p0/j0JOnjfyO3yYQzXcMUa6ZVtI01pl4RghSQcQQlM3s04oleEUl1T3jjOUf81s
env1Tx/VzePxMdnJWciSadXhHEBgNlcmOOGEyTtKf3hgV8dhC3Vydjg8UjAwsnt2jz9TZJBXgfjJ
NPsLE7U8jKG1yMQ2Y/n0kPrqC1LA7WdD6ysD9P0b3Fhv+k9ydhZy85V6azBCAMOJS2nb84y6wiAO
SLvdENgYmq91NwMEznm/7XRWdTJpao8Kc1knWflUcapMIoHmU++qaXDqfh9WBRsjINgkfA3gtjPr
YRyQG+p4R33ejOzvkKFTg1WRrK+FUfJU7AxPcxbTlADeMtEQjdYILIyZRxmO0czxZnpFCOIGe4u6
TLUBwJr2oQRTjM3/kLY08vhH2MhPls8sVjw4vj4SA+LGfB65UldwIwHQS9SeRZB+X0dJvylI1z0P
dGBrUDj8Mm1NmhWEpgD5WhTnm4ERxPddqD/7BKz5PjDSimZ3yJZtNbgEtjJELyl+fS4M+Hx/RMRw
W36kpGRNnMaNJfusBLzlSArV+tZjCRVZoJgTqmtHPfwCUpLF7HGZh96biyJbYawGwIZvGU2LvvOV
DQuNKQJk/ySdHdkpYwgJRxY3VaNOy0P933ZvSCNWvQTWesbLA7ZMXDRzZXSpFviJa80/QfJkCrJs
ZL3J3Mv5raIy4+d5it7p2v6+9XI31L6KJ8P7/pT1mHlS14BEJqPefYoG+H8TFTk7er5BIcGaqNQj
1NQvalzkdhh+HsB7AskXMdD4JhF4jxY38dUe+KOK1sYHScgxzO2KYAjUFmzJK8KVYCHtlRmuAYFA
3W+cy2aqFmBvex/FP7dssO4iY7MIc0koEKQePegwGU2IqX0hkbSghiSbeHjCfObB2kLYKlJLOsUX
UMnR/nMFzqbh1we6GyculbtdXgQyKS7+Dyb4u6G8kBoHTuYE1lj5wRYkFKjfTqyixqYCmKqGpgMc
3f3y17oGkFCmO1/fSPFNlXT6947w9MMcaznP//vIgTPJLcDZ3E+V/vGUYXMgDcv6wjDNeq3QU8ux
rSAHWTr1aLgPPgH2k1qmcuG49wkT8+bsymvjY9ObJsmHBIsciRUZVjIsleulu2cHHDgbEgzluxzC
83EoD6XDV2h6BMt5RGqpzIUa+oqILItTWv1r0JHVBFie+X78LxzGGwzdT7lErg4HAoN4QrKVlW9d
Y5eFMgeSPQxcDODm+6BLpeirnTnC9Nxw/VU7WADmfuCSX2x5G5gph6/MMuH1JJ9HPNvKN6ldT4gs
UyADh22y6GqnsUUXCgISqLb5HB7+HiNEK0a5b34/e5B+OZ6Ef0yL+UP540qIZ4z4YJKM6f8upSjd
VvBJCvPFEyfnxW4tWpf4riItkUvv2d62vOdsADg9SFFL4pq3ivIxhZnldEZ0GIzRQE0/wsHIf1mu
mM9yev6+iyojxLS8DTWWR660KJ0ToQZZyBtZF+fRLC8Psgn6kG8OMvbFD+Xyc5XsQkyW8rB/aAa4
GBQoNyWSwZKt0z8eHsTMfbu3i8BF/NsidRPoWXjuxZjkmsD/vIVvHcE6loJPmhjLtY3SFd8PCdD7
vOIiwKdAwLiD4mRyOyXaKeV1qaHQy2x4bTH92FgD1dALDqN+FAssBXd61dC0qJaagNsbpwTpwidb
OovMJiEzejiND0Ca/7/jBOiODe/1aeJS7MPoL+r4prujO9YV/eQ/kVXA2uE05+y9wTY/6MLHzi+m
m+PMlsOQFWr9JAIZvfgbKjjGOW7X0YJkSp95VwWsPRQza160uorNW5XaOSGDtWTq2SFbJX8icLgk
KUzwH3wZSHghaFZEw6UNY59pvBlzEkDZK8FbUgqzZnTT2hgwgvpMNvyQGO+AOHqC4mkfPZvk9VoE
HmZkFf8OvQRlJRynoXbwAL1wFoIAPnK2uSL1BZ+/INlG+FDtl9ZOP6tDO6Wra0C6nptzaI5DGric
WBfBsLLu8l0VJtAtLz+WJeww7241KWMAIrf0R1lEfZ7I7/AS5vPVy+QfInSpAwdO/RrHJM8eeks/
+A2yGN/dR+vG77T9NOIP8FWTroX4XPxXPU+5ywAnQeoYLVOK8WeeLJPXZn7oBQhSyr2YmiF/SX5V
syhkGDAuLbR0HXk+1yc2VLTdN2+jve/5lHbhQysxWAK8xc+tOV744m5SxQGP1LTNU7YG6Jb2dSS7
xaNR9Hv5GNc3kMIQUX+wq/H2Zo3b9M8YvYKPzERvl0la6lKrgOAIJEQFdaojm+cMsD7L+8WtzJZA
k5QEcck53ltFsMfiQ5IF0k6HRLbCWiVDO296iQC8zl1wfJ+/NRLyHBZ+MbYnCzhbPaVNOp8wWP7U
ONRAjSWWiREtj4BYSQtoCnMI+ut4ueLjomTc1hGq4M0MI4SJdB89OTnVA2Lc0aZluzflpFrVgZFL
Fj2di4KI10Uaf6qRIY/NjtBg0Fk/c5i2U9VwiCmlFXIK/S3smEhPVnuyVKiYFQa8xJKtkgxn5M+D
Hf8O9h9UrKIEj974eD+YhYB5lasblUuwScnp1fYTPVH7TiXjiJyBfLSpwxQczfmPuVdZpy0k2kgh
2ypZW96iPFyBayXIVgdq29AjQh6MD/YT3yEwQ6PjDPDK6qnVXo8xaqDPy/Jt5n8DklGSRnIPG31O
+R2mvha6lGYI4OknC1XBzep6isVJtEe4DNybDWK6gXw5DazWEF5OmCHiM+JQedsHYfnL7pCVsXaG
q1bRnuNhC87avL3pmXi4hhaWbA6w04ajyNNDOWVwD+rFMSyMHFKQvGnTqRSo1FJFsycOwf9hiNIM
JChPPJGh5gR6WwOG1puqCe5erlkdgwrafW79jX2zkOGwxJ3wQURtisELIVNYNsOSqLKZAxyr3eqS
jxCm3jIe1OnDpC35L00lp1Yqj01YMyxAhxTZZJFfNNc+UHddOIv3+nAtrxU6A6yM34e72p0t+nxw
+a3jUw4PB4bzJUP2LeGTiDIFAeaCNYO1UWi2bAIfBr/XTjFB/10SVgUEs1XbgJ/9Av9vnTvhdViU
RLF+o4KyuLu19anaNUuAcDqt5XdtcKJQ29DgEfvroViRrmbWjirifFzTfieA02XrzFdFwKfgq1i5
0Tbo1/zj1v+oc/bYJscmKdXcKpC38QfHGTVdha3WJo99tP0iR/I5NXEAbZ/NkAFOx6OTVOUlbNBb
Rozv23bzGP3AnX/LZjb42jj60RRjGEt31t8vpXKVvfYPepqtusX0RTCyr9Yz+uC9dSeH99d3qJ4U
TTgMPWJ9Te2EjiYmg3rGRFVoKUEEL6DBkEcoSicTaS22FTAtxIi2wRiVJsCx8nX3QuB3yyfACjUc
eKtROQq9ejJMC96zu0zhYnfat/oQTc2n79uBNkrJXq7WrvqiwMmmeSQV0FmdsbicIh0oEbxO2NaK
UFkStntLrBa7wToW6IDYw6SZhdieF2vDSbs1SHZKRHQrcsoNMPBt4ZFUYM90Q1k6jEPg0iUZG1Cn
ZgVyC5rtR2s+Z180y5U+hEKODmAF9vtEXx1wkCEwpZDgF6HAzG30Su7R1Jwz5FYJh6Tddi/R3jv4
2CCA6ry9BhKJQzSIOBIIz0wnTwGc0aTIflnvnYJL7M5vw6kbwxE5I4RJmYIHpcUjF0gaY+f4To21
QexS2zD+fO9dqiA95/tx5T4Cf0pL63347Oh1IE69ddxhgYMXovYwyAnRBXK2X1oj5hJJAe50ajrs
6KlLIwmWloscfdelosLmu8egoiBy4tQJ2G4fqyK2hxfXxIF6eCFdJW+W2H7KghBL9IjyUt1miXXf
Di/K3njX5X0A5XTRAV1BAidvP5DdsuCc/lsmbFAttOcAfBC5YKCBSDIFiJjFqnT5Tmuf8dChIvlw
KGh7Sxpn4UT1VJWDFYg0ZyU/uidjOPOB0y2YqkX7AzFo8ZWnjLCOASi73OBuS3sJtmyx60PrgoQF
JZo/zUwABUGSTDxhY/lB2c4FGNZ4K2bW+aL7ckPFijMxXFIAoqNt6BF5+AQ/9fqL9nhMJ8Vet57l
H3tMjOOXEHDs7NmcEQ3YbyVYNBkSiNK/iCepjZI+AZ5udUyGLPjug8+VF+9jF6GJD+mPggYx6AkC
++bFExiD+Ffe+SpziMjDhogKkUR6tj49pxKaUjXI5EH+wWZ+mS3uX9//qz4Ql7sen9LwKDx54a4c
SFPz/4wozI9iRBN6Zz55LnI+RciGmALS8BcszQVnxr5zxwpEq2xIoCJqKMnaIJ4PobLpaTRbuGtb
mMFVYIMapFxpl2oz0PnjdXVFj7528HF8R7bFxhve01azH6JVJUSq6VUXCiGEMl13cFd3Bm+TjXqs
iWqY4hj3N094Bxldg2PC3iBlBKYud8g34fHwR87zx1q5c+JXLQIfF/HKybaB3ox2zoHii3/Yr39g
tSPGryvQycDIHk/8jZu2dBfGAwKdHyAKM/FmyKo1IG/qGvH6OhXznclwIkpOhLzbQKonjF9IrzdU
8N+erpg/U/XTyXWuJnTn8Vpf0HbH4IjexVOHFCNK7GRiGt/CiXIlxs5HWM8/MY3aqhOotMlWIdjw
INiDDDxkZo4XNfgf6hOleDQq3SNIFgGkc1maeeevBUQ2VtDV+QjinrtfsGUKk9L00cJASUG0Tr1C
2ee2V7y3lN6JHqTz8YQpXnvQKqbDWzrmDRVV1fcN/9yv8YJhaEgsZYtMhh7UPVtTINKrpmJcvtOt
hcNSqcYbEZnd7xI8dKcF6lg6qXw1bqgAyeaKIXAIvDkmK4zZ3jttCBVIGDF42j2M+7HCEJ+J443r
UerKIV4My/xY1O58+4re8kv+e6y58Max2VZPzoziSsS0HE3aX43gdaholH+MwzUGbu9UwRv9YtQB
s4OS5l0IuQh2fWHwHUSQFF3p8YoIkGV8TZ9ZbApejnU722a9A9m2dJFBAljqp5CuizcNd1txFcWW
1mmgyo8bpznqith6cK+zRwjERVm2D5FS9JvcOCcZV1ocTnENuCG7Ef9bC/KZItiGUok4IoYhgVOF
yolgRfDb8M9F7xQUWfGq+zaXb73ugagpcVHgmMZB3lhJNdC5iHgud16vdtfBxzgoZImbwL0a1PJu
DnMFCxPZeT5K/uGbtGZ0lsCYG9dyip20pf91X9K/Kz0txBFa3GRi75/LXv8tueR10hcq7JjK6tvr
XVIk4LoUvHWdqbLdQ7yMAYApTxLjB17TTaRDiZIuLrwdUyxlsC+scZginHfIX397W2+6QjttfFUy
2x7MENLUaDgreLqavFgmpL0B2Jnb4zQQ+QhCIREElGYj4z46PbrMohEaEUm3EKVs6mVVFyOhg4Ck
hk3n9jLkOjbWpoLA1jyWDNIUpJmYRZZn2JjtXgpztumakSmHEaQmuqS1bwaG1Q+R1zi5yCya8YA2
BFkZ8BCSlGlegfqU1bSFWVPDYCjtJ258gQQh+z/3lzjHY7uxAwYy0rW47QWGIG3wAiIBddlZf0pF
CPfq1NoGgxxbtWPMn1J3vrqaDFVl+MXzLgts2WTMmRX7xJQpbLD467JwKa2ml2rH37Hq3SH4+h0b
eeBrwY4HIpduvycVCSBGY51BP+w7nw+rR8gyQ4HeTipjEouQVTr6VyVBrBMQtYVYHGCs42h5RjQO
NdwSZ37CuRTGKxJjPWplrshQKcpFRhym0PeKvhCxIjGazJNL4rT8Q+KgiaeNQFVFNBzzbVvE3lhL
T36XXNUESeUhyGiMFvfc+KP9wIupy0LyjCJngNK3/Itjsl9zuqWk6UE+/15zN8mRr1V5Amz/XY9V
u5WhjJ98l8Zgm1s33K8nxRdImaWFGWhaLeK3R19iG1JWUy/VDl8PdpiK1LQG5Yb0oNoqASrUNHnv
j1in+XReGsgDkyWTPsSGM8NCBDb9z2qe0FahEleAFMQuX2S38uT+vbQ4q71lLkf6vHv2hq0lYkyr
97LNsqP9bf8oDAijipd+eFH9/ag7DAWlFPtOKfEI2PQB4FNXD7HZjjooKrLAHgWhSM18YMU3pk0z
jS4SklLXoRJgSty8ZVsYXoIBRiwpoQuFIydO14XlJjI9NwA5sL+sAA4CnKWllDjAEQRGcGGaaIpb
Q3I5sT0TJPfUK1r70VFFVxntnVB1LDiX3iJ2Mi6im6+CkDyb9v3mwak6xyUaBEEz+49e3nMvN1/h
wZN//enzPw0J5pqrCv2meoboOzhmcOESInmV8zPDzayhwZ9MAYhh8QDbBbyBRGpkdRbB7OvDSS4L
p85HgC0OIglJ1ZQwqrbE2KpVXnZKn4SU7AlXUxEqX7l+qF7Ej3Tt3s3nk4uGx+h8NeHBwZu6S0Uh
COW8Ialn9DvIrcjZv4KvXnAd+i+QwDd7kcVOMZgKJCQ0IGyVoeFJxmpsODIPizOw7dyf3ELh/1Rz
yXxszO4zyB92kUj1DL93UT227kUMGiHwJKyFAgejozBz/DrxMqv+9+2WSJst95Yt2KI1YQEGRZVc
9TWpJLLHwJLufrPclyaSsnI5UbsXLNhSaTMbacandyLY03aVszsdXY6mPZN2pQYBgktIt/Wvec2A
XUggHOEJxslRbvwFDMNoNN10un0zUedxqGg7e2JYEqA83tx03tiVtpg1fN/zG//w/zgCNwTB+nZr
V1/OBrpYTF8vY9hEKwhSv8RbVlCPYjciQuvITtj62SuOiiRPBEslPOMuE4P4xciLOD2qcWDoMwvC
7PGyaVPbq2VHdY9tEBQfg4Z+6LMy4LvICso2Jzgt0QUlv3/HVGtiFaLSNjej6YUrUcEwqE2NcRGX
wz1UM8neeFtTmesKe61VwSjWjtxJ8jVoj5jaR1Ch2pimNIR6gasqX0FSgsi1JWJbQwucdRzyt390
ZwTwYbipTb87mySFdsiSPL0FB19r12mlDyVvLhks4hla5syeyWibrrVhzPQ/2QQV9LVz+qBP+Uj+
p8mIOqb4o6adKri1mpMs4UJ/cb+uvhEBuRWo90MLYa7d+X7Qs1Gsrwu0UUKRAF4Gaf5EX38hvatB
kPHfxrZBvDCwIRh4EplAlR/km0tT2zSzbcMuXPMDUN0WYijcMAN040EhG1syY3LxXsgSIwb1iaGQ
qYKanFs9NosZOR6XPlMoIgsVqQmITPhE9wm8OlRAK75YDg6WfbB47azoR+26lOibKIdrbwaxVtIr
skC/CIThGz3be0auiXq7zT+nTbT+97YziRpUn56o3RU1w7EXzPBOpNyAsdQgoyZ9mKpWKH0R32Hn
GwFIIfiALCnL15UREYxXlmccH/NsBRua6eaXxYUf8W4sHNbnEhan4XrwW1qlfxjJMsarPqgvw+Fa
7YSoMF/Amy6r9zaXbRGBEK+g2f5ymtiial34Xxz+MxyIj229/jCrAoJPd9vrl8f9F8A/b889xUVa
fG9CJzijskhoKGCGc9RavLc7ijjhiQkukv87E1v6YhwOEvL6f7k0ZXYzhxtQ1boGeqVVDz/pOwa8
hblJzuX2LHq4vQpc0/6EkmQr4SvFWr8niEEFoT7vcsn7sXeTe9UJs7MW2dGgoCv9goBIZqR4E25q
Ph9Nar074ZApjH7nncnnQvgN41ifgTmNOMSey2rsuJ3oQxnFcUFxVDGHI2lToY5t46G8chP0V5uj
easgNB3oJvj31xnFzK70IpJD2aiv7bI0WaeWNzJhUSDCdXLc8xiwSPgElJ+qMiZ6tSp7Hy+SMvYH
S/l4gCLd0papnnZsfhZ/TsTJAI38u72rSyN45BpdIlvccs/nOZKjRUXtu9oqn4jRgRHdn9wB1hfr
tEJmUd6BGzvk7j+kn6u8h99j1I5Zqg361lWjxCo/EaSHoWpc8dCSG7dISiqvkDYPVq0R6h6n3pLW
18KLNnSOnC/BSFbuqRx4zQmd2pLWCZqIzhVEhfb0CK2BD5eWX8LmIyY9QmMjd9jtFNdCZUYUlS/Q
S99hVaGXY8t+2ZUXWKAu3nDDb5IG3d26Po/qtdu4YS6FkfUgxumw9XAlAK0wEc2pEMlQAu9/Ahpt
S7SvRHoUUd/8RwUmqx2y3YPSlaQpW/nf0MA+u5g0JTZcFAWHaRggcqaidvlzGWcvBtmhpr0ieKRA
GZgfhYnRExrHExDn80fb3n12qJybyp3OQDJSSaWaPj/1tqj2J3Dh+hti9D7NaDmRvtClVlUn6ib/
4xhz1zKhvB8benGxHQWmI+2mEnM/vea4dG1ZguBP7Ub5P7ASx/Hw0pUk8Wb8I1VALophM7OIgLR2
BUDUIU5l+fnEzJxGbC33KkKsxcelNgxvqhXq/BW1VToBBA6jG54xu8XmmUeS8wCO7nvEmJjSjY8t
QYPxD+xq0VyZ8mOi4hZ83mshQrchRqnmm1+PplQLJ0BbrQ0G66ISgGeoMPrk5u0+JWz9JH7xBfiO
XeYjO/7F/DmPPhcfFA+cdUWi2++VHPBog6Eix1B5V4/WCcbVyVElwR0h8inhQNOVHobCa+NAhyW2
jTpFkoo1X53cmhMaZ3cTEdIQHiyPSUtaSiI0Gpr8NueCON/YPxUzaaXIbiZAaspo0QU0cHnf/aaC
Qhmq8RFJ8jRygyXOpBMFouJGWJAWc1sGUm4ZZXO7EvfYWIdN1FoBn2juB5ci8vwxklVbFZGWFgYq
ZFQqA9OJ0nEnx+azc8k3AzbJyjMpmarSRHtJiiBwYT9vftnohMA+ld0bgofa9Nruq/8F4D0ZMyeZ
ogwmZulmIuyD7vvhoFumIBtyc83y17N1E99Ciypra73/LY1n/xvJNvILDlY98x7VMvTzs012QC0p
0RCfn4oRfQHq+SC2aN3TrfQUdS5M+gBPHx8C25ylYiz0TxIACPmrA1WH7r0OLAwO4il7vifKaKTo
rcHtMNFZ3SE4ptoYCsq2638fZLOrEo2CJ/4daeNX33oi/W6pLj7B2X8jLuAkALDdNoqI4z/NqIJ0
XwiC1/To97U57Y3WBQHg8ywxJT1flB4etEgixcolAGI/mUO0dcqOHKK5McZUMSVLXrTP3hPEdtuM
RYeUF8GQq/u8tRjLZz2c8OcEC8EIc0lPOmWnYNck56VUT4RyTrLZQ8/tv3+npGsnB3oP3j4/YcuF
QoI6QosDXmgVqjNZZ9EuILlHi6XaicVmXjeAbnBer52SHbPFdf/82D/RBh9l2RByp9baX8e22eoZ
H+NpTMJR1oh89/CIlKauU8xtkCIaohg5SY6YbNqIyiG38V7+e3waVT0ZxyBfKrKTVhcWVtZZUCTB
CEyFCkrcciG5AiWgQsw5QE0NL/HbQsQcBEJL7ntT1ogkuP1kfqTPvtB0ZnfLMrCtQAwcBWuAqVkn
KETdNkZe9mfSbs1lUn+4hGV7LsMxzh6+sm3N4vqdBvnC5JLsg0Lwqj2FaArTD7B6rPfD5e39Dycm
Ndk2xtp8jAi1cR6lhH657Zn2lpT56GIwMrJT5pYmLbdBMK+T2/ILrN0Tu6meKVJu2GH5610sISZF
MiSBHASSUEEH1jw9ca+UBkBG3daWRI++f6Tbjntj/rPihXib/WuSjO2AVkwA7IrQaui848D2NHoc
ivooscu08Tawpz0PNkrAyP86TIUJKZ6E6zMuZQYuYbUsR5f0UM135iyHQLL+FFOQ0HmkdnthED+X
2P7Wzvdxo/hGZAHp/CWe5dBvf579QbZ94caFlL0NkLbjB1vpBSm1OYKm0CFKrxXNKSEe2KEtmvaR
7qXVkI8uJStk5AYnYmT48VDsr5cIxu5lTbqrCY17TxvAFib/l3e9ZgSMmp4VMBlBvvZr+X2IewYn
C/Ot7YdabUq4TwNQhEaKUOQWD1vFXyfzW3n4JahhUC0MG/VSbSvm4LiCEbSXTUYW1I9IugPDgc9O
248Q9S3EXkx2wFJhRPTruRlRRxHPjPkogTY6CjaaWw536xJSdBCkDjWMUNecW+VbPQYXjxVctncF
ZBvmfPxXLb0lCd4SfvY+Wojol+YmUs1fvHZZlupYw0Cmw4L4QNTh0TWRcLLOMpzN4mR76mhaQrUv
RcqchJsm59e4yYJ2V8AFb6q04mWgG/YnHovYRKO9GEeXqyLCTyYtm6drI1bt+HGyO6+Hf/Qqt4Cx
3i75hVEX6m55ObTxln655svEjpajuT8BuQUe/R2xdnbCf15Avuk+AN9r4z+Zinw5pPxSGKI32uHV
LVHpYneVr45hCybq+ypR58BUu7dpNYUJKh9o8Zox4VtT1lVYO0BJyxYzVU69w9MTr6EDNrZCksWR
RdA1OjAm4yk0cvRiUHKz1GRkE0DGoA8GUJwkqkUvKuT3qsxSCAXVhBtZznQmQYSLlkWdOSv9+l+7
AMbhsznMEwX5qOOzLFF4d0xb9TjZUvvrPxFlQvyHwqxG4I7Vjm0raRiMQ6i0aGuRrB2MqASdVcyk
OFUAB7jzgQfkKYTKPcmVUeAP2ZLDIYWmNJTYR1UrnOGbJt+McQBMEcZqUtYn0IAxO0y50yvv9Co7
C+S9zN4HNd0Kam64iv32gjeWZEmcp2plNGz31DpSuYZeLdWf9V6i1iikVss7QHWigPZfpaR11nlS
lnxJMv+fmMaXZEoUs3XGQKQKSOevok+DClrgVS2I0RhroO26iyvelL5FizM4tPRK1QU+YRT0losH
n39El9eD5Ni+qCGr/7BB3SLB8y+qa0tJSlUOGnQY2+nr4gDYhPma+xus/fEzE8/MWsIhDrr3w3Wm
Yvr2318FwrgWBw4Cb1Zb6R/BeViirszatG5M1cc/oydqTUH2uE4T+xbmhyW9yO5aRuUclzOwPhut
znWr3nrdJycbneRSMY/A29WE/lzibr/xx5HBe2tUqdCmcrmgptWfy5jAHOEvr2/VXEKVIxLCvYYa
axgPu29RMi6/Y4v/BFt5mIZmRoBeiY/ZIZTbakRDbkT7Q10HGHa7xymEBsehUDREIwujRkWqgFBZ
fqJ9xMDus9fC0nDDF2K9pb2JBi6WQo7x5zeruhHiYvSKUEnCzgKd8UPTLODPCAB6prRngvzbGLCC
hE2z97+7Ed4q8TBoTRnpDYJpw11zgIrO1XK2Oc/aghAniXD+wxJbACtuJ/hcc89B1XIPAu8PqA9A
aAf2iuRqYzuEcSzJ67Lq9BaVG2lEZiL9Bp/GxgWJNpA4fMWm0cOKQIi3BVH/DZnITpb1cadysLad
JG/uHpR+zfXKcOhz+EYx5sWu1ADNsmUmSCE2H0Xe0Wfqmo5BeZU2Z6m2gQlE7EPNvuFCowHqLXrj
CCBD7XAxuvtBEo5B5h5pPE4VROEPUmd5J6Lso8puJ6eEXgDgaMJQvpkf1U64MkJpCFz5fopdNXgx
H1W1i3jcq7sk72tKrhZpX6/p6ZwyypGp33ByRIYUupxPIQ/r/tTZkugsOjw5ywXMAfxICm0EThfa
bxCztDohVEYiHly0g4VcYGR3iIxmUdx5qrlv20U9i7gMNGGx7FpJ2K5UgnmU/6FUANwyqaSo4sCU
o1ex+gN65cpymukoz6Nx/fdBY4kGpF22+CvlcR8PLNjnzSC2YqutNV4Javxq4DtYXXKdbxk95B68
XMUoKfsKgf7oQR6yp88sIntrajPdFF1Z5zcr859ibyBHM3r+jeTz31nWh1OsROC47lhYg+gpq8H7
zxTxC652eVMwaY7H/TKREG49AC3K1rqKHJAY+2QI74s+lPhvZni5r45wWYUxAV4obi85NnCxt9ma
oeqxyhf4GBz3lgRJQXLT+TFpBmt5O4823Yq90yLaPrJrRQIZHBrcML52giE6EDKrwjAnWJa/EiVI
voyto2OFn47ePAraNQOrH3ObhIvejxlQ+Aenbe/nE696EFGPFoIntv2p22Vm2F6W8GVw4ylmX1Yr
gV7eIcw5kX3HhFYp+4Z8BO4DFBqHyrWIsPrL6wDjyq/AwwCca4SlZJadN+QgA16P3Sfx6rEKTISy
PixQAlM2sIU7rGPn38GQjDhUW2ELEAozxm9h1rxYnbI9TuLk1K0ps7BhWi4ZTRzNTeVR3fkh/4kI
S5OU4OJjLiKEoee765gwCFQvN2DMczoss/WENDMYEJVOjwqAuhf0vA6VXOq+nM+B7F9mbwCWCyJR
mrtnP8X/VwKqK3Xaxyq7pWEmMVWpiy0G9KPtU2oHh44HywZvsz45SUxo3JoJctIjnx742CRyHO/p
zjAf/d5qDB6lFPSv8Nr/FpABpn0yrwjsJrExAp4bMJktoD0vhe1pSV9pc3q+2BGe+2D5cIKE7nzF
UBQD280vRm5Q1STQSBE7+HVHnD8YFW6yT4aO4/0Y4SmesnZfLPPI8/h+QHeN6ZkBVvpHiIz/aE5D
0IXJvKQmyKKm128sI7fso0BXbz5h8lKKmEGw5tgRPilKlmMl4581aWfIWsq+MUfFzgn3HwJG3wO8
DfsFrCWHqpEjMn5f/NFwfFOn1PUUQYPAqQF0FVPyfuTmXdj2ELK/CMpz+bqv3RsIWHD6y7YfhdCI
ZnUEjyPxYp/GmD9Z/EFzr9JV/9j8xj7acmEBK+WSLp+2uGrD9kVVMJ3jFYF4QFuj5ui5Slk4RKUv
/yL3zcUzCemgH2YxQkfDhfDplq2V2mOWVoXz7PG74AGXoSdjofdCtvcQfn11Tj7U98Aq+v+DGOJp
FA2FnS1FJ5R53rCOY6KlFBUvCwwrZ1GtiJr2o+8SR+NZ6rglg4pqYlhgbRvU76UHDwvK92gAKihB
1R9stuw2/nz9K9Nakfx4A22LQgcRVTTeqhdG+Mo7cCYKw58f6oZ625MbZ4YbQdnZao2mtVnkJBpu
m8K2YiKfxR0iTmxUdW6305aQmm86A44etS6XenpAijCXlWZMUsmmGQbKwEO3nRjCkRSuLt7jGXd4
/oKiQXk0LklZa9FvqwvuSbxb7waVj/cY8abnstOgVVtlVBj0cxxYsIGmtL6yQ1R2Xok2rRVdiu7j
tiyosnqYhmS3rQZ23Y6PTff9HXvSfZh+rWRXY1xzInf9ff826g6TETAELLPywUOGORga8Ebqf2Z9
cFnL9As8absWd9o5rgHtegyDdr/Ylok1wJpUcPDnpmW9yDWqmAcL6q6sk/6Ilsiz/S+KcWj5f7B5
U4XVkICTIaYmtdNxDv8Leg2PKsgOY60jXwHJzuaD2IUERYm5eDLBeWPdUAbddSdOYykA1wRXt11E
eEpxZ7zys/zTc1suyPI0JSZllJulxhbDiYzESfn9q91o90h7Ur208DeXOdPO3EvHAtLBnofnOk6u
/w5kZotp0LnLaEGPc/oqRriP2J5iTp8UmyxiwfFoNjxpzWKdG8yWk6a8sT+oR2YG1TYPbTG0xlJp
nk2IAh7XThqC13nTE7JScvozv2EUoULuj4S5Gm7XpsLnekHSHiLY+tXwoSgmZlC3LmLD8cTHTxdS
1ruOGhVSKeez9HJRgK8kPdqdsV9y8Du6CBritG9wDWXLHo/Ki+Z8Tl6P//CQqwbeQYYoi+z2TJWv
SIbTXMbdZcw/MAdV/WIuBftEpAhnHQMP1oCOyg3HNKdV0kKw7Biyw1MYbLZMkwUu3U2nq5rYWLpt
HsaLqa9w8VZEVQvmefoZsM4h3zR0C+Qp4unYuhmxWv2ECHwbfmE13nw9p0lmncFVk2Uy5j/m8l79
c3hT8Ei6FIxyaFHdkqfimZYnxTAiLeaubMErX3KbIWFNkkycU+S7eUHrSDtEhyXKImVgnCVxqjwU
rny1Zg98RlX+2SOH4l5Fa2z9T2F8te5y4wsds9B7gDs5/MIRFPWtspkm5jUBSZvPsTCLeMnmp5Wk
8x0bQv9z4cTJcjZgdGCg+WDSXTzcial1lWMucHfMBVHiWpCSE0PKTnCldIiIUm+MuSRkDVNxM1zP
ifbu9ULMRzCjREqc1DeImCuCWyUzo1SmVXX2QV2me8qwHTkFTX+XGaTDbrjuxWIs2lxDbhhxvBIJ
Yo1/fb7wwfGflgzIPOLXg1G8aLdN6yafEcgOhVIpYpkVD/mh3So0ffAf663HR05UkULj0LUL5dFC
Rk7eWpGE8o24enrRSyLaLixfphZpuHUVPvfYZUamHhaAr6Ywi9boN27Fs3I/aKn0UNILZi+RRlYt
dqvZyDsGpr2lf9Yo6O6s5CeaUby3MgYyhL50p+JYb8PcprnGNt7CnhTho2c5D/0HrSsK5b1Oqu+k
TKdY7S5rqBR0WfNI18pUFfnXXrOzx2Rj7RkARQpr+9NRzRdtOgRC9SEAd/gHmLDBqaETSWjOp8dH
6Lj1pDHviWS5YSRkiY0iP4VU1l3LaRMtMdE9Lp8JUE9FHaHHeg5E9ryh0j3oCB3XHSnK6RBndOAw
5SHD0EMCWo0FZdLRTxqcRY0a8EU9X95zpoXY8g3xgSJeZppt79WlpMhs0gMqhcvSOAM5kGR7yK+c
IAggiOigzleA6jklDDk2IMi4NH9he1i5TsY4CQmmeNdNOCKl0YfiV2a/CPnkjIKy2lmgBNcv1GUB
ejqvTckg8/YJysJ/36kqeoM4mKUBz1zGTNqARcHXEx5HMHBjLa1ly+Y9cev9azqDDYGuXFloopD+
c1eeS1/cz7uW/+1khbA1UT4lU4RdBAdafZyHeuMmAMaHvG171eh6rGxDe1vUDhiLF1t6LmqJQGJJ
hVTvznLZn1bDNVOM/4800F/R3M3y0eqvd349nVjzwPDl6Y9g/VKHud6IuaOSUVfF3wU9bVyaknl8
atfTqwti859epvbM7WEBiWKKyXJCrAadBrmmDZa0z+LoV67IAl/egXVDDq25IFqfmx4xZ/XPQ6H/
hZ2YtUAGIxSFo5EXK4CvpF89VuPKVUCJVWbgZypxPrsnfOqpEua/Sm+rwU4k7vRbspoGkxKomL0p
mHY7XSucFHqllrJZtzjjirkesYwBZWbnjsS9F77q5JmxUXvdGyW36bVCeYGBzA/W/3gOlLGvT+7o
JbRlI91kbrzfY3cUhN29HZ/+4erOIjqdy32wcHBegM9Vo0W9ZG9Tzv1AZG8OU280kqC0Pt4zmi6J
Yb+039ZUIVQBFE3zsV6KjJYSDSc/eWxpfyyzzz84r5K1D1HPVHky7ya46M3ZXKlyNKTc1hlvV/ls
vxxn9xG82Y/CnyMDu1k4ObrRIsUvSgMY2tVwzscvi5D7IZO7hKqd4aHAHdxcjc3Rir00uV2mNrVz
v3GE2PB3jCBVWrlC29iACXsQSvg3ayOU41ZTgje6YTdh4VnQkUeQq9ozvJ40YnAHkP9s6mlgDE/D
FY7VLFqMfKK/jYTPcY9TqE4XOP7v+x6l8uZdNb5ya77iXou+GdEkbld5onOznKHmmPrxR7nXQ1ZN
hNQV18dn3BD2mRKRMBhYXALq+LhT6seVFEYvOG9udDaTLYkp+6j2f6xdCgAVJcfRwdkcPESk6/PQ
2zysv+PiRAntEMbUUPISqEI81yCYwjkNJRHZTmpBT1XQc4T4SzAWbD8xxsLkep0o5IW+R1s+/fqJ
1pUEmPTOAJ8guY42cgXqN/cEjiIlz8Gy0xW5GL6YoWxyXyhpqBlj2YJx6sjSdpRmcVuk3sDN9CxA
5tXkpiat8UMFtKvyGcd5xui/NWdqxVPXwRRhKVJmiVKFwumy1+ixIofnxAUX5jwLKIFw+3iL4WB/
i6qa7XeF2hgtMTeuBQBNYr8JtJBLQEgCvpSKBz7I9ZvUNTKLPKORohyuHFactvaaFfqeTavPNIch
u6UnQ/JE4SUMDeSDMHbtb14ngL3Fk3di1JMCOMUj+wxFW5iMNNLV1MFhSdIQBFG0e8kionYyKq6a
EaTEsGJBQmV5E6+JFOvzs8CMfLiTrQ0aeyIaH0aw9ENuN2lbdXpq+dSIPsmBQMoLYXu5xGffpOKe
WHotMjIH7EaGvIXm7aQ1dAah3Wt1W8w/YXum3G5bjEr+N6qwfHL4YnXREw/CvTwi8g4XAs2N1MIr
pstUOu5CwpSFZwDAZjMbbxnHVHgLxs+G7iQjx8BNV9rWIh7hcqHvEtAMv2p/Xy2dcFVn8jyOz9kU
8x3ChArlaAfCC2R8x1dActFqrda6N7jm7SKaZbJn1x7XvJ6SwstfYCf+7rOH2Xh7Z4YRzublt1q0
uC1dDejogusIn5VSaLROn6gsvWGNrYyKQa9IEeXYG5beR6crklmm1xCBPq5W+2OPEsF8SKY48AVl
607pSuXjRwoNbGpYb7FqFIeJit4KNnt07Lqlo7xsmaokyYOjgVYQffFaabwua0raR48XSlgrNCZ8
pVRlxzsmGWwEPC2A6+pxemBDeeGbhwkcY/hNNWGd82zmbKIK2NRqxJejTV4YSMWgf5ZL42JiE66U
152URNJGo0FbAP2uPFmiqe7/g2OKKR4BXJr/mtaeiD0eIN7pio6pT2cSYIr3ffJXzfSO4o0UANHj
PBMJqChbkiDHH7rnTDqCrVPweGJUjb2QqjfmImEgHe2UDQuGms05bsDW0ovLb1+XNpgohnPwSMT5
o+sHHKZCior5GqMasWkOgwlmTh46GZ+UhrysKs1zRoqHnmblhWd5StIJ1mjM+uzWAxrD+0zNehZL
D6+J1l3KXrstCNiXy6CNdolWKiarUz6reh0mUFpTlKfvMtLvx3Rc62XlRkkuWFKxDasS4KUrZXKM
sLCjzbZCVaCBGSx5ChZUIgirCcLk2PKXsuEin0qSrekIgW9ntszMWYj4IKDETDVTkio+sdaUcDun
0tpAn8GhOuNz0kznApN2VQuF7Zn+cZhsJnBVHuvRT97hDx19Jro25C3X6AR84x4qQc3uWdtoUVcR
l0wlo0hjcaUmQ5XsEbRNEQ/0BHDgUN8ftd3Q3GjCOWWSxtgUzO9wHYBiEcPdTpiq/LdZ/dGIvakW
+sc9ipU6KbUfsNNuLbEaDgOdjFyEnym7K2xaatPzMbPXnAq2HWDq6u2/hfYGie1uW7TLcqcVJRSN
Go+4m2YHaTh2ZUwL8/qZsAynEKl49KKirup8ykfY70okYvJ9irGblz6Kcaqr4wnTQhtmUP+5clLR
+LVJrIW4aJ9W/KNHjyzXFn+twC/aY3FBWlBkWFdk0JYWWISBrWSnijXgofFhRsXBTm9tbrdtBag9
S3ugRfLnyDNDUuNKtNbhc37u0xa0ERSpEr4I+5JHVv60NZJC+IkP0QnrMkHbBJt6Vtu56w3yLDeT
oxJO/6v/s0xrrUxapZwyVvg++h+JvkTMQOUC0ThiYSwIPwYCAd0Rpvmx1ZcaU9LDWnOVl3g9zxcj
BZobmcggd45SxXYIAqUg/zyiCnc8dGKscii6IluUkXbfK5CJ2juKAdW9IhgfS58sGNH7qULQ2cdH
fQ/9pQGJynjt0/Q3iwVR3ED40TYKYDp2o+/6viPDUQjZ13QedieQXXht9v8+vc7Jzth/gThwoIni
nET5jyvoIbENNymejE9D5rO8c/Lb8eLiiQi2IDF3lroPL6Ap3eAWq3j//VqwxpbSp/XzxSm/bLOl
NriqDv84u2U9PuQYEsdOapd9A9T8BbV0PKkKTkfHNlz+mxD3YKE8mBcb9rmnmBgmPbtO6gUD2MU4
XvYXCaDycgDxclcndoco6gadU0MD2Ql5gzdTAQIPlbuPuRVzbzn1wORiLmX6laFOYgcGTMxLA+KR
Z1AhkIVskrPxl6IgZjCsLdTVx+xYkFR75IpkRKwKL3dkBy9t4mNbaPrFCECs0tTh4P6umth4d/Sw
/VZQfQmPocsqVHN92dt9BgU2pdGoL3p161dYVtG43hRvfECIiLoMc3OAIS7p7nrNNAnCOxIem+Nk
z34zajj3efPGysRx2QATQ57YF4qfypdoIiDCbTvM7rIbPwXpujGSV3zg2vcICiHU4qLTph6P0wsj
hTZnUG4KrVtVUar05W0pLDpnpWgENTxqN7RVk3AKLEMaMxcJ+zurP2y4P+VYc99u4myRYxvhQy/Y
euif+zEDKFxZG2lK1x7kd1+K3nHlpvSLFheCbZxbH79lCalNkVnDyj7O/Kd2OhYwrpz3G+nr+QF+
TSMIiClY5hp3g8UMJal/hPQsj/t/NyE9vjjW+XJEVl5JCcTL4fDNT+A9qOG/6Bg05vcgYK5W7Vgf
SjBMiTddEIqAAwl1fMkCjI+VNUAD6Tei8Q6Ay4vC1f8Kqd5l3tqhm6pHwxpnYidbXtNOkSwsW0SY
KyfwiDLzAKvkWynmbbRXaczcMuqumBKsUXu83utsL9uxgklkKINnaXtXtj9Xl+2/gpwtPrXHmtD0
hYTKsfk/Ao6PWHNaA7EYADRXIqgc0GdcX3dr8o7cukl5HOO3YSfXnFmNgZMde6jUoBKs0N+NKAYK
3fvVddz5jMQFJpZKYZiTmtoGNrJlGUpW8DBn+GtEeBCNlfP172ZSsL/KcWNR4tTHYpfE/QrocKnD
SWJmZuE+SqIG0c8LznsmALUan11V5a3m+yOBx9MU51hpwTX6O74B+vje7obEowSBjo3iFk8M9iHg
QfFjWszVeVaRsc0Tfaajm1lJDIm3xWerYjODo5K/t/+iSHEk2NOMi7YPNgJD/9ywNgR7N+Bl0H86
WifH5Xdn2pGO9/83JP01Woy1Mrg3tPEhbLmPbi4Nd/Q4aNNJoaDbZOPi5k3JQfAKppnVNKTkK/XP
stHxj6gRxIcWWJJ3PhiCFiTNwAK7WTObrTF2MVAmAZ06RQloR4X31m8PLng93JHGPNKiaq0CxL+Q
xr+AJV2OFlmD8tSjQLdhBndQ/1N0ZUAEqWhV9OB8lUsIaxS6aDoxfkBkwkBg3nOa1NWkAOWsDnT/
613BpJz1KmEqphgp5W5nN0HXkOqxzy+EFYZnAwrP0yjTaQ9d1YKQA/7ixsyGTOzJABqf6/FfelZY
WTDsgQ5WyYnWLnJVki23o8iSXaLVbbjwg57qjq53HxfD1or06hOZPKOvEy0zJ/pIyIhK2bKW0koA
lmK5SoHxHPZIoeX/fSJeIxFX8u6KKYSTsTH8tveWvlOqOlSyYAbjwrdNpvrEE6r06AefWlVL6jzl
HBRKUrsAH7JTcN9ixKc7UQt80M5cLyfRucRfcGI8+rnH7TI3oQWkK1S+ETa6ZZZH642cvAh4td8w
6fZtq/DYCJq7/0fvdBqb53EsrQFF5zRCOh+45SNhRZPOh43cQx58r5fPCNDm1YlQ9QmzHOLYvKYU
brgMJbqDZu6IfXNy+Z0BP3tApacm4Qs8gYak4I9HS3KrVOIxv4f+HaRFwEuWwMIoboDgQVgxuLpH
KrSaikuhhEDid/Q+Bh/hG9nHYXmcOJask9YJs5cKV6H5bDRV6dhSa32dY9+8Az0VNIonhPB3NX2J
n6cOACELZqC48hKiWTdVDSGYFd6I1uetJv8eoTvjM31vsNyQOKZbx+x9PJT7ItOmlFBXI3YGJTOd
DvTsh6d5iAV3l750vIa7wjqQcozHtyUQ1V3bKjn3x3o3R+hCj+h5XAiJFk9caH7gC+q9dYybWPOZ
sH84hc2emonLYkgNaZSIgSYVfIy7T2HAg0VcEkHqmRMpN5ZuluhIHuM45H4f/EUwbXaAJEbExoPY
RYxQYL2TiPekOQbIhspMaXE6Un0uU2EpAorztkLfp0wqDpLn/7WpHRbNuo+x9JOCgJKQSmP/v/iC
js4Wzsy9wVk3b/CUlyq7KyA+cFcJWjWkO5SHHokxX0kpju38vjr5egcCLZjefTAfI1XU4Oev4cYP
uorYuoh+bqUPutDkihTc4WlcU67wxeYaR6dg48hdWsLQzHG29ZBmFG0XK8sR7x6j8/c3Cli/RZKT
aJ3JqE6CkDNcz76r950fCIvNvXvuxWPBezhkBPIk3K3fCsuHwB+2+AmxLu3Fs2NrrKDUpMQMXHrA
GE05r0l4yKyefOhL2Xt9ox9KX1OQgNEWIvYVQUd8FDBQ4QHHKtqDYPKBkNHwuVN5uifgeYk43r+G
XVyMEd4ibm4S2D+WYRP7a/v3WOCBHR5DLiV6thRVOUAkeicfiUBsjulzQKDc6fSXKvk5Y0MmuIal
XWBuy2wwuryCrgWaLb4na0zMMZ93FDgGI+t0mJVf0YPCSjmJ6ZJcUsM4IL1+QlCQ/ZjnQ8ev32zC
YezQ4p3wu8w0V5QHI1U5/LQcbBPPy5YKEFM3WLOnbctNJtG5wbmUUEALhSZc1ofTKZUXRZ9hjqJs
rrYFF3DlCKqEDOi36rmfqvcWj94fRtjwpbVajI48H4RMwtT9QkRJk8D7DeI8fA9Nj9nSG1Acg7st
qKMrcFWjx5CMkLrc9sT8SXHo0C9FtYRtMCgwdLko1RjbDDLnKQpLYWwiKCrwzUq0n6MsLmzCNVPf
80lT2Cph7uKUkfx7QkFi0aO66eithFQa1xjRyYBRl4JCemVUi15+ShgJ1UJunDTPk6CsB64geiKv
TNFq0skzp+iWOui1psQhcGElbcMZFpctQRy8QEJNJWTPOL33+z0sAUf0dfcTSB9YRzDavrwx11pA
TiKRpo/ev/03YWnPi0p0OaRPB1HMzPdTfQ5HO0862uTxoE+NuMuy4jwGlkMJfnO9MDqrAg4yNhXs
P6rawibwV07j3Iv0AgZqDPNMZuR58wcg3RhHQVGtv11UtpC/RWBbzqi4nIRu9CvtnN/7sy2oPOdp
HfvmHzXw9cDhK74gycEi02pNWh9SSfFC5XiVxkaybZk9LwtUF3kw6SaHbuqluJGbRdM8xZX6CUmo
Z9HGVuEYHIVPEU1kjmVmMeuL9QI9MhVHHfTnftubdryj+EUJO1h+XXRkJuTN0NJJGi9ATxLVBz1P
Xn7cPs0QQWOsz+/GuOWwSjtRbw6xCXXpK0Pdsb3GxTeBBbalMCcontmAftHU0hLBeZ5lyvpZjhek
FDC33D6FdUNVN1aJnO1+TCLWvtXvFfht8CjCpF9iXuzJHvu3q+TipDRdPXdbLE+y/RzR9QCDOi3C
T12WSQbt6hQg5S18Y9yGE9gzfYx85hoRuQxqgxbsDx+bGeRdHLcISaQd6Qhw9eWn6dOTv84+6D4E
6/ag9ccgjNnwpxO5IAmDgzqYgv0TOUmcXy1ptQRHQawVKNwBi/Gdc3AnL9nu23HqUP1064Mxsq3I
ek8WCJTMmD03OL4a8IPB88xryRWVuF7pBFiUuwsK8n7DB/x6X+LlsopjYIiN9EVo9E25O5+M5yHh
VTgD53Vxbb4H+htNmyLt8dofRXowAmIUn+krXgJARBpJafZLFEz16AdbailVPe8LDjsOoxvydf9o
Ut54gY2Fuft5AuGiTf1e4eM0H7UTnjyLGt3C182lWrLcniCbmqRKdjg2Iu6rJ4Uwh7BLJCm2E1KD
wNEiNu5Va4d0jrqYXjqOFZCPxm337bs3ME3NV2ZftldXn8k4U6wO4bkHmck/em5keBGOZyDzYudt
XGCCILn/7qjamDxyF1zRIsE1oZRjCLHNtW5+MyeDut5tuJPl5fKtCDGHOl7SuLo14LHzbOmJc7Te
84Fs9yw3WNHJ7rBD4gqkH7ulz5Io3bpG8DjUHEfHHCputYRuzor2hTBSe0FBhNKJ0AFTrezZBpqy
gZcT9UAKqj8FWDU/2lDtwv5vfaoB3aynaARmKry7lwIhDgH1ZHs2AuT9VTLTDeEuoPSpOf/S8SHm
7q6LEHuxX4z6goORwFxzlfZmN7d3d0h7TxHCUmMjl/xfpOsNJmQr1zJq+anQIbPvHCPVZXI/j+7q
MECctobn2Iu/NCBIkL34W7wpwRC+kOFThzIUXLvrIC2VDpBcD5NiUyK98aV9Gjais6KhmvFjffeJ
/kK3NcGoZaaCzfguDJaPm0DJquDR0vjZwNKaAlFCR7jv4u0LQbpG6uW58452Q9CFQmp5LCsU81Sk
Ph5JB7LEX+9PRJ3O4dgmQ4iTwcFbidpv0NtBySerFISbTn97DZW2tupjPCJx1TqQd/yA13jnzVWP
20r3unqcLn58+sFlGX6rqADUN9hYqyzYy/wy3BH5HLMnAYHGC8+xjp96zQgl+qpoZtza734GeFxd
mkXgS5DDw1v+RUsDk47YazYSJZLnt3yhEAQzUT8WQvlhk3bDV7FzKCEOBQj1OyfkLJFzZzntCiKv
m2DMC021gkZknfBtYYhfHwB4LM5ZWztIAFbP7S0Y3fpAn102Z/7BDgx+4NX35P1XBsvtBt309XWR
o4Th964gIWmU8tSQDL3McfX9zRWPON/9ln+hujj5egj65Z4obAbm29jeypYLqqkQayVy34y90sS7
evoFJ2wn8z+jcGePsLtaQpfrJMiGupQI5PVC0JbUKv0eIn8IKx5MFs8202+mreus+A5Esz0scvSE
EaQ4DxUyTTckqrExwETzVSKvj+lbt5RCdV8vN0/cj66iXUQXo6r7054fDR+UEl0ez2QGhJyztbqR
8ThmwNuySlXqSLsEXiHZ5i/k94a+VUbGugy/tlIy5RNM9d+WA251oqLbpfr1/8kdajOqV4Y5UpDs
CSBSFcgLmvtf4vR7kCMv02g2Itkjc+eDRHSPbY/7U9usui0H92yXlHHe1mR20Hn79QXSt3yCcMab
JpeEU0jWBFY8an3BuBf4+t1ddeLonFDVr1wVyx7q3Xb6Dc+yjNBcUsYpbovvTEiCi/sXiAEsgBTb
QKTb01830kZHI1l3gyhK3SaHCQVxklDBXGUpnmUeNrHGOIbnuQugfGgOxi/KcalIGrcAgawuntEd
ahg/OEQduvkP2yHiTkydU2DZNKhjqxcNctDlDogThNWzi39orCP48Sr3bdtp/cuKH/LBRbXMSp5i
XBM0jZhdNIpBNtVbr2/j6lbOapU0NjMiq5B322v7tHFkhcVm/8VoYjB0Dwb3NNvu74zgj7O6pj7E
NyFUiYolq1OBoXHspf9R7wK0xv/shMi5lZNiuqouvr453Ws8snfNspFpoqwC5s67WDC09HOQ+Wcl
aF6tWYKQsV5GzzGstS7kjSLwgZV9piFSDPSSJb4+CwbafDG+OXirS4iGO/p90JUbyFnIMWtYXXSP
ufhiOpc9yWDZXkDNJvrMO0q73WjjxkNQJVPxiDYKO4t3HEQS9ZRwGbDWO68VP0Rz8x9aoyAtyTqU
M/eAN+9GjVGQOcpgGE7uT5f4W07VnJboKX9t45MPmCyamoV1tGjE5M2G/ipNABOItLuw/8ogaIcA
dM98zDgNMZ7pqw/58OIjOj4xqhT/GiWTSeLP79h7s7+h27l/JuhQlBGUIXdJ25/0Y7KIxJtfXtMx
DlxUCdYr8nXObElfu6QzjNtIrK7Q+48sgXcXKcMj/3ahR6bhkGW6bFFRSP/hoHmeAp4k9kPuVhW5
4RWrZrvTwIkKtdn9RbwqY0tC0FMzasUk9og5q/VWziQlwMCrukx+kt+BYHwPv1B82wdCYLdsWYhx
TTMd7vDhQjT2TtCwpTUd67AlKj/2AMcUy1oZdApNQo1Y9Ehisy1aU53a/XUunIa0VUGCZIlxCxp4
G+Q83IorKGmlyb7YJ2poSTMgZdNsKPtcsuikjwU8/5mK69uZejA02jX5egQhYEnwpNprXmhaG7fs
/BlNTWvuZhRdnDb4BfcDH3ckk7GHxPX5rWNa/M/CUpcvvnG//a/yie8CWt503NQgFP0tvYgs0vAI
XXn6iXOff/4+epSd/RI17sZOnJ2W3a2YLd+B8tYK5rfbhgOCJd9qn03R/MZzAT0qtPoSK6EUsdck
X6UHJHKYiDXTGr332UYsvU9SYWN4DODEzxX3muMxZHFGAY1DLE1c9zMIqgDIT8fU0T8tOSWh8g9U
l2iLaIjSAqSA7IF6OEd3rvqbgN23pEIG+2QEYfTooKHmPR+mJihvAMnI8RRDgRnaEoi97opXuGrX
ZVSp/u3oJ6MufEqpxaaKdSO52LHg7CStEVo1h2FKetfAZ3omcW/VpQmW52JmnK9Hf4MvchDilUdC
d8ekG0NWhGTN2ReAcF0Idr3mcEgbQRXviI1XUIb4FTDKuA5DhN9gx+VKRjD83T7tq3ELTe3euHlw
EPXETn/R3v9nhEoRW4T2Lwgi+AQJIPL1DmoRjpAT3PJYfMh9u1smN1lFxBuEhbxgFNWKyxFSwdrm
QFeC0J6vzVpbqI+aE30Jz57K3sEhe8/WXLZ51u8SujVnXYnSrzACaVq1QMt52GSJOkgS4oeJlL/x
TCt47OhinLqkUyqAQ5X3jzwRT3PUGzt8o7FKzK4XVzjlh1Ml+ud1iscjv9SiSJcm04MRLEw/fiZP
Pv+Uqc23Ri1iJJo72KApVQ4yZzsieJQQu+7xUWNxu/98YiBBOLORNFwGRST0DZKOVMeFroZ7zZeY
wFJg/YR4C3kENQ5mgBkVg/BLNNTg303wsaJ+l4xaHOze5qf4GVtFDT70EA/31scFHzwrSfgBHn6E
ylE/B1ozD+b+8vNuoRO7QxAdhu1QqdAyhxUGptUHMwT7CbcIEQWtEjug3Ah2K6Had/8iGSm/U+CU
/4c4PhE27Q+zddGJJxZLM6DtodqIzDchrNttc2f+owAlui4qR1DAdnGxqiA3G3ExAib8NcQf0rra
zTnoTh1foFwi7oz0/mS41o0sTGdJU3T9z1/omZIZMuxYzsw0DdOlYEK+xQGPAy3R8eW2OM2s62eY
8ycoPG5fwCt9KIsNdSXYyUMkWHLbVbpCASoackzC1l0GKMtBcLqQBHBAvHMyI/OBb6R63wgRV7uP
qU6+IcOzqTbrmKCxntVmEBuDnR74CKoXehb0JldFSmWG32vZR/C3pBq3yd9dlEoG1gC24wY20RJy
9YY+Dgv6EcWe4sujbncKFH/nxvX+6jInVRhMK7mjzF+jE5LyEHg3xZke5WBk3n70MIuqRSLXflPz
sbsZ0f6BS+81J4pl0RrRL0BGzuLaQL7wvgkBq5oKw6b8RmfwRE3jyYUD3Ni+3TZMLWveEicWFs12
FdOd1zwBxIT3+UKYXAT/yXUZ29OgSwGLF8bjgmIhvfhqPnI4u9vjA5jJY0smi3aS94q16ZM+PvSA
I/zj7xVCTcbM8CBLZ1koo5fJo20BE+H66RNnD+2V1yS8jTzgMWGJTye8OpxfAt5plPFWwnxPrJLe
xTS2SBp4/YlWIQyB4TXkv3XA4k9TWyqdIXbwb9JcAypsD628lzE94n61AktDUU1nzwWZgb3B3xfO
HxOjpRcDiqVz4jMFZOjQNqABlWVEzleN11TABmfiu1BCJ45P2Wuss53s6YMMo23FzU0ntXLfQL3/
k2lK60OprfJ36Ly9IHOE8jTOVhRvkIzYW3O+GNeMeH9EA+xSdmQvofQ4jWI8CZdtUhrsr9khb4ab
8AI0Wo6JHZ1ukrl7UAqV3fmSwK9bdc+cLZsQ0UPNIqqefn1NgMVmfnvO2qX/XQPVxkcr5C3OSO3j
B0+5tgN8oJl8bZjgZJDSpbOXjpNMp0mwHOGu+zoIhu6gnoXcVbZmdXP1ONHmB+wjUaWO+rZ7SYfo
fuCNnnRf7JcZVtvmph/HDJA4CfCvDyEVQDUDyqgkBCnIupdcG7cjJiyA7wrm/MbjlC9ebbTBh6ol
RJNJx8TI8IhgF0DQhxLekY5gM8pRFSLKhxMrHfgBwIcHavsgv32IaGGqTf10LiXHdQcY8LW1SDnq
829ndggM0rA2O2018XLLW9DuYnkbeVWM9BCRjkOJ0XSehhDWpcqh7Qqf+M6efg4OYdRVjQCMvsah
tUUU9cWg+tXc/JyFJPISFOOiN695wlK3iVt1yDGywYUnc8KD7WMRF7fNwCFJ+Oc4CS1fFlR2OHWJ
WNu6sVOtkxlc2QlB+7qw3Nx44UmFMNnhrG6X74N6v1pz9hIC6T1I1Et8NhlNqrIOCdawOmRcz7wF
pqp4sp+Z+lc+i2Wd/6EmpwSHFToQbUFl0QF7cDm2Zf+wmWF5yu5wnQdD/X5h8rfdahihl4Qi+1A6
z+/cwkO1JyoqMDtE5dbU9xheWrr0AUz7xf0+YyvpAM+P1ff/B1cjG7tCb4lZHIhJv24ZVy84Ckbq
UEg+0w8gZ+hbFkYoRNvEM8JxeRDsfB5+sBCNReP+QVka7qbMiiDeqpX8guPipmBwJHjPKykEds5g
VCOdzOXZvCfcgpCDSzkNeue6KEzvCJr2VxcCzRz7hKbkTmGwsSDtFN7EdCIKo9FnwDeqalx8GcF2
4yItU61VQZANSCjHqRe0zk9YSnwbrlKJkeiMmXR32pmyrZSkZH8ySHmWp1RQBUjzqlUEElGQxiJg
9Vfpyn7QIT56kWrDfhmDzVdkumB2Jr80d2eW4qNT/YiY/ypF50GUfFq9Xeh2cn0lIgokadJscYDp
qnsT9jS2eX6rm7aWanNso97fA+2ltc4W4iNdw3J7w3VN3yWZIJOy0llmsbxdigtxgj0tS25tN4ZH
6nTxmRi3s4fzvu3JYkohmBtZk5YGMlSDNRaKbWSecLixXWD+voyGkI78rLA48YZR0lI0u0t9lM6/
Ig5gTkFZ1Mfq6z+gHJKsLIwnB9maMZIPzViA+lazpbTjwFDcHapo9FJ+PSHIcUgSMiIl6k0jG4If
QBrLDNFsWX9PAh9IV/3eeW0HFlq7zlc/niKULbIFSFqm2L0auJzS4O4b68ZIhwhtvRaMLi17M8zG
BKtFFLqN44AgcjOx15ui8UyBlVue4me9l92L0uuZM/LO7mJfytefYZ5YD7YrwjAqftF2Da9iQgh6
oc6s11C3N/OKG8EciT3R4d5GQVpXag1sR9FTQEX+iIESr8GpM56u8dIcFium04pd1v+GSgdOxNtS
p8T92uOVzIfuiP39R55/rW3bSzvomSLMPs/z8jOg85ByU86wDQRCatw8E1PW4D1MfRrH8RGt4K1w
dsxPBUXNDrsYroVHelusCJxU4BHyE/oXUUX/ViQBTZXvJmb0zvdHkgnSInWgPe4F9yn+K7l2EuZc
mfgVZ8ykhJ+RlqlSWBb3EfDhfxy4/SF2MjHOdYWtHZOUX19FGr/0IPGj4RgpzdDC7fdfAcqxiWFe
CMnp9NgebLkabCNGIauq45NREtujpD/tVNHMavfGA1cFUbK3wT2jKGM+EZAuwTC0qPNlaMrU+17b
kMiBTeSvQWtE+446v7XoQnL3NRoVsf1nWVL8tFmsK56AwUCCXES+pAMFGtKM+T6+eXdqnY533tHN
u6X3EypzB8Vnu5eEL3/rTdHBJ8AB7E9RksOqA2K4HounY+BV6FCVRUwDkvnYImx5H5ogeTsPEUIB
nOrqFCQyjpvf8+H1Kx9qaEwSNM8P2V9S0ptllEW6jD/MXB0jxmUqQfRpVBbIwXoxTxGNsJ4DqXI+
4YEaN2TM4vID5pFmMK8NwvlFTEsHtLiJHMQ6CbA0RHZoR0pENdBoNEEUvS+RfKvRwqTeRVRZwodj
RYLvl4YDADYn2kgfERjNHfI20YEG7cEGz8LDuBZfnZdHQ4/0oY8XCcm9n6huO2AD9P4xpPB+rU3q
zIjrSha3TTkSLeLlSTBlERfaGrQ96wQ9RHskVyDcaXGOytE8fhdKiE1nCeTd4E1Sou8FzX+c2sk9
Z+Iho+AykYBx9cGY4B+oQeGUWFRgGfAvqz3HgnwntaZHI+7HUUlAaJkGH8YYjGCA3ybnL1YxP07Z
WCg+VhT3uxDj1WOv/PnmcN4WismYcHKZGkTcMCO6bwRhwniRemp29pqbQnrXsG8jG+EDrOUavzlr
5gunTdsnEBJIdmEEwaamf2BzcaYU8UGt0rrOUcpUJraCSOX820XlPfwCa4ipfJ+j+g2yktETN7wH
1w+VjcKPDsB6/cknV8wPfCQ/6D7Xhb7C2V6xuJNQ4C7u7k5Njw6VNzDUtMwhd2F37lVYeqearf0L
nfrfdvQ+MySiT3AYFuS1kHFFkUg+1o0w8c94+U1Ml5TtP2jH3av2elVzES64zT/5YaRS6nobLX1o
4OJTEptv1n7zSk4fpUwXXhMONM+yoLujFXBe0+TdExw+n1tOaUvyckKiRnbX29IWV4LPkUJqSbe6
rhqAU4V8xErJSZMPafK7M7r3aIiQdH9KZa7W23PXS2bYIya5spR/qM3eQoSBQ+hBlWsF849X/RvE
24gUC5PinhxYugAr9SY05P0cENyXh4rq1kNUt6KzAuyUxpetoBQ2NJ2UIp1blaJIYiWuzxbPl9dZ
vYlIbp7m1nvdoBvi9wogEQfl8xXwVm2NDljs8PgGrCjmtTkocbUGn+rzdlw2EuUQi2FfYb6xX78e
elixw0Tdn4qRB6ejeP0dMwAmaqR6GqD7I2W5a3zBXZyU0kg993C7hmF5OfnYtjTpmffgBYL79MG2
HohfotNztiPzh/CARNmRIhFE1PUgpAHr3jigij1y8+V9rNRFjqln4IL/uV65pQ/YDVGiUZ8slmyG
o2zWrW831edKZ0cUz+hU0r0iOVG/hJYsBppqul1K82LWO8anN0oIyHAMXUH07PzL638fJGuae6I/
rvEaDZsL2NwYey1FR2Dx0vBl5ofBRsBjGCjbGL6NwMUX4PhkpP9U9c8DgVfOaPOSBbwFCSbSsu1+
yUwh0czH/Qhqu+FiLCqrjVCUI6tNaNjRJiRdOBKb9g/RS0Ng6C9y/twT7M9PMP9ODZBwxUX9hUrB
fjcwjZUk4T/m6HlWcN8aEel+/or8awNWSx1eK0Ay8Y6it1+C5LUW//ucJuuHwTtISsFC0neKorsl
Yy+JqbBH69oBvbostD4lqz62kVBRTW5tfjhm7XgzNRmHpoF1SeodKHK9yYSG9cIf6mgd94lR+1uH
ztMCm+CQSoUqbFjNcRvLdI4nBhn6ixAcWsFEoa0C81Shg48Ws0OBaUdq4EJoaGnol7Gjw7eHADE2
UR6hw3pP3HIMUz/5dAmo9t38um1R68sdI5XXuf86k2kX1+UNTbkukRHmlAyDFo8Bwbqp3wKxVT5V
K4am9zXMiSagO6TU1hkQ2u511VITs7vEZpY0Fn6uYsy0VVvEjCu92FqDKr1cpt2ZeeIMxFub9M4x
lN0xGudhCarq9+TO2kLFBnSbjtSiAHdDOnbZM8UAPSJHedYa7F/iy/xENf4bFj/39wIhQmacPtiU
Gm1Ti+yV/yyIJht+X9qwW5dsHR4bkEOYgYEVAHJVwsufWgiAkFPDF42tOOqxJftaYW95naCxCDwB
mjjgGlOAb/IJSX4x9SerSjUBIb1q8iguw8U5VeTQfjptTWWizN1Am3zJRooBaORzRQAH8f3bYtOm
Lw+GPRVI2kKEUjHNCGvhuqeRr/5MgFzsvH6dUx9ajovbb6XqJAxPc/79lYh9x55Y10TK1MD/OTgM
KWx+hQVox+kIQ0Uu5p/65qWX3GBY6SOz7u02Az4iFdo6cnVpndKc4yTKv33YpBf6aZpxDH1VtS4P
vk2HLSNmGJZ9iv1sM5eTiYOxVE/6IpcIu/U1YsABhdQT/EZPKZ3J644IJfDrtdj5kf0dmSly5Cyc
YzElpipC/UAJUimiRe/Y/C55/ZAIIgJYofuz/tnimeQyRMf7YUrjMtatz/KdcAvX6eb3KKQF08PB
W58goKCyZtp/K7Os42l0ZIL5/nYlAC3brXDGjZjGNk6c4KZGWY1ak8f4LYFtilm+7Jeb7nGwyrPn
rYqNbeOhEtLbB1vb382WSXuSGgRRHi81v4fkcX+0qOCUX66ZwVrNzBe8kJZoh9AtiT7BeUdwa4ke
Gva1MVe4O/PHnnuLmPNYeWEwrT01fRmVC4FE4Q68xoXBPu4cVic+42p9/EGj4p/E70ifEqY1hmhf
ptNHNtjNP4AWOi6+OW2RJ3OhR8iy+PNNDZE64sbRjA5Tjo/d79H6zCQI5xXT1w3lRmZqWVpsc3BX
a+K5U4dmZfqHFs313pWyqPp6G08tlipiE0MANxXo4CV4mToAqCeTNA4NQULJ2jtXb2prO5sYLkFe
eKfjxwprcJV+7Jca/numq+HN28XqXv8UAqdF1obkgQyZ3C8icVe1iEFbeSZTKbaRPZ3++JIp8hTO
UmfTrKVZ27kfgRQ/w45AWf75HdQi8IURk3eGqyuMOu6EzVqaynfdgIkYqhtDuj7p+O68tX3/csbB
cqsRf0ORNZptLY+WK89JYsi6qICFcTm1lSqKT5UyKr5w6TgoCV2WedlaAfwXzryymWFcbgb1yo5I
geqFRwM61hcaL5cCbtCK9o8HPnF+61hlEF+Pc+VSEAZ5QcRULcPaaFIium5qO9fT5rl8dZHi3NDQ
yzP+p9rAcndRXEA+tdTNg4BDebuUkVfY8AR0TY/jQFQD1W9FShS52AYDIpS061jYVhI5N44qWRR0
6njGqk3MIhQT3iSpgLRwYwTwxE4beSOchp9nd+esj/9ivpR4YN07KXNgLe9pJz1Yggd4MgxIZDT4
jIEwO/b7Ou1w1/TIWMy7nkNkli5HMm0+AtzBwbwhSKLZ3uMlg8Jex7nkeExRWVn7wsieP1Lzt59l
Hwxnt78pN8yO3Ut8Q+t03MxogObTGW+6lPojvI3gsHvIJNPPyv3ILD/zzyihhlz9yRLsBFWr7RRK
9bSreHQ0xNGHCg0MJDoEkPtb/zZN1SFaPQV6L24bWEJYf6gAqIAyVvE7/G/LtIeqJPW/t6C76ow6
YtDv+kXpIxmNcp6feV4ueQ2P5Pp0FYhkfHhdN9CvB9eLMG0jJvJ2QHHiw5gt52uGgZ7MTyR5tBUq
lPhSintWfVnVNqx3xjZyZdcj57aCS4DLZN95OluVJz4ahW2bysXCspc4y0FUWy+qpYJt7rh2Geiz
KiJB1/qe+SqjCfZEOlk0AuwdUiuJjUF0vdSva395qrp6lRt/3IRx8Q+SV2alPeLPP++ZtdIIOnph
/z/twFxX09skPXu7JABmpNK033qTDen0OZEgmeIp/CaYB0+Bl3WfLDxXyk2s3ckVm8COqr8c45pU
E6tX76zEIVKPqvG3be3YBHDCgfCg5Z1AsfBcefSYXs1+saUOBqSXb3tY7x+VQ3seXJSW6P2ZniY4
vFI0aMvJmrhrZCghfuTmkyV2YENEeyZQI+Vj84g57o54iSyPr3Rkbe/QvZs9qyz/urL224gnYZM5
bvoQAexjuDVS2xEaKvyIbezRMTdm3H5K3iEzGbCgMMxKTeIgUqusynChdpKPmQs5EyZR0s5XLCGS
SuaD3gTGaQHBON8AdT8n0JFBUjFbLKStmAZDCv5j6u7Kc7TzW1YFb0e2x0ugvT7/OjoVrqzSRbT6
N+ICoo9D7v5Oko+n/3l3Jl+R7BHbjA/deBuqgusrmK7ZaxiJj/ryNGHYr51Ak4LWykzs6Qn2ftcD
c9Xm2ou2oX/LtLZIr6xmfBzQfJAq00RprdiNFjZhyzfu1JOaHoSZmEQ5YGtSqOJircGqJuYL6bh0
CQYMYDpwGOBinhlBK911dQWrCpldef7C5qyxFBFCxltjSDtE6BrYOCPPeD8Gik1wXkydtYDQ1Skp
1WeAuhj6ROAAj2ZADg07f3nt2phngvpK0d28sZETyOTrKFPK9fTJkQ/tB4jpesRnL5z++RC6EJQU
XxRwXER9SOT5HBg4pnb2W8zSMYPZsRiwI1YHBptZPaf9Rt4cNrFBGWNeQ+suIis5MOHQxGiQlDKG
7P9erFD3lCpbtWLGoiFlprSoVljsoDK9NTGdZmiGAa8QmQmNvlbz5VgkZxSUKCBw7dN7DLjRcu32
4XxrZTKpgzupEK+z0ozLJZcXgZUHxF5frt0OwPYSNcAYspmHYzpjie98TU+JAD/1+NhzoAPveXFa
PhWSIUPC4Czp+Gya4q1iz7lLNvyK3nhduRPrX916VJ5HrhZ8mj3lDKSym9F3e5sW9tUnFVjA2RYF
LW1ad6IUkk9/Jbsxn7s4OC9EZRFl0BkNRmpzCIqT4aUeifDXiRLMKOaYxor1HOvzcQ1n7H/+v/vK
+di5ovrb1JB4cdWtB0lmPN5tp3OqNU0M/SsPTjpaHUg1X/XiqKauZar3JcifuK9RdsPxtgQtSt6t
O7xglxJrEnUyh5IzaKbhOh8mSK3ELAe8c1t17MWgXGE8CIbGIE1bICg5ZOxkYUxd+txIqtxVsBlr
r6GARoD9g13WoPnN6DlAQ0bdUuJAQbTeGpXXzQUXBpke2qm2Hy5VWO2ay17WYu/nOVWW3zJF8WL5
Gdv1O+QdFXmlqt6Tnvsv6v7x81nuewVNslDSR6U3NqxPXy/m6D7ktWLSMgb0r3rQ4WWAQEv+7KGp
ZwfaOwrPfskvf6eDjhtYgPrrrbQw3wRJt08bx2rujYtkx/6SP4lX4tB05BeGrcuOLc3dUne62nyk
F/pyrh1/8Q6VpbycfZgplzLnWgfsS6U2yO3n0QSQxRLeB7gWQpC+uLkcid8znjkjdYb80XDfXxO4
N3JwQRL+P4Stp6HV/QRb7pXvxIcJzl10FsiOia0ZKwcs+9ycoayjLcDkdWX58PEXCL5H4nyZWyd0
CH9Jhy81xOxJikgLrSduY25jvX7irulR/2UCAF+KkHadb6VIixfxLTKQXIrNjzgpsYj4rZCeuKUT
P/PBu4QqDLp11fGDM6VqBnm0mjq5dn2mCrmezGXUV2JUl6Thh6K9+mnlUL4ozVMuI/NytbEZQLy1
/ZY/QNrneuqZerOZKCamHVjGQY6mRucvmEoY6hl8vU+guthxZMXaVmObOtVuTeNfW/kTpB9WfnUb
m3AUxIyXq5wereixGQXN+8CIxH6MhURm2MvlsqfFZ51Orjv5/q2PHgWIYO97vZVFdEAUDemjsWSY
6CX4uF8Hj6hLBb9N6wr/cyp/YbsEis3hc6pF2gKIFHjJtOtr+etNW9AOFwXELi8N2iPS38I+Jq4S
RBJD9S0IqA4XUCAwuS7+s4dEjvs57NIKK3yOhwwPBx7XYtuFE/jHa/LWqiZ++tWaG3zs8Tisipy+
21xw884QKfXSZ7HFJAB/10E4mUSypoQG4Uo9A/wUGBVkkZSHebbTmI60ix9zJS8GrYvOR+si1UpU
emwB8UX2+0VEq4ZFTTbsEdur1RIRpQYQd5tSh3Xqe6z/c0khJ3Y5k+VUhWo25SZgfNhc6PoVJK0S
sN7zWut2Cn9zOEPATshCWABED0PxmUSu30Wu84qBdVQj6DzucG71ArZGmVVWVGvJivBn5JznL9xk
nHr1+HZgewjy9upmgvPx07rrTc12W1tj5Ogwph/BF9s7SeW1wd7s5bkNu8si5xk3kn76X51tjv5a
HGg6N0AqkhXhouGw2BfssZsoWmBM02WTRuK0AdLyeEoDWIUIZxKeTQ7ZC+GEJDK7bVgQsbamMLHC
3xRebYatkL1mUfJiBSp6A/E+NHm9K7cl9X6mVVqhoUJrOO4uSgmGdkuFOD9YzYUpkdkDF3L/0fGS
XQLh67g38uEAmvM34buV+vY7mJxVGnP4Yn/wgc0Y2hdIgjx5jUhU/HGqz+1u1FFq7R6Talqib7Q0
8qsWCndEdjuaMGGbiPZlCxODumcY/2V0z1yfbghZeF7L/aICnK9inaK6KKftbGkQMOqWl4xXecln
LbSfFFHbLe0zQQ3dfx0dxJGj6mjhNomT63smDMC1ZhLVDWhx044gQ/ryvxGTgjnyBj+B5Exiwnk6
6bzFHvgD0/EExwwO9WdJWMKaJp8yNWNow09eR2jk9Fcg/dNXC4yOe/M6PkPxILGhHW1GPW7ejzIS
22jDUat8u7bQYdbS4QLxFU6mkw==
`protect end_protected
