`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
P+5ys0V3gDpeppJWzbbcg5x4Et4BL6IN5B6TYx9R4w7tmtVZ3OVS3LOI6sRsk6EcEhafO9ZfAn+e
+zWD8hgc8Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HCLNwdh2w4ny/4ZB/a7d665IqrnEGokAOxwFUQQGrGh8CioUUGqc4u1EQ6phQyDrHYK3NeCFaUav
5SRU/JE3vPJSk0n9BN0dZu+QKAInT1rhzL3Gb6AP9QZBT/bOOaskNvBduPDfU67rIf65jXSzrdqw
RS9VGidO7S91s+cpVpY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eb8DvioM0ppHhQt+iCNsssd+y5ZcvmEUDZUim3W52jCwMHqoOHhAsl2TqhSeuhnLk5pA4+vxw5iN
aasMB9ONSTtbXkrnmuTPEeMUKSyl5NJPytLv3SjMQuGdnTJ/X0NbPJkv7XlDY0i1fhi/Egz1tC6e
EZREfE8bJjQgj9ZQD9JlZTJIqMsrzMcoFRrH0A+wgfiaFSclcnXmlqAgiKTQ8TlUSmoL/ALpNkjg
wBcHVQErMzNCZ9eVVuI66Hkw8pGo0Oj/T91Fzi1rnzvwX8s9N4+4HGhfqFL9d+hB7SlbY0iswovN
JOd8KVYL65yJtADLIDxfe6A55WEhIlh/nA4bMA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gFYJwS2gS9caVWWzK7hFad+crZTFvR63WxK2VEswUWjhsDL7TjdgBM8rIpdWnVD29QscXO6TuDw3
Hd7twnrjtoLW48hhHvAk1x/zHJ+mC15KJxSs8hxgJcHysHqGGVZS+wbDoj5UXxIuRQTsbP/H51X+
8ACPQjrb2AHWEzra9+Q=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rRWk+brljkU+cdzTo/W0rlS61KjQmks0jYbqZxgulf6ZAH7sMuf0HFycDWlWwQBtF6LPxbR2yvrI
EnCjpR0chBoPVOPRoIgbqFlemWaL2ZNBm9qHCkj4x79643u4LaMnf77OhfKk7yLdrzxi8zwD7I1Y
+8aUAXfaAdMkcjqS3ZY7RAamayVdxOeSuSBQpPm+WbcV0kkLhdVTDlzLmI6lo3vYKcUtEWHLCn0/
j3hnqR2JzHqmQnL4TKRQMQfC+oJ4wzzStNeb/P+aLf7e5CVxfmiV5HDUHE1eWLw7qRXFFsEy3P1l
PFQ55Fqgv9jrikJ1BsGqtGRlhQM0jlSCTGcWbQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9488)
`protect data_block
gF6Yo3Y+eUTYM13sj+7X2x980VS19y+kzLwkQVqyTyNG+r40H44UK1ypzssZldEsZZBR/iVus/NC
xUYRRo6VMzsaunMaQSn5AT7kKxi9tMGuBfwp8r04M7cOxXEt6vjESbsSX4JDgR1Co6EVIcLD0xW8
KzoYW/bGgGqvrbFnjq3XfH4pr2d6O/4T9bpMIeYlZieJj+0otjzhjHc51CZGlipKKjjJBwrTA/od
cAhVDxSrh6KaHnPt/0jhAX9m8wDO2s0Y1IRMJUCFtCwkFXXvF7cYea+OlOk2Mfu62IJbm+d2Bk60
VByQWeAITPCoCE88VMR94zaUmK7QIDq6zmwXXnv0pYjAuAw69HUCPJjD5Sr0yp+pT2axhQjBhEDw
x57aSmRZtpBk0EWOmDpOzR5m9x6d4qwf3P1k/W3aD9rn+FIisHyu3L9nR954Dl0uDE0xZKL6ktXO
iBnn69r17VXt2oIIrz3W9wcazBiAaoa+8BF8e++JumHw8fGXZ0z0i3phHbiCf/U40Fegg90fz6q5
LiJfLOW43NfDB2rb+wpq9TcXTLDuho29Np9vy6gJ4i6swBzJnQRX32GFbcZZaWJgaCbIQ9LY5Hfm
B823MByAxYldTpdDk5AV2skKUP3QbPjP+Nym43ukW3h2QVuSiS8fCiQDRsDCJKaq/omLUh8EonwN
E+Edh5H+FcFxTXXyN7dEtopIz+4GQ+/2B6qHr59f28wd9APrXWLzMSwfdxuD2+uJjql/X5cI+4ep
6b3shBxakEDXwCIiAn5Ej43cKYa+XOfkyMl6YhUN0owrplWGIxIANsBZ+v7MNOSmucPfXv/0dSXn
kaEJl6HpL/GbZxyQf62G+kMMaDc424um+RN5lDrJVJ3KBZpUcpTHlyO54kN7KjYBRXeTr3b8eDVp
37b6/mmitAprx8ByvbXJ8X2eYeDo+TtAPMreYLXm7m7/yqd1T24xQMK/J5Ic1W+XsK6h1FIsz5zq
/2EjXH+Y5TaW3XszsjNFuqrLA/iOfaF6kT+AUvEcXapRxozg8tAs81ppqtlux00IiKE4Hkn/1S/5
rgcUD5akvldxRtboA+0n9FzlC3fbgqKEzSFi1CFyi9GgGpYSMCvPPnSruzoiePDAY8UuKBiL7itz
JImfcYPS5ZugkzXb2YtNM5up0oHj2ikga6umBOUZQg33jIsFSWInHhqy9Tsfa/RVSbSRx2zhk4eH
YItniX5+NzKD/1PMYxH838azD7m6oqBQpbSzJLCuks5I7rDAqB9VzCEPGk0H++ZuaMY5T3LENAwm
c8vV6vum9M3k4MXVoDB+tpxg+hmYQfr5/ZheV319iuC21NrQ4hf2guqZmakbRfHWSH880ws65FV8
o/PtYVNxUOtJNMEDEvGA6UXPos5U6zA2q0vNu5OfEGCZQpl+lECeqbucn1DK/h7dJftaJ5SzD5Hj
74TAQtkNmBu1onD0oJqcCa+37ak8v0hiy853J8BNvLx9rlMtnk70o9QhAStbjgyN1xGPuGvq1X9C
IcVhLnKR6Gm+jqaPh+vuYPtfJW9UKVgirYaTJIaRuM3+DGMlASPX6rlMcn/LyLO+G7HC3D/7Kpqy
GunW9ehMk1ePkzoRANSjDO2kNSVUen7nqGqr2qus3lExOtNP5b3NiIOC4S3zyJvxjA4+COfvBO6d
FgNoT8FKus/U5eobqfswrlxrX2aCSn6hon4/Avp7mjHKB0TmayVPXw8D79x7DIjb6a8OGY8uMFjj
IYkWh+eRWDynbnhwqNmuf9+4xDDcQbpVLu9j/jcOQTfgxBiRiLkQyS2kpB7fOoPWRCcE14ehx3Oy
v6/tvMkcB0Vbf6LVFu8mZl6dQZwNhaV/U+RpPPcHPS4PkggpGPpy67I0DDObxcVmVvhMSb9MlFNs
uEdgAQNEYzjWvnz21+GH+nUhZIWHXnsG5rNsEq5vU5Z+EEYcM3yC1MphOemp440rp5lfvZOIBg/E
uRrfb1ziPJZ+Z+rng4AwcXZ2Kg4yMYgSnvlANBFOmD9o2ZZCqZf+ZmAMbSbUNL/v1GNuE0YxduK1
p6Yas9cPSVPTTzf3pl4UngtcqxmHEDbFZhl9EkhRL4A4sAHTxaDJ20nB77acSdyubh5SdczZH6ux
rXAkS8MCCseiIz4Y2a794s3RhYXuLBOEMFz+N1cQh89Poqka7IZm8kpwmb7+oYP7lCLJVqPhpBVH
f2oWhU8UecgoGu2Yym+K+Gfcnw6T+XdA6dSTs2BYM9L1O8OXjZVnBTFSpufiHGsEQUzTPf3xwugD
x7eGQs/iUjHHqpjqIPfmMHJfwAnrZjsU8l6RwnBnzh9ycSmE4LdqxpsL06W6RbLTqqIMD9ooP08S
A5HD5cbZvYoF7X6nU9wUbYVdLBG/SRmFn/QWpeuYo24JkgkNf6lY5ids9r5FGLgcw79cfhwjYrzW
t3793oKrTnSntHmGEHGr7J3RjJ7e9o2ZjHL5r8oz78uO08Dx7KvPFDTkuT1HwrfEdXO66IhXX1kC
f3hY3YRDmffnRn4DNmIbB/TT3+r8zW98h3lGaY9KPaW+6VFQt72r2fEK1mC22R0CgdGu7z2/xGLg
DV1OzuPpVPx0US/Atw/4qbLfmrVywp13N3rWtLlCZIsX/+IDdim4UzembA9EREhptBsRWQZzBAYJ
DxCDykOo8INkZFCUBkZ+KIBaP4HTbEUYAxYhIDLxZ7TVNG/bR1CyxxkSpS8F3gY25F+zzbRGtnYd
dBloCQLf1MmxL7KQXO9jSpezcQQKcRHj00/JGJxG/GEy1ZQIS81y1D651Cnd8lh/NyIjw29cntxG
xfFnFMdGmC7Zly/67gEgTHESxwBwqE46lWRz8M/Ei2Uh2i0vder6y9I6ci6T05kOycbWgBGYwdSk
ykAcND3cLuzxHhs9jjh8AzjlW94Xo8Ge56JKCPNOWBEh1RR5PA5QkOE5eA3+jszKAPfjFJw4QlGu
FnPIk2yRWD26FmvsPHZghOa7wMnfMuDZO2ETwhKaqz1aieklUI6nHSODkST7hpzOoEn1h+isjOdX
mM/KDMB8xs7ZEy12bm835FrAFAu+0OC4ZNJU9GLoAQTT70EAfDfPx3Ir8YQBm5tYR43jVClkSDI2
jOjmJN4PcEv2p/mZM8reKDPBLjV8/1Ae1JmvY7LqX8Wzm9gsMDwIoUXKdKrd7wPn8H6bibixoKIL
nRSdcU3+AxCE9twkSREAe8B//BIfnHtRyt0hVDHF4nx2BQ62x+pwSjXgQDYqFU1ol0LYBs5WzSlC
xuzllcz/05Eo47zPFrTV5kBydt/EQvYwE8tXPAH3Qnl/5eS0Dr7/W33BNZCrCaLKFeBlx8F7rG6J
xlSvQZ92Fubr07A43vizW+UDGReEmkJ0F9Kr0LwcDYSWwaXQsnqdirWDpYIEcrWbBc/qPz7vXWO8
BMiA1EKH0pPa79srR3H7LXG4y0k5oOlbn1fmZy5bpAhx1RVXo8aEPRRg8UJVMuwQWC9lxmr+jhpQ
CZ84qZlZObhdz3EgVqq6KqDnZodv6Dfh41ae59ebeu44KlEIzHuNOvcErzJXR4193bWVCvOBx/Xl
bF5TrHisofsv3eZGzorICftIj2HFCC1VAqZD8XAj/2M+mjyGjrJjLGI03PInj17aDefLv2PvUMgn
C+4u4WiGZWU7IYRvQycRpJJbhvSaBCjW5GhiMTZHRB5LumlEiS07Y4LPKmU1VGnuwO2oGAA9Oh4t
h7+hgH5WK95VbbEo8SmyJwKookELlkP0ZvuU9YldtDBruql3jnG5MC1YRAKWMlqC7aFr7Sn31sB+
uBWLI/JAwZUJhg7diam35HP6o0WBP4Sp0P2Q3Qet6/+9oG99aYJDltlq4v82M7AOQOyYyvOeKCON
0AaEIGGmRT4Qysr7UsUY8yoIf0iNSGZP7fNsiu7iE7kR3h84aQj9QU12UXf4kYo415d0sQpIh5Un
FaMdz1iClZQyKO2D3234C3gYf7kuFvLw31DOhRljkm+mIay0+W6SvCZAWKytMlFD808hfVMAo5k/
GCIcVUwxkQWmuDyH8LQlQHxLUK0/zi449O5Yr4Io/8jUsxb5nuGumop8Foi3a504cHPoO5Yia5Ca
UPQ/Ge4wqy1BI6fri8g1ZM3ZgAFWL//eksX4Gp4Mh48bd0yoWtWM7mLooqjqQC2+pVbDdV1C3B2P
j/QSiOyc9V+ihXLHSlf8TRsHS0Tvgb8ePLIJhQBHIksgVTDmuUfv6wzua0yJvAYSnGg1eM+tN92a
udjMt5e8BT3S/aai022wDAkYtoAGNx54ZrXa+js2Uj/Xpy45NhNIbvpwB5mSp5HJzfNx//BhD3+9
qUK/MCgTp+t2yviVFmh1lnw7Br3qdvhm3AU/qCE1lAo1yRBxctL+zx/V6MQq1ht6t6Gxw521DHKe
MtdEck4+lRK8TXNgn67AkHNVUvL5ZECUTzIhbEo08jsEjpV5wuq1KE3QnoV4ybfvtxObGawboSkt
Sb4NWic0TUKzbaghKUMw4kGjsnzQvRZdB9v/NMV96fRpqm7fnUQxlz4WpF3rPOsUfDDZzk2lStBb
DYtfQ5dXR7w/bJuCxg5mJaJcWAtIYvNeTVVUHGBKAhcaJRGyFlFMDEF/wiWw3wP3kohLRzraMpdO
yg9bGMgjsZmtD7KKx5kTr8/W1RmYUQe+xnzLzcF2wPN9fvb1kLcm9SO3SF/IH7xivU/fA/E/hvGU
Hp3jUAxf8k9tIfamr5xXo4yjLpwNc+J0qnFtkdYqt73W8oGuMPRMcWlPM4502EfPQAc4fxAQWliC
3DItPN7hu0d75+JV4oLE/QJ06DUg5zMrRFHNQzo02vz4bx6UIs8UdV78D+rDJB2NOL7trYW9wLC8
5qCj/6JvA2DF0bWhGtrH1LLMPDpuW+XUE680cRRqRty3tzsPRAdCrREmsHl9x/5I4o6xoTKfGr2S
HINGZSUfMNza0JajsCULfr7UB7vRTdIHgYB70YBojSTviOTNReZDJ+jmAUmtCLLHMJs5C1FOqstI
Kbx8qXJGG6NLaj2fZZwep9M+WluRmt8RnPNGJsDltIc1VP0KjKZ4sGuPiTxs9io5Xw3iIRwPbbTO
4qZlb+3G/nQZhgA6ckciu43f9zpKdf43UKx03O8Q9kHJ+NhuL1Fh5UoBXlh00cifNKT7Jwyz0SYd
mG3d0SAuni3BkDAx+g6hUbdIGUc2KNlrX+0eczpCxrZi4XPi3LpDqZFWFEc30+AVuivpX0Mk+wi8
X2sH1hWxbZFVBGB9hbY24gogx2kK8hybC4pcsj4Kz1oWe+e5RSkKLqsmMBIMCF8BV6fGMu8sm8W7
qvBCwVlf8qQmxl7hdEUJzNuc81/xrhzB+cYK7RVOYdk4cBaKHCrdlZ651QOeeVdpLjy35N0ohr0p
3N/eUAbkDS8gRQZynTD2PIR6aRjPj6y6DblJO3n0g4byHTn7DM67jrPBKMb0XC6lCIftbsoQhTIh
jI9/V2QWytzhkOCwV56vFGrJ833lSki+pvL0oSaSicFWVz5Nox0VS4FCm9dj10KJtyskZUEhgZhD
bxL+Hy+YWrFWd6/Cqv9cbE/G4rPkXQMu+clkzWDnhSBIBq5b0RGZAI3M2tyvfkUIAdGRvLZMI9CB
7aZfoeJOfgbhtf8rMhiGondBXxKwXEHatyu0TdI8XiTgpFvzKjEULx9mWj2CDPTj4Ghymr4MKGJd
hyl8Af4qFQmUOEvWwQ/e+3oHHnKiMj68QOOXE9zRujjM/BaAAYxuD9sDAHH0yB1DQduro39vwd7P
7VGuarQlXIwqPETiGYy4BrKAyd+OqyvAGPGjQXETP3D1oH8WKBTdXVC2C/SKc6LBJYonDR2RsAYg
u7kC5mnI6W+xvzOngOF9SpuVhVD1TYv8AgYFFJuzo4HZZnfSv4mMnhNGRmubEpbxQIBYRfGJKRiw
CRq05EpXO8Crn+LE3342VnN9f3z6TyWb4IUdX8BuCya783PO0I2XQlfmtiIUdpPZj2OkvldyQTNE
LYM51NlrjE46KozNcXRZJ+bRWjI+zkjdx7KfoOwnM7UFsl+VkSeMCOu1gEwKcAgyVbQ80mQvnD1X
RGw4mYdqIG91rcjmbww2gdlyPu85MNDYQruynm0qakPOLs2JMTwXoPLO6g30fLZqJGW+H1VYYCfU
FNAuxkOFc+Iw1Ip1FM0nmCe6hrdcvrysKEoaZKwXPfvZdmuI3RFa62Vfij8gbqtSosLXfT7SAXq4
6XhUiQ01oz4uOl4fdmXXEZyd6ZVznCGvh3zRFKXKx+iZJcAuxv/kFka1wuTfx/npH6O+EMjuT16a
PzlowF4iJf+pp3A8XY/4LMmpGJRW0sIAEgCHatlmIbpdbeozn0EkXlVqUoq3Qd9NSHkrlaPR9rlj
9MD9qryjVn4N0wO4EOhrKCmGuiormnqPgjcnKJvguB4Lxoyx0PzmQTpw0kQxGu0kTYX0CqIuLSG/
GOHebHGvvlDbXimbHpNhHvAWbpYtuKXIU6qspk2KzUtGzztUk91R+gZDQrm+SQJN7mpAI2FvwiRl
zWXbetvPzkeCemuR7hDQaCKPke9A6NofxA0HWS2LEMSRm36ZzA6hBtTke75U5Xj5jG8EhX1LqUzm
WYDPFa2c7GobKfmBsVdV0DhRZbNxWRMpYzx3XeoStW/Q0Ra5aWxiS85WvsJmdMEIbuIK4kokKb2+
A+u19D6xRXidsJzJHIoucZxerCcieyDUb4XeNZpujvulebBQgW9YsLiu77QZkDBL2l6G1LJWP/q4
N9zEWisNbPtRFrRPxr7L1R01HC5ulBxSbGiu097W74xtyWgL/AEcCkJXURl+zxknkUT44/of7+oc
BGbZWRSKPSgu3g6D2EhWJNzi+gUJUQBvP3hCpQUEaOs6oHwD4EcY/yFjiFMMYh/9XkNDb+PKCaS/
qnSW/C5GlUnWj3QtIqQeuu02+9AfONUnRxH8pc/HoYk7TcMsG/xEHjsKuuHFSoPWyaPS4SeWwTUe
kvlNXuh4tFDVejdfEqEDGH+22A0cFvFIQ4002z25eTQTkYJDskSVublaYYJGG9UiBAQYxa/2nvj1
81lTsnXCGAqx0nXsdTjO+1xXglyOisF4BT0kf4OBX5Qz2w9IKngKqkX+4eq1h8EllsAqBhLRQGQl
oQNKG589JoEK3vGp4Ga1w+eAjP7oAePQtqHp1tcxS71eQFiRyejV8qZ0tP0xf8TQRiSbbuEx9Ccd
TH5U+sbI+Ze62zY5ZRVG8Dpcsho7/nahHm8CLjf+h09CAw5YmFaofheKTZ1+bXpaht90bakLtpnx
BMnazwFfpPRH2nTQe2pbFpIp6mgsEiMkDFiDUNkNF3qQC4e1iiidU3KFOnGSMRI8nAFC9oyK3Gnb
v8cnKCsoTWnLiXYHFQrtflFmPxNvRJvW6XwieMnh13j2TIrkxZjdOu1BkVk0sc8h+DLk6zGnKF9c
K8M/Vjm/XKuDmxJR4wXelrHE1g6zv0yfIRGVYU5uz0cGEs78q7AV4jAWWvAG8KUe9+LIJRVq592/
xR56J3oQfOqxKVD5d0M7IVZBeXW+iLcg9QjwBl/Wj55fbA7O1Ykrzrc1yoDJ40lW2JjxFlaxBPzu
qDZoD+IkX3qt+E49jnceOg5UEiPZB+UeSmbwWm0CLIlFYjkWlCDwVaaNrrM3E4pbz2j+8LnuguAS
xD4ftr+NQPC40io/Jsq1PGhcV/Nh0OC/DIBVLxMikFTb7N9qfL6pxe9V2wpMeweQWr63OFLJ/YRi
ZZupMr2d9YxC/teu2+vpaEk1Ch42eZPY1JJ8D/kGzaJaQ8UvRtjwaJYPSZecQOWlSIUtvtXtbWQK
xToAeusLE1m2gF3fPVWwNRSZEstNlheuJQ4UUeg4S4hNVFQL9cwavL0AzDllrUYf+8sG+J+YFb5p
vcOq3Kd7Qx3ct8jwnsXqM/vot7xS3ADgCZG/gfA217PBcXSt+8h80x41hBX73dCbR0TKag5CklE9
U+gQk62Zmj7tE/vRsm4tprzlE92HHMtWr5Pt3hGR4qKbMnDy4Ua7Bc7Eo/ZjwsA4m7Dz9jocxcSO
vmTD2Hhx6H8AQ+CHI9kmmCdJWZ0WKXo6+sPSfc0jILo8l5DX4J5oFTU2LXHokdQCsNu7nWjfKbOj
DqySp4i3DrbOm3Z+vpo7l5FLgfF+TP5yVQ+eMmw/UDHyxpQLE7u+xWMKcRLcitgY5TIq8chiOkOH
VlGn3qsnAfkuNPDq5eYSObzT2/xfnQsLDJni/1dFB6AZpZmWPGeaSlMdvNtP7kkXDs9UAOs/38ZK
57W94KafEpzKqJC4sGxUq9JWfZUa/UHWy+KzuXXfuX0F7vgkbij0BhjDRfXpyrb6bCTGkzo+Jic9
9sfqxgRLTHbrbBbTXFab9mquskGyLxhVjOxJJqpk0csy0jIu0WxgfajPaH2SFwqnbZBXGdjUNAZW
bvlpuS1Ry9caTfDFuTQgvFRwrSzmmNg7/9ysiIYhiIUtWecLIwGcckBjNJQXDlo+W05P4W+xpUbW
9uqH38cRYeRRFJT9oeQXp2uaQ4Y8cMUjAwgzz3mDQOSdb4f2jf8YNKV1QUSKU8Rj2KfNX2AJ8uAL
bMFq3ELrmLhKUlF5yDh6UsrffrYdsrh07u+x976K9PPS77CSv6lBdvDyCxMpCdp4t+hy0o2weEHN
uGSPpUlPyjgbV5JHTyk5ifHyGCAOLf9UZSH+tpg/iwbskmZc7H0A+8G+ts25Vx1BVijFyt8Sjg6Z
0BR6JXeoKp9iuxdAOiYgGbeSMQRfRrErOypB1pKDtJEF04TEhvhiLarNCWwkGs0WWoxjAaGN5XQO
cgykZYm3UndANOgeu5R/O5BBXyJhpU0XXI6YFW1bfjbbiysyGzw9PbqfOiAFEvfjecvCsRdB4g9e
Ml0CFsuNn7SyB6GW5sZvmnDAWVsAUkCcIhKAdo/fTqcg34Nh3ugVAM8ioBJlemsSHFwNleG1A0nO
1MZ5vlHMdi8zp7FPEeh45BRZh4+94DeYoDJWurhOHNTEXPO0g10ZKrsq0mMZrMHQl2n9m3kAZDJl
f/SoOJBQdiCYGlFbx/KkyJjDTE9nPARj0L2cFiFQtcU8LNNAMHTEKNJ+4JyFmuhB7H+TY1wNGXqa
Xqho1q3CxMbYHYCq6gp2e9rTHdwBA1Myic8FGPkp/1b1B0TUxOnvqWeablsdm3vOEe69iJI9qdOV
t7/L3UDC+tc7ohULq6mfr81reQzH9MatCUlvc+HXL1gH/p7F8ueJZJHo3OhUMFayZlk9x/0nsu36
6s53LoeBZhKCeXdobhltv+H39UPUVV/etD1bJDxDL/jQ0cQa0y3sNGtVddUK77MuAzI9txgeynW/
DfEEvXDv53R+TcnyIE3kuvaS2+cE1iTWKMV+o2QXNro25n4d91FiyQHgy/66s/HwlmE/fHtLyLgk
iA2MoyPE7tw0M2Uxai7+TDGjffPzq0nMvPTWTFjkRbgQKYiiRWyIS6z+NYPi2yJX+qZCFPRUAqBB
OvxZpsXZYOFTdvefZZdJqg4bTM7tvy8xinoBZLruTD3oB2cQACeMLkFT7Zw98OEByvByN/Opsigt
ao7EEE6aLaMy1+NLGvfg9gYVcQswSJ1gqTvODEH9Cw6rNz2c53UeeCzZ788AB/0spfRieRVZH6F7
jOOpuj8ezUTvwJvIr59H3H1ceQf2zb2t6xc9Lg7emyVz4+8OwIxFxItiijzqPsnWVWCiigI/Whdz
H7EfaisYpyBpTXWGaIDX1dYYmNFMzOFzObd2OjCSniwYHTt3He0YiOmy868mf95p9iI0QaH154Wy
Uco/XJf1Go6bltHsQCLqpbAcGuRwAqSQVa7u1BuR4MlzkEA6DpN+Zwg67pwSvC+brYfhGIoS+vD7
lD5zz2kXHw2EHxOUWIeFxB9VIJZL7aVjHkeZS0STsFy+DSEljkB/FfZ3+k/zO1GTz+0lcL4xs5X2
2w/IVjfy9VVCPGflIH6a8psx27Nrpm6pGpzUMLaGjAIUpsmT4J9oZ60naakOrH8F6PXKcXLRg7kS
Y/8fAFu404Q7kPnwGXQQu7+SNGpo12QybPdV9MSIS2WrfApSSYrWHjZTBTlmnVkatl06nayUVtRM
6/HqFBWPjkdIWBi7r6WWKIAgcQ9Gea3wfJvA7rJ8vvLvHkSc3KfLdH1VEUqXBqaxu6yZ8S5VhIPV
/6N/YZy6l/1PEgr6jSOJ75/rrwsgxYnrhPTmfvbRcvAxHhH8kPUIEUUzVtWyk0EEr+r+JMCvI0Yd
GZyjvOadncKYhJXZmNL8F84J5vZQk265pfDFW/gqdi2cVtp0fH/SIp1aiT65rnSZBy/NNwedkyx/
lHyHCGV0q1FDaU9RLE/abmFQfnMAcGCIuo5VxTsscuDenwN0JTQiIxhAWNVn0CQxQOYV2adGev5j
HKsWB+obxaSWXId6DuNNfDVPRYy2ikUnBHyjy0Kx+fmXOUYoYiM7AnVyEGI9z0Zflp02YlqtykMj
QjLVQDoq3X1jR1ihDf0Q6xvCZ2WFXh21qVe3NTgk6pprF0BHdEJBzdKBiWLESnueb/09AzttVTws
0432aVxE7pl0XB7n8Ti5K9edguVXmTr47zJsz8LODFpisY7kJuZVZ3Of8DU7NUL374k4WMNpZ/8O
LH/vKqNahZczbNMQSauCZ3oZQlBY2OseKHdXolQ98b+Kxi8y20zCtOaVXJRW0MieXyg9pW3KPaRH
hvCAbq3klukQeO64A+BMbZxVgF3pP5hWM+hG85OY3pm5+DpVhXHcvkj7YIyl/vQ7x3rbG57qMuad
HQIsBg/OowxkCe60x92wbmFHtWSlTYoKiQ3YnM4DuEFijk1ukwug+t3ExbZklgvpAYt+XSWCfIbz
4bkrcmfuRy+8dzlodiS/pLMtu04sAXUTwrk1gPTBUGlOq6GzUWiq7bICCwZfdUUaFbShmeCM1t6D
mlBpS31zpYoJoDboLPU4b1xSba6/a4okIuwh2k2QsGmWbU6gkQjAyfnA5vicoyvsO6uAXgGTlkH2
alUStcrGLYre6Q9Vv3RS4RpSh3cmV4PFzPB9OTR3Jm11t0Tvemyz6duGepUtb4p/IBNFc9WqX2E5
uNm2qc4mkxrF7R2gqwcxv/72h51G8yhYD8h7D0yfiFRkoqIlfv+y5lwbtNaCEIC+mcuO+Sq1+iZy
KKrlIEbvteDdJ4KR43tcsTwdEX6etF7XqoyQTBHcOP4/seQpQ7yutheWaT/7671JbaDmMWtzAuul
oLVNaKehSGzoScva4/HkfRLf3hkXOghuBxv6ttgsDIyM7BIs+XcQmPQX+Rjamczk1a6IPwg4Cl/y
Qm45qbkhAc626L7WPKm9PKWPQTWNClFlSQRQTvxglvcbnGA1hFd8wxlUetw7G5oLl2f4SJ8/+BQR
iMI3WDr9D3ZWy3AKvJ8GYwhEByrrBcsePNYPeY4PO2IId55fQLHkZFWFuMbj7x/4s6ERUxLzx1zG
PIMmA7HcdED/C7A1p+HX7RInh4D64P9l2cYEby2IQoMLaTRBvbuCXzBTsqcIZg6xFQE+xfIreuhY
6Q6iRS75ckHbfezn+QEBTGdvjQt9nV0Kg103sfnWfL230qhR6DDNTRWSDGwiZtn4jNttVXsP5fuo
zERBLkIwet1qQk6KeK0/e0IJ0SajsS40snxmRF+6RaC9A+/piLz/7qB+IXZaZO5UpwHpzkee83yK
rP0l4LyyI2AgJLVz1pjZLk5EHv/rJg5AiSkDwm9c5imM/vKw32wssRC13sMd8dpka12qMxrO3YYY
Veb8NdSFR68dAoPTeuYyWjic4/iGbf4x/d5aybOeHbt7J7KFZTqt6YEBAMPH254v81YEdcoSe3Ia
JJlpVBKB2SkKN+9LZrJwprt63NL1zc5TdEJ2FOTbCopnwKrHV1CBD8vjRMU2FxbImelzin0YVBFQ
z2poZUq75dcq1FEeAxIjA5q42Kz2/eOHE2mvDNLrx4eTf2dPi3vSkDb7DxzS9dwTyYnxzenuBTu1
ZjU58SWIbcAKvjGsrjyZSUXfyGgjBAi5spX2ocAbU8DKw3NP0FrMGB9NO+Qi6Klv7OIiWp5Na31C
aDA6VA8d9xm7WUUbW6Kgq0jqhe17ySAPdrkSDz3uV59do4aeJ5Jro2rUX2d4F+0M4H/f2JowUpZR
/LbW0WRmZpMY8R+X2joC41MZtD34VR38mJEYgEm3EwjMMG2bs7WFK5vXRlupIwD8CrKRiapi1/YI
ifePRCte2s8EngzVqyBTLAR0WJgMgJchEtXfnQrPpyufRF+7gAb1xW+QVIoFniCTqR1Id0mSbYMj
Zti3i9vjKeVHYHDI69/UtvOYFkpQlrrHiyaH0cV+rurB6dqUYOTeBDNYO/wXqyywV7rCnKsIp11y
FO7AxYG/BEosZOINGd+pbHzMBfMyJSKpRLjfE2QoQ1tSbQZ81FlxQN4NnIQ9YPsiePBATP5XMwYi
yJ7VV+PFNdPCnb5siSUyllGfBI530n/MdU9o5ymdgjiBmM2a0r3gOIj4p6jlhouSPqG4T4CoZ+12
Vz3AarsMkflxYUGIcOurZjSgA5sri8BC4+kSKGCSF+57goMKYPCe4V5hd5Nj16hzemz8jngY+Uak
vH6kSLBJ7JgHlyiFp709KRC5GoVn2m9+hwg=
`protect end_protected
