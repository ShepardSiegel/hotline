`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fipyxXBj1iumYrMxFt/PKn80JAuqnTEBENk4afcOddEctjojUhoEt3iZr8sZK4IEoJ0cF/X1fjZ5
6KxpooS1GA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
INQ15xxT/xfMzRAsHSwCd/MTQ2Pv/t/xfVcsGTcoiqq4Pj39XPy8wIECGmoA727ViMvmsJ0edCQY
t+ZHq41/4q6rlmgJ1SfkgrWdvV0tBBhuWwt00Re1Sc0BnR6Q+qrUF/fj3trnu/pHPy2ZG5RGkD4W
wsHiJfruinWuCDNp0rM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NYHy05x+/QfVkCKOkCKLjToEjJcxtba+wf8auULf4255yAOLzEQm26LYANQOedOetKoKSuR20TeR
a0E6XBueqaK9oXGibfbFcLGPUrWrw9Sov3TslMFscrmS/yHXwzA7T12fl7oOBGZfEly6ipMhL0hN
kUwwwgK4cXQSVy3ZWSQivVJG3lABrQxayQFOfTZR058egsRDKIebrVEIzg3G595SikExyS1LlTxA
O+Bp7bzbmq1eG6jo3zy/U702yoFTX98Y2Omhv/QJTpKAo1Vqovlz2bwxFRGkhj2/c7TPfRGfkRvi
c1gd/CJdrcyG75bXDm1VwG8OpBtiO8LhPk0zbw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
M3HO9oasC3vnBkQM11WA6wMWQJJaaSV1YAzRflW2FBHAMWc1mX1l3usmNpOjCdcQzEiIXDsdebMc
NDRBqrXYp6aVytlyrC8DF0H6uvGjBR4fkC8LTqtU7orSBzF1uDWxt5syaf3ZdheP4qUiyuWYs454
WdqT6doljGP+bBLjr8c=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZA4r/i4brfoNvNtGzBuCpGPAvgRIlp8qCC2uWyo3/Obr9z+HTAAJ/iXSt0ISlgifamQGroNZ00ur
zuOm26/yMJz2SFibQgCR9orM3juJdz2+HUaXe8KADbghMpUvrz+r4rdOxlXbA1B4ThsVnGru/Ee1
KbFNjV45mI2PWozPSVZPxC32kndvukGVBYL3v24JsrY2RIn1cY9C3ACXgwOhbCNi9uKP0trhq6in
/vm+qmsH50EcEKLAJaE53gztjvfyU7roV0Wh4jl+ybNzua8HxZcE8pxWFnbzSq6pVn3DQRmiksjk
eHCsjbv9cIjXCrCGcTN0r9zge3EvU1UBih0CRw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12256)
`protect data_block
EAmLsU4JQj2Rf30/YTdWwtu2PVYgBOGrGboJt1sICelApNqMQKv8yAdfljNxdh+ikIv1Iu8dtPKv
ZTm5KkY+iVdBHJJ4o4BBGrZ/vWtF13nt6Z9JQxHVpA2eh/j9BttRubcFc5vYF3B81F3t8hndIkh7
jcPHcKxphzQvgwzyHZlAKce+ebaIKYAArzJISYPTuF3ixROTGDbqBPCHqY/GV46rraFjYS6wvs1w
ec/U57rKVuqgBda9WlqNJfEhx8w/ClPq4cfLOquS7TaS1V2+YeV6IYtvJgG0SLkJjtC+tIRPmypi
Vq+q+X0yaivfpgsepcSBOGon2blBnWTc3P2dqTASqNEHmD6Sa5G7oFpU2LYcCuqSwe+Cva/WjILq
IzAJp72MYE04VPtqzw5kPRVOCELwFwZ3K33axVo2Z9d0fPkODSemGuQ+BbDnwuj2cBNaCI0SrNAt
D4yGcZ9770orkdFLOt5rwiKnPBv57R15r7bmDuKSH4VtCfx7fCzppe+ImGSW+8qCiYFwXCrN90CI
LV8LpZbO96KQ0UMUkAAa8NlxVl0Hqk+8YGAZC7Kn9Xt+T5RHd0/9RCvxSSfXD1DEv1gxp0IytnE7
Q26pEyEDxsVGVv5FC613y9begOZNVePSoN4ZqqeSh+jok7LLOyiaPpYzcajq5P0qMTQyToKjxSrH
S3FFPyGBoTvR+nM6NfRGSF1VyGHblWvJGX1FumN0/4PRbwUSuZfu+sSXxuhkqHDK/h0pcqLUmz8x
Qwkcl2nYBtlTAKk+cBjVt0VWjQaZMp0/V3KB6gnJKY2k+SYWtx2z4ZeUg3KilgRze3j3+z3+AuuO
GKlubMb3nbQ4V1JIIhLnMl+TIvN0kwIVzAtap5BSPDWESgT9+Cdmlfqx9AxXpW0scfPchHxGuGRo
Kaqi2gKHkKM7HY5ytuxtkYOz8KoFPm59C+BFAavsjCwQq/aFh8frTimRg7PY+mueh2wXvcSuzySm
OVYcVMpXODFR5nO3bx5buCTSK8ozdPCvfg+LbhvhgyXBC+g/uAlNXt6lxjB/tAjc2P1NBQ1hTdCU
8MU3rcrfKiy35oYBlvF2IfR3qEa7cwUl5FhwkbcPZ6IxTHyhMSgS/sZiksR3hz98xguTrE1NADCj
4nfzlChaEOfrbD3Q099eqPx/ni09vwM2j6dr/r5rE2YOC9AmIl2o//ZYHVUxCwLIk0KXLdWcylLz
sg3QbLDle1o5sgP6SohnDkCv+mfIK3/nH8laxH2PvpCmqVRO+qSCNkpQYTr5MipAu3aPmlnnN9IO
uBZizCXGddt2L89Zbt+1ARbulE76y+OZoG7I3CAm7vNtWWGD7qbyNBHyd4B1/qxI8GonPZ2kUHax
OjQ9cFf8YHGlX3uDdkZZS277MMt0xEqYx5hSSBTrOlHo1UEWJlgxPNXhJRUOHf1HjgrEpq2qfe8u
kAw5pnDY9eVaEGzBxCMewL87Yjl3CKFdsVhwSOL5s7eIu6kjuBQA21lS7V31iiLBfWkWxl6+ag+V
SNlOD08a5vGuqDu3bOkeg/0hGGXlHB4Q3IEmSOQtiYv1O5JbWIiOqH1FmEaMyvNiM73J9PItL24m
50aygAHtiH9o/BBtH/MA13k/7tanOUqRrWL/tMgldB1dsTvfScs+WjpnOn22byJiBKIgxgJcJzdS
tsrXykd4VlTcCRqlD2dXhmFNc0VKXGTFFMhTAH2Tr1dGmZSf0aHb18oD/rUXnuskx6k1ZjBrALil
LYn3unw2Dyl+BhbJBuAnfcILNTHGNNO6yw91BmGwvXHEsYZaBIUQqGExkoUM8zVkQcKWnWPEVHeg
7102W7EnJUP9Xsp5c0sQQRx1xWVcDEwo81gYZTP00aK6ZMiJaRlYJu0bM9QGlUz0jplqd/RFupJp
A8rhIUgAAyF8kB9CrSHFKr27CL19W1AO2zhLBEXMvFE1CcAWcZKeF7r0zRMI6xig5s1hJPAtncyP
W2nDofCw2AJHgH9gms5ZQXreQ6VinMSKN7sit2cUJlZ83QPNDc1W84EnRi3zIyoNggNfLYYmL5KU
Xk8Jbr6cxHakNv1CYgpKbeGSZxJmHUQQL/Yp5GL/hI5Vy73lDAUxHV8TbFHwclB+24GmlfErdGrI
2g2ITfPgxkC0+vmIPNqIDikBW63UmA4k4HQKl0Rq03LJnJ1ZyFK9d8upd91gV6ShQ5OW2GiSLmbo
QEXhUZkFCde9QszmGkSNMWNmrZtk0VfxMRnuKk2SYn2SlcMNqfRW/CMGyv7rg0hpJjGYh4yVHOuu
rd6yxZ1UXniUrBLY9hEVGMUbvHKtfbxVq4r+6k4mFQOdjlfA3Qj7p8XScBLZQcYQCfge8L6+XBL4
6FGeeBY0EEDYy55Qx7m87qNM9tzqVSOlBHDvNiK7VJ//4LmdgDSM6oAN+8HYhObRenWKzZUdaPwA
q6dxtnYW0Y6iA1/XS+gdHdonnl7soujJTKqerHYqqXNM4eUgM3bgE7VrPb6q5nA0rlO+AxlEZWXi
tyUZ6JQt4XyG2VyBurCquKt3DX98yxuTMD6m5fZRczrfCJWXVDMM3ekhXh20gzjcdb8RM23VhapI
pivN2UAmnaI4nXxJBopSxoa7J5xxbCZgJnPfiC15OoA/LB7gu0mz07EaMAALftUfSGBQH1sTYIgC
RIzhygmEykkCG7y9RWxVXh1h+eS6gU8n8w43FkS7wmM06OTpITX6Y3Yql2Y1qDv+A2MzSp60ByBq
LjNqCjXK4hbPTm+KX4QkBuFRUhPjgB5PBKFSFjNhwyqUDS31PFlt/KC0kud+/vMjn1IxCo9URyaH
zpiUdzcm+A0KSZX0f1xulYbryMCOs5iMEPrPA/fIDJzMGNYjAdIRvA0oAaoNKSOEf1W2kj9ENlBR
TA30yHoLJXCCBTAH0vTv+xA6rlxAvJxoJ/ZKWshrrpFvcH93NQc59KjbTneCia6q8lyzHfhRXMpI
G0sJwoN4Nd81kRGiMG36vk+/ItpeajWm9dM/oUtS44S9eEXC1Y+3Z1us4MK/Yf2+nlIQsw/NNpbt
l49lBrJGpzQFea87pcd0OpYSirkVPhEawL0aO9Ak7Qu1EV/YmAQdwxaQDwc2V5nG3xEHsKk9i8OF
HmIvLJzu9t/k1ANm49/EMYOvYDjr+1DF3ugd5KuiOQhupGBvM+UUHc+pa5X3ag/a0XeJm0LQAB6h
bXzAIWWEFLxUOv4EQuEhoaGvNDVSl1JpUsvGuavAF3Q9Wk9yF29Id+6kLmgGLzNmypsucrIg6a2O
zKi6ywMURXBrmjKIMwjQNja37kG5rCNhrZ6+be6T1RmKKcIY0PtVmMppPyW75NFhcLlO/IBxdQQO
Bejn8AKRAchKkEC8TTfeuIcHq+T82LDkBt8xtp7y5pkT1X5UUamMOnDbm5r92VL7ScJJsWRMdR2k
wlu26tIwS2iKHsSjucAeRvjfCRTmK6Q/ZDACBC9tF3op98uwycrw7WGDRwLvfoZXSOFmiOgeYdW7
1khlrVS33GWj1O1d85fcamUDnX60wAtZkFw4lvo8v0mY0Oaj3/90FzKTcZdQCQhDq5Cki61sQBu9
/ePRK+bDo/K/xp4ACR29KJz8LJcj3AsO9ftsZOtpiszb0lsvEG3DL/adE4YKfdvvuSrA7bGZsYhH
jNjtpDEiVWJaxtvEJzKwdPqvHy9cttnq++4relCOqcuxUggr/9PCKM7PU9zhfPD0LOlqnhWpNxJz
dykRUZXT2CIk4m1JxbLljXxZM7C64EIzqju1UwDh45frqzFy4VL0r5gcJMYlPzp9kAgAfr00XZGE
w3tn9xdTnQ+l2ucxOy5XqxOrxQkY0D4j0D8iQLRK8HOUzC2+u9hVLz4nfcMjCYxpUX9blc6ezbgE
rVMYFW259Xwue+gnGeoKtFqgNFAoIV6+U14HMvcFFpRVuReqDk9m4o6BhGNihmcWOe44tD6l8ede
BnqWplp2eoJP4tT6NHZ6rGCXnkeBv5aeF4UoUaMcpH+gSXBTC05/AgFr7FgY0TNgZvvbT3EQ2cvY
G7GPDb2v7S7KiB/nQyTjAGk1wHz29jXNMrI/1UufrLpXdErnJrTusdACkcVb+kZuvF+3hLEihYxM
OGitpSQ/bbYYi8IE+ZgusuKH4R/iOH0oAvYRjODTBjqFK29aVNDYiCSIpv5C0B0rJuBy/7vMf2ph
3Xbqc17QdL/3kzp/peepnZTRfVr60fFHPQchsNi/V+sCJbzfFde0JRmxHi4AUal0AG4+ebaXxffq
tkiYqTpHfKxAObbOlLANqxnG/2SaWIoBqeIwt0133RbGMEcfU7zFiR9cvBcEj0SZxLj0MkLnN4Ql
sbFCr8o0anMkRlU8kTUpML9FxNRPKXwBBM553v0SNkO2Dt//+3IJ8nNW+cB2PoSbUpzWEocsfneg
La7j/kBymEdNxU+s70agflcXHqwXQuEhpazBHuQQA5F3h68RtON9Wa/IoS3zREQfmP3Qlc4sb9Qy
Orr5Kg6XHBYR1PEOGM3z7Tcc/g1USdigEVJNbMUdImwc0UBjcmNQtQcu9DSJiPBwXXhJq3RdFYkQ
nxFjaktRusKnnbjthbXfDYxfUAOaNODl+K6PFrV2fvO0RPGKpXgZmHZ2Xo11KnwCkebI8G7mR43Q
zPaeQi8eI2sUnzSyafa2+lFdFKLrHcpgxn1iVe6XPb6F9JNHJjUqfR1Sl8sGgKCfUum08eJZ7Y8z
nqeK9c+koB7kV1tNgngi9mgj13CPdPVp3O8tOeLDoZLFtCtI0eE4FoyJV2h2yztuUSJ+52OulMkV
H282IPnMSWZ5c6BJl4d5JHqzgDD//qxrrjQ7P5a2wEUqxQgoDDoqBwHLLIiJRkIXUYlu7DhG9KNZ
A1LhPLCgCj7kArTLN9GQ3QhkZdS2EI3Rye2i0dClhY2yX4oxgZ0njYhRbOCB6TtT3lWZQpkKC1X9
EP5+qsZ4fdl2aKXVEA/seyn/JuqKilbxgTl43jVtph8uG/UTS23O66Knw7ufcwqKnlzojWUModZi
uExJmB25Ck9+VzNaDe0DrUmBbyYZOXhpkCP6hSFNmg4Eh5R0u/tt9dQVuve4jzGcv0n3IOEuvrc5
BhiTdLjyDw1JYaspa5K17DLrtElIo5QYNyEo1jLWBTbpCHUaw1GS9Ko0Zgrny4v3x8J5A+7f8Apb
BWSsyS3cP73M+P1V54TBbkmshYsYdCttRn1OtaDVOZyzcss6BWshwRo0hAdPxfsMvlIFHNJnj6ET
WQqt6tpeV2LkXYiFv98ah/Shj+0BUopyObQ22CzHjESq2JzzlH3cXx7zriuaMyAAM0+6dp9iOTOq
gU74NNeb24QTeQR1PDhYUxDnNOhx0FoYMfjtDQ/zEf5BPSzWbJsigjsQkZbwRFXrdZ/Ydq66nYQP
NSvNfkPkSwWF5OokfQNSTNUWzCY3FTh7n5avnb8zUMkcWSu6itD8/wZT35+NikNL7pOrA+wSQljz
dUHFjn3R9jtzApeakW4DR2Xfo5b0JjaLhGmaizL/vOkele72sbECuN2Cu5D9iwU7i8Pi+N5jag+Y
tWhPDLecHlEnIGGQuo6GiwvGE03rSIbG11N+9l0I8+AQyv07hMImXy/ll410it+ncJDGFCx90VXe
XVnFde9xOIh54wrBjd6XRZ9kU4me5yG8EAHdfVwOppmpga3BfUdRAFwGxgMnYL41lz+lYo5cetWe
UcYUTY+AVqoxu8PldJL/+UY/4z10f5WIy10dvm3n9u1PoKy2TuxABnfgEuMcC/KTqtpCE2R0h2eh
w6UHYtpz00rT88yi29OGtSA1QLYEwxuPxXHIFAY3d0i6lTWug/Df1SJx+02ZYM3sKlL8oGwK80O8
sBumOxKbDPqMQB2SzHZwh2AMprN5xboobkHCOwkTYD2uj/YNfDzJ/xcMhgznyBrU52jmO28pJDU3
DDkInZ3f2SMPJhxQljmpB3JqMT1+Xz/8EwIDYTcqbL5gBh/xoDj6NMy9Qnf3qhpID+nszZDfWkFR
tQznNT9j173JOd8kMGpIlWMXhi3V1jAvVm9wIhaTxCGvncaOYAwBLs3BVReB/oAJ6WOx228LZORe
sJQnuzdr+JpsuX3530YBuaDb8YC68KEWRFEplflDolr94ePI0TmIK5N2seBEC5FPuI/4GG4qwEQz
bzOIJRuZo2iXU6vbvXAmexCh6FcIk4neh39gCYo2dmxwzJ9xVpYogFJ4qGua2X3hDiBx75AVUTQW
Npb2Ys1OehwoDFaC2UT2HI+fNXsBTGVeu8Y5xNRMmQBbABkoX+1G1kwBFoO6ewlQ3T4jrYa4P3FV
GPAsuBDSCSgbO+HQNAV6IRmP5tSGM5LNFr94XXdichAHhUBsTNwMMyzFCKE+RvuPY6IW7CBzn4Xa
NxtPKhKG0vEPotwwvgyoQTrYSQXPJwgjf3l3GSDn+jKpslUBAY5Bft5dMkfUwAMwStc7KSxxMoWL
W5W4vh5UeW5xgO9DGHpsHh5/ZBo+50Qk3yYP2R8P5ZYq393yIQzjiz98tbTb1IWYQdiGY1K5Wi9O
hXU86F+zBjOLD/8Ytks0ODojeag2QhpzXhTk3lxSFHK2U5xlKyHiHmMwHm3+SCgv6JgmzxtyvBDE
6jM1o0OZYSy/kDKxveppfYgVKhObKQUUTJRkXxGyximlSBBZ7YzFIvXLAgdbLDXQ5TQ4COJ5IxY0
uOCqatOiWgBp9V+c5VoUJfKoDt+g5utsWwXNBdBMeXsEylAbAgwcfu17/mjKIHRNuXCLW3+mheVu
+GN92iyCi//ywo26aXOHfLuEwDOV+h74IL6XT1fwalplfNuA/LlCDcWCNy04/B+imYlbSn8rsnhi
8dxBEQ/xEJ5l2ql54CnyXXypZCmM9/Q5xZIXC0fTC0SatZnst+B6J69FBVW/PBRQAKNuu1jWZ8jL
EvummMyZNJTp/YERsdNAs8j16AmS2eNG/y+yq1/PjmqIfyAJ8C0L7aKGQo3RcC45zBS1qUrGLRZ1
PNLfXB6a56xpNjdtLn4SSMS8ocxtJGS8KxMPJjjqwJXszHrVgVqhXQtndq6wMccMgVtUOY8bBvxZ
cpdspib5ysG3NnN4XZCDFg0YWHZjb9v422S95GrngyEI7byHViBhWm4JcFdBOZ+7+2cOfLrj/kMe
eIzrkG5DHmqUkrNvsdWFnLg/jfakd3W1aKlbkfufohZ0to3g0rWXY1OjL24GnhSkES4mW3O8Xo8D
CC7clyKxg6r9F2BVtlrbKitS3krPmgwN98p59P7BRtoiRzvfluVew+qqDmfB1rcS05OMhK9qJhuQ
ag53gQXUIm7Y+ilY5mrUhJ88TW+zbbZv+NMrKdFOZ2iwMJXsEsOfpi30RCvRPGdCzJQfmrnDl73R
sls74HInzxUKGGr5thImo6e8PiUodfX1NBn5w3CLetEDGA2jnfScSXvwMPGThuYl+XjtKsRTm6i/
dRkmPJ+fLA1oVIJ8Ny1uW7PgZznyErHCZHhFfhjOXmvy5n4dfydGqaJs4dKfOEudUn4ejsz0E/VI
+q8RuFH8hr/b6uxptVJfBQlv2XeUpWqU9xAEZUVqdmHMWKVXExezQJpQRa+HvO3OYKxf9NTw1zZY
eslPa49YGulv0mmznzieyY1+d0EZhLxQ6Enl3h7aX4arPBaUYEhLhCjLNlTUeLfpXndpTDpTQf+P
Ywj2ujfMpfG7fUXSqMGp6qViUFsbBrSZqr+Fp8EbYc6krhSaxbEdcIOHeSi5mcSmng7erHqQo6ZT
buV3zcltoSlKi0aHPpN9oHTOUp9v3pPKfCXJlqWKuI3ksoZnvPuNFqwbVW/2c3db631KiR0MIPes
dH6HoBYW5mGe8KKcXNZwpdQwFbbQPhwWIF2w38Wr3uZDHKWVcSHYVsHLslUDLVNr2CVqYz/xp2Yz
W+21/6on+UqN7zZLwbj3/dBzZKmSLwhz3XBri7dMAoFsdORBArDd7eBB2I1yt7uu7NwY2kXt1HOM
yMf3LZTmGyv5wYrbkzSUDjc5Du0B4x44NMqCWgt2L/nFJHoWIvrwXoOcMKbU1gsc+rDDGx6zZ7JI
W5rFE5QQcSm+aIRIe0ZQglH7uugSY2ZHLk0/bJIarV+5gbQEy8//I6Tu7DRM0bcgVJoZcVXL+lDS
+mFQebXXmfDkjKLfQX01wKMVHocfvi9g0kRg/h4qoTtX9BKTs0hxpNh7dYXtsUl5oAcjlhQbojDj
XEXB8T3+aoMqDtieNipwUmeElrH8FccXXDxY40fFj+lcKMMcJ6Gh6x0uDugbqPKnHCs0/bbYO2tw
XGEQMn8oGabBqM7g9JTIEQbywbA/SwHQKtQcaOeffPSI1jVx7mTMWR+NOuaX5yyFImS5wxViSj3d
L8TJrxI+5U72M8G1bQCWWki91IIkBHT6iINggYvfjjxRB01MvlPm8X5Mf2cMw/5GH73mBJCMbzpj
6Z7w0RaSt+0nE2fTnamBuxnjcia/L+DED6wB4gUfiVKZhLPVT+fayHuJ4dUxjNERmL9hSxnUwTFN
aFWIkNHbFzFOB1B55WJgC5quI6U9VRgz+yN+EzdRkwNjfX2KODvGNRxaV0qWNyirhoxm2DNOuTgx
+2IANcVscWn+917XjHVQ+i///FdcIoevIT1kv4BmixaAyi40dtiEJQcHvP8k1cVDwaH0zauJ3hGU
sUq9HrPHwR+ujXJJg10pFLXwJ3tytdeoKDTBn6oo/wGTliVYCOx7Gf9KZN9h9ZIvgd0Bp7frtjsg
cpa7/6ylIQXDMPoiKAF56a8iYwWVA5IZ7vTpDMQIa8YJuYMGi/mTdgRPACo7SmGKl3S5jDnCq4vz
CDpXrqcCIm/cnTfh2vrGCEa98Udl/nMfrHmTQXZ4o2hFyXgarou9jBJn6ls3gdiBqOvmDhDJlyiV
4Xyirc/0YbrsyiYWgUveOuI2MRqFx38Uv/MArXM+6f+Jqc/ELjuPr/gCy7eRH8yaox5esxgfdyZ3
LatgesLlUEg4cSPvk4redNR9gB0V0TU62XbcB2YxJD2m/T4vlzFH1ia5p0uyh/Qihf11gPsm9Z2b
xycm/e6YtG6Hs8vZe6L99cRjk83YVjDyHJWOr4pe2Fr6NyIJePgOByZDZhoTxqRLY4lLCRqhDXgD
muPXXVQ78k1x4UYTdLbW6V8dsXhcu2rosAC3NYx0rLE+oaobNWOusVppQD5rpEtG0SZhiverGJ3x
m9SKiUvrDXcR85k20yF/Z67v/3YRFgm5l7Hsyb3GZI+oKKqVdk/DtikgsAFKAt+l3eYJ7hnmt78N
U+99cR/vSeB638AAgeIdxA50HxbUAHxOa6tL/NwssyAGQME4C15mswiDbzsG4zcjjBqTrRED8LJQ
pJsmGPudjVoNKEvIlOdVqKSvIGG+TbDhFCOiFHKmS8ZYNAkOygVOypB1KHsgvAJa//m9uyw3qx+5
E7Ai9kNFZGQnebDuZzkPSfmQ4TOiguUO91nJjFQwMFuK5I+RqEwNvbS05nLA0shEW11K4p1MHXLg
qDfTGBWo0ZQQvV74qch4D78800q/wlw0fm4P7gkowWmJe6uLsuLnqvVN7+f+jpdBwJ71eomfSkvd
bN5FIwgf4zUOMdJShoWKDV/OOXyt4QZrKfSCy+c+HZ+n3DS9G/vFrC3dr2TdSMuU2UViPpAGWczT
bBQX9ikGLC0udExer2aOxBbxkKLYrcLtzLG6BsXj1CJW82A135jvPLU0RDvEl4WerdKVK2r9/48v
0OQU0nDVQg+8yDI57uXV26quQ3FzcW+jbRRArVqs/JsAimmat+5POzI4fhbDn23F2aZwQsShQKx8
DZ4mGQSGNQ8e4f80XpdWqruON2dbuK1F6tlMFbVQ8IucGm1M6bqz31Qh1uRdpvpVosIuGrusuDGc
VZOA+y+EGDZSgnOopI1A5Kzd4hAz9mZD+YAROeWzABL2nb24HxPkLoo7KfSOgSd+DtqW5pQLTpoy
WdbSe+kUFViI3sJDYuQzxrpuyP3RXwkSsBM1xvKA79ajtKdT6hd41/REpGrYXOnVNm2i0zeWnHB9
rKoS3ucoVDwEne4/ov7rXjiVcvXU59uqJwMKe7oS8Oshf1Ktyi7xBOSR8DswLZ+GhDKk26FhSBt1
4Z2/7R585XPU3khUnwAcfscDEjEadPMZKemBk+WuhGN4U6iW7DYrkeqv3HKP9Y5Y4NvCZRdwli1O
FgB0R7h0havuZn4A4o2pm3z/cdShW7elJhHp7cAsYM421+rBFMNrpcH5kQxGxHMymKftKeLlfeds
mm4ghzVAzS46slomE/2uboiP/WrILnFuiuQFLPxxdq1gYC4oyWor/5C05JIw3ApJbZ/YKDkUVEEg
lgjxZenA6FJwkZxAhk1pvzzu1SDthL2jWHcf8deP46xiFEIibFAAwDrj57lITSX6rLP1khh4KPuY
vwFRsw8q5F1kVR9avp8deu2ozAqlFiwQ4XFyMlo2NAlp2chYBDMzW44MkeO8ltNu9skzTZb6/cPX
j+1vHQYNJs6Mjm1Zagu8suAHoAhvLNmfVK7kctrJ+kGnMdEJjn7lxi8Y0nWodRJ1ccvIIVtzYZKV
HC6UMvoNofW0ytVAcS6ROH2ccf8BbKM50WgRtNwdNEQlq+PIbbd60xXxkCcteLGNKlxDTyFPgxzi
xqPeZNBB/TKNlk9P1AWRKwxI4nYYr/FUGnZrUrRZ02CF0JgggiXjMRVDTsAi7XCqdwI35G3YN7K8
3LzHYm7OTVQ/eqqVfJwkVEIIqbGaG1vc82JRTh5cwREtOu/1uJoB9gdpGEF4UnREk/p1fePxzeVC
/pI+xCvRjp6kVYx1eBffYR79UbSJF1xsl2HCB97W5VTj1g4BN4kb56ZlXfRNwUxYu0Te6xPbq2PI
v/gQNpcv5nSDz9u4ASjhoucU3mASz0kJEPPnEY+9HOO68AUTgimfAyYADmJPGYFy816wlNPgVOPi
LwISQYjfTESTaI4q2+ccuK/Pw/hSUSMHARCDodvK7ntmhiVbWD/ZzxbNqDXc+EvjF7TTQk8Y+6wV
7r4vt8aaBtrotujE+/XDn3zyWepHW69d6idkbLk+gerHl7/SjxQqJnoWL3EUlUR/N50aFd56vML5
G2IOMTWmTAmxeCkhSI/HZMoVbugYb1fNvpdZVHfXQbf2puTzaiUYUtDqbnqR3N3J2qZskaMM1PqX
tTba29cwqqLvKVCHy8utz9EEXgjLOVWRdEtNVezsw32vhfd3uJEsEnpJ88l0h3FiDUVNyoqvd5rb
18yHeRNVuhQs8aPL3ZttyFK6YFtMgJY/jUIoD4+FBs3AqnSrAQC/IVjww+eKVVgMEwrMRXaEMbeG
u6G65qYLY+zN1Etkpbrvyli55nrMadguuJWRrmk5bb3FAUMHNVXWGGNPz567/xSZSQh2YGFG42BG
kqJyTpdL5dvvrG7rj2tpv0oHcfZtQRiDNl40ctNU1effY2KwB9LqqrdunnXaYqLhLhEZJ2AwOyeA
xnZda0ruy2vltAt5MEGSspbVp+a1/jjMKRA59EM4sQvaIy+ZHqZkZIpdrPuOLnzNYxiLEf3ZBK54
UMFiknQc5ulM+w8gRh9yWNWcZgNKpCyHCTef7m6OUa2R0mTppMUr0eyLbe5NBcrSyOqHg0RDsIG0
NSsumxrCnIULTxYAESdKStpkx0i/Tvm9RcFTeTWHh+md9Ols7r0LQD+eJGpQmjnwIw5keFTMoyap
vo3du8WvYsfBJraqY0RhzJaXwMkaL3AB1e/4YTIVPjQbgrGNpSb3kPnylCgv7pZlPVJLGKW/fMw/
RSWYasIL/AFqv3s3OVekicdTov6shBL8MXx4RQ94hrQKQ9cOEQNcKuYa65blMAY2ylQH/peEmFzr
eG4ZGKyS0hJm6Fqpo2meVgXkrS/3pgMDGGxk6ETM48Ne7ssWUAMwpec647BPJCbIzcxmuAP9MpFp
PivXZbuFGrg1E4kyUpHzASpyXw5rPdw7tMhY++uXmIvqofVSvMsbeSa7Wn7ktDlFDvMbEqYnlZYp
bM5gY2l8jaeL7LzMkULblib/EQEbk0W6xDoiwOHZnQwH6l9hgEJESmjy+R4NtUNABhDC8f4VWuYe
wR86gsfHd3pU69PXTLS15l3ckLWE1WH8IC9A3qJOIGeklXzUHGKHYGvbM2jNOXe9771lFEdQOIFH
OEW1eV3egweb7zTHpEK/t3z0nQBouqewXvKhlu3VG/9l0oNfoI03URYsp4tD+9czL+QRK0NctCMY
2jdWQiZOQbOvixuuYbp4Yxyu2zW6Yg1OWwu6MAihzKy7CcFr2rT3h4fqS0tN7N46dBjmHDfvG3+G
d1bBhqqE+lEGypmF4ad0RmzHqvt3AMWsoajsLesvh1JcF8Sm2InnASzAmMkPLeV+RXW3wwxwsDSj
52mYjg2YdGoTjprUgTlTyFKQtnONWO2lWG/gHtOmnLwswvFRhGt5deiNkDbCtVU+qm5qlr0UhiAh
qLn+s4MHiP8p59WBWWRNChoYUBsDVxLeWSwnECig/aSpBeEooS+oqTuuv9Dq1dHdzs+jYaZ7w4BQ
k//qXMqafgU/kTdtCaKNg0d9U/B42l/xjZHXFj47cT442BOoupwks/NIc3pJ1bam9NDPYRcGEMlN
PaHgFNrbYMV9DQt1cuslL9L74mkkeCpsZDZSlqyN2pov4bqICeHyE8j97yx63QWqcgofxj6Kq2RT
HC7G9zzdGqbhgHHj7j7GHmPPs3tFV+xrIUknzI1oA1WG+kTEXoUFR22Yw6FJn3p3P4EqL/ySNa8a
g0dajx2kxKC/o38KHHDEAAP88+r5viQ0wapQysZZS2g72O0v+9KCihSAs+9zxFItsXkqmyWL6CKR
9aP9Ge87qWX00Hbmu7TXgLexnFxRZSumOaU1ZZ21UrttFL0ioN17kgBrnZeiXnufTsIRCmx87cN7
GYk4t1MfZAhte9K2/f8pZQjLr/w3viKnOXDQSLG8KIggEaad5YqFKXCMYDzVKcwgpbnzoNbrXFGx
9Og9r1//PT4savx4Ue7foW0d2jCoX8ClBNXkLmB68v+RJrpxfZrbAZ+tLDxU+xmPAUN9xxjmHUyF
HpGZsWIhI4BRdSPVQENC6xrnWJjA8j0i5DnL0uV5B+Q9tluW6oh2TsXzikrEVFWyXgp/gk67bXIt
UsuXGbZSDkjUpktoYsp8+v0kCfJW2xxAZmaei3TCheFPfrgAu3ivJ7AYklT8nhzb3Hqrbqk0+Kh6
WqqZwHXCbkblz0Z5hLNzK9WQRocIW5QDl4IBhoIk4SOjv4N1/XUsaSkzzOmmHMAP+FRHixgr0uAg
gcIWxztXPipvQhtWQglRLVWAC8iDIDxo71EtgYeIEmVTI6SlMc47pMFXbc3UWDR09hQVqgl0jQWO
vXGjtKAPWENLZ5zvoIRZy3o84jA8gs/y0VDNBAKzuN/9wEtl6NAdVsM3ASusubNFG8YvElGx6l5D
icZzWCXvNnzyyS6TA3JWu5wgSFiMdP5G3xgNXrFn8x9F4mDMh2qDNhGSjfIHGAmYhv7mSQiF85WP
mQQ58opph4m9uR7cL5z7JcjESkrBElNwotX847Q6YMk4L86TMigH1ExIv/sReBcAbQyXrdoDvsW+
LVwYEx6k4/VgFfdQFJBC8mF5y1Kl5LhueghdcMrloVE5e+1S0wN8m+6N4fLyMSE93zSiaya+dEWq
TvqWc1UC7DeZUdwXBVxr3fbRfTh0RWRc4dKVpAk98XM3XAOE8DuNbzvWHbKFxnO9HKYi4Kd7f5Bq
zj7+6JhHzPwkI6Wekz4279YZBmiCTN+6Qs9jVIWvE/aamJrGkUfq+xLUX+a6V7b8jrAomYPAZawz
QJZcqIByQrKJ1G18Y3laPCdgETksEbVm4nt53T3WY6D3GSKOpeCw2wC5CH9rskeXzP7wI16S5+10
2LWKt2+XQOG7We7BG/15kJVFhpGFd8A6odY7crDA5dh4MDhHlHzVsGnAUEWjTGnRk41xf+LJuVEm
07KjhQ9TzZPwmLms9otCerZrfb77o6I9FPXRSdEbFldzVfF+uPU2AcnxdkPO8C/sz6xkpiqbfYbq
ekmkDZzChOPVvGct2Cu2mrm2ZOfT/GsDIT+uFumT3Kd0SC8g1Smigz62e8sGYOxxWYnh+ElE/xXV
TpxJ9izSojtmVsrov8CWrgyRmFoMGuMq1xaIr36AjGN/pHxa8BaF/D5MxINCLFIWtj/mDNGf8gzs
Na7ZyjcZpfF80yndqynG19kkYQ2Wc5z0+c2ubpdSbEIIdnBtb5YZgjYLHRRukTwW+MkMAMPYEQVN
pCZdjQB7wYHRitfqfwn3zs4GkloxtJBxyLyFX7dyEtqtyk1YjE+zZ7ucq+o09XzngcFdaplJG8/3
Yntr8ubau8jY3pgxrpJwsVMau9ZuzsudCdnCdgW8vo90i3PyT5HyywW7O2roUFLQtFnMzPhZ8/sF
woZAAWe5o2/RfTz673gQ/s3euulpLZm6rx75IOw+W47lGtwQiI64snXKgv3vQQvwmM7b0XDntmvp
qthHvhsL1AXADN29QR1h/ffvuBh34n05g5YyEy+TaOFKCP+FB6uhNBQ3an1m/DhXJ7uM0aIoYMWd
L2RA9UsaLExsv7kz+nEg1mORLz5poFxAbktWL9wlEj+aXyEwzG7N484lQCKb2EwyRjhsNbY3xa/e
aG+tZZ39T8yL+GN8Qfwg3N7YuEVZwHde7uh04sM7aNgi17017HyRrHcpUt9y9K14wGhiqeZNmZ0c
bslLDL2NGh0W6YwATGz9CSl1mQE8cea8deCsEZVtZBdfvHe3/raSoEku2KxMfKK33bN84AQtqfmc
LsszKW7NjxkULbLtzjr7+tKAhPuRgVvpszitayjaFGVbY7bl9sjj0v4Akia3dQdfh6qb2g/ZhJtd
7E6WW80q/H2tUhapnbLNuYKHoleJI2HLK7b9ogQbkHkE6vphzHS9RT3gArLb0IXdIhsT432++FfZ
ZPim9KRzLksiMtLeoi6tb/55X0M7qGB3J7u8QCQBvLMnwHv+KmzSiIOi5iYsK8t7OBstZRp+3fcQ
7kh8jJvYNs2VHoYAQ3uF9RcnhUlgYrpDDfTNvr2nSzF3PcoKcEmQAjuVOMzpbZv6L6oUpKCeyPRI
hkjZbMUcmEfJzvuj0WuJSMpQlfqeJ2ItQwOmOU5okacYFyKHR9Wp0/QJsW1S5KUrmXROSX1kzu7P
lKIudlLkm/ZJ4/LYjkpGLSdiW0CHyZQ8oAeCxMndXhYnut1JvljwTx//8Cs4A6P3AMyapJY92df3
DjtzFy4Vl4XRUjz4VycBiRBE7M43WseZ3oONPYfW+jTf7G0sqwbnr7Yqoyrz5R0V3QHlgfyKMlsq
PESZe9hq4zaf1vfKlgEdsSYGYAwKXu6BQSmzwZFzBTPS7iyK+o4djnMrrYb6fETpbnRMH2BTpeEP
fFb7REnK0WiTg/ggZCts7fk4j/vv7JP68a2pwQT/5O2wIbIjKqlu9ygQ+oIB6frjF1BLbKPJjFII
zqlrfwJda80NERjyLTjlbR7DwyQS3dyoAfpwVHfLFHz7PRVp8zINFZ06hGkMiMiD7YuuqQyIxZ6K
+YpjdEn1pHHH0ow9AmGzGnVNNIw0EqQow9y2E6wwOmQC2WJKSUErfnTZ2HLDKEr3xM3RBdfCkBul
gjYP1B57dll50kU8RJ+85Lcs4VhFoqZcZAW1RQoXcA+NKk7GY5O8sK3BFGk7Rdsf/8tzqdItQgzq
/SgRSEl06dtZYV90bTio4i4d6WpeGKHpa+ZAtc5KkZjrzr5rHYUl7zcYF1ugNwtTekMgz76ObCaa
CJxf54rDybdotqLYMP1mMCiF1yJJ4qn7O1U9Dt7VVXJLIw/RJBTv3bB32HN+jXrdDYeYLRTfCiTT
/NHam1oV5UzaibMCthyxkUN+YYt8zv+84rGoMiaLFRa/532eDXox1BU2XDj/mRgUpz1Y8T79VRiJ
+7Cl7a7OLMXB0MQFFywrAEOOMLuxeyGdLzh0MJA1tdSmrWBtyW5O4jUSthF+HFjnBm1x4caFm6RH
SXBH7m3y0NnbgnbzH8ztV4IfrkVcOFZx8kZRgdiQ+5XgJ/XWGuCXNiDaabK513GJca/h+76N6pkP
rSHQg4UsjEn02VuCl46Uzza4cqc3cyKV//2Ljw5a4zk+cymvvdYGBzcQR/e5aae1ihTwgj2tOQ6e
9Ho2qgyRkodyW9uCvlc1H2uqupfqr6yj70o/6bhYfvyxjO2cdcVD+OqEIt0syEJ0G0ltRZwe/sbX
an0I2G/WyQGqv+OPnXOt18RE60073GcdHVNS6EDyU5ZiwlqzlxKTl4dtJVa5J9KhRH3hUUJhHMcg
Pg==
`protect end_protected
