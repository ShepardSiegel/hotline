`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZAERTISUElexK3YLlFDheF3UYAk0o2DJm+t/UCD5T/V2C7IZBOY+dp32X9VchRjPy8z+rdwGpLjj
Wi62pG+pNw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mIoci8+H0Bw/hZchw2xSxWnxLghMFNLoMdLScEqBxMlqV2bWvQFqNUMifYOmFQRWKCiuwn8v2oNK
jwGUAhkI3Uw3hz45IBb9bqLsnCOUn3LGka3sWsH0VX+JCqI5UovYTUafBdQypXCXMvNFs6tu65VW
Xu4pUUPpKTQjX+m9inU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jxh901GHWjjoDkNTogBP5DHYqMJUIZoXl1O0Qj08rE+WbKggjl/PA72SNC+rzdmjG/qfVwQhp1n7
GIYrlaKJgp7gKaT/bdktvFXjrsqD/W1Bcpla3T57R73Gmgxig42dBZ48Xx++6KzKANBBlkHiHfvk
yWgTKfpPARoYQJNC44lls9Ke9eFJncrvZyG21V3caHfidnGnHKOF8S9g4PVfRSEDt5f4qk1XfNxo
/MvR7QbQKQo3kee5FGqOIrr86pWos7tsDndVj3KBjor6mNvAGt5aJPFYQYDglJcnPYpLvY9ngwM9
vI0iwL1OvCHdy1ebZUVseo6I9ZDBVo8lrcu/pg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dUdIT+Jov5FUjCCkutcj8isgFkreXHfmELy6XNxJUGHShhsWmEBhsgV8dWoWq5HlrS9V8Oyz+M0Q
unby2jk9FY2wevcwAH6gL0UBC/dnJQJAcoUZjIl/4web7Rv91N+nD0Y0sGFss/ow4MRpTEwdk5bs
9v7J/1R4E5ueyBeZvBY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nD3cONV6DErXbtU8Fvej8doo973oqoHBjcCxqRqgOzyA1s6n8KCPjtU02xfmnHsxrC6M1kHfFjGc
fSDQc0b2ArAVmBGStTYwtEBVeIJE569UCCqewbO7NcdEUEUgv2HXQQIYQhHPci+dgSnjpAsCgMOl
Sq2bEMunmxbDYqldZHgAF4H4H0GEHR1pu8I6U9AH3KgEZLM9MPOe1fQhscCKEGVugVo0YcRZrMbi
y5rR3Qxd1rpJ4A1SfW3LNxHaB237MGe545+DVfJ/jOIcHCy6IE1ibT4uVAx6mGeHJid/Hlh6Vh+g
sBiIS2vgUiGVep5lXhekTreHu3JLgLOCssYO9w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5616)
`protect data_block
Su7NOkkQ9YMbCLVTa9O78Fxu9IS0rltDrPhEE8zF0BwdgGFV17tz4Z7aKDTEm9XHsODK4wq1wHn6
+V1jHuiP/dDgLoOOS92me6RKA5QRAVaq3pNcyow4lIBuxI5I2/erTnhpaykgMIgh8t68qgcq+GQR
LMKWhQmSXjQp2tVyIcjDZ2QnUpbcc81+EFBrWjAZYJ7ENfomb4WYMqFwaZ7LibKoYQbdGLQDhEuL
6gW0bmAcXT0puqo4OrcI4c6Yb3JLcBFPZbuZ5pir9Zkt/n4EWkH5cqrQ7enFNiJn+/G7go2CX4zH
1/Aawtq4QxriO4qKjuzZtR+eArUo1T7RDB2eOfiMtQLW2RuXSqSbXY5mY/5xhbU+Hcv/ZCk2v28+
KTQE0zwlPY+EqSdZcJC5G6d5vmSj8TWzich1kpAh4iMei3+dzGuOn5VG8HXuss2FlvNsp+ARDQ0g
5J/3F22eYPNsMJwrlnerDkskDk7FOocttt5JG/wHS8ti4pyNzMLZOr+0UOPmt0CmKXwpbm2b/pk8
z/EThdnG76pcQCzJWpzNbxkMLcP5sRjuZr4mcV7CydF02YpUg6hr1u7rqRRGeVVQdw5g6hJZ93ov
mcZN2ABW/V3V9f7NPyzIOF63nYZfLDDfgqfJGZIBEVVkfavd3GKHARo3gOAlPmbjPZL2aT6sll8Z
Es8olse+S7cnORYNoOp8Eo7j+EZ4Y+CxNNavLcgsu7hhR2U28fy/36T1KitijLY4ZMMgsSdf3uaa
ZopDHMrD6Y85QhVGCPVMnDnrRoUosQjmpfaH1wB5hklQExKG8zS2e52nOWPpiI38hpBW+Hsor4v4
aDeyRP3cxDSimMd/QzMsIJ6SDyLD3cGUbGYR9ls/teYJBT/MTbZUiyFfNRKEbi3oWoYU6AmuDyy2
RfHrV4pAZATDx44jS8c5lJwlYYe8NddQOCQXU22neS+wFHKRc5lTl0ckq8bGaQJ/1ZsW7IMKB62u
VGrIYUaqhygr++cJX2n7jY5DGEMqwGaSD9OzKu4N/R9IEct74Frb4Gsq2OS3UfWK0HldTsNQZE0f
nyDDG9sXLgIWwrExWv3L9OV9gvvOFxKV2ZognH8Kma8WRtxS6pIbtfllOvfyBiCKOOhzaI4k1SeY
9ZDKHQZAYXJc0SU0xwRpLFOQGZ12sHTS74wrMQfwQHuA9ki3YwR3O4VflxwALwmCLH8D9S2xljii
UT88MwRBvgYsEd3bVODAtc1cCbyCiyemmM8paYLvirLO30vzLVEEwOhdP9GnHAgztzNt+Ly8ce6F
bdJI7zkLOQx6buR/h26+i9WqxXiIvIrW26YjjEohZ8mGaBceZHeBlCvb7KWsdYrnd/B+B1wxfnux
1oZxmOdilUoMeWBMlJuhB/U0AbMCm10nDfAgZ6Lpl7dWTaKgxr6Q/GsQ0TXMDvcp9uwrhf0wsH0p
CbE9HGTw5+JVRywxR4Fy22/pcpRBHl3BiGrIiJi02nyA/wsbpYzNou14pQ7Uo/pBnpmzchefc1iZ
VfnxaMQ//uXE7NKzf5k1KK4WTWy2uEjvUzKk38nyRnBqi+AZmJobAnwYvbeOqcjofz6KNu5/u2OE
rcA4xDvhW5Pz1DNpSdMeRxc3+QzRG6Lqt0gelFPzm9HfczMdJM6K/enKRq//0e/YCGVhUp5dmdt4
7wCrQi1zD9rUqsAtWp9omRQn5MX4yadqJwhM6wVoQx/PeM046cI2D4ePG5TqDfC/v7YXJMSgyFFt
XDC/sVff7NK8/ijoXCjsMzPPqQdRZCFkUHPqTXPmQcCaLT34RuDL3XovQ+NKqKRNO+Z9jof115Be
oZt+pWrFRN9GdHNgzbstTJavLKm7KEZH61t35ZznbiD0mED0bXsiacDVth8kTEwTVQEpuaENIx9c
2AcCcKvTXDW6sk7SUf4E4mQooM10milqF1gIuXfN7sBYGEhjP21bd+Qy6r9UmBy+XCOozxfL2QIi
vVDcvDK6IsqLbOjAxlQ2AfX7dUxs6xvPHvZqOO4LIVWRUuJl9xograe9h9ikAZLKLEdvi3Kz7R+P
OAnHlHf+j3z3xwF4zlMIrxa1I2PrXiDn69iVzf+f8g4LDD8qWlFKrFhQKMIxtgg9JKQzl805yNd5
JnS4K3V7LpQaIOEoQxE0GAh9+1HIH/lR4S4E2UXK40txBqufgLJO4006Uqillx+TMp/ZjvfKwI1v
RM5fbnPT4ixHlF399imG4QunUKqVNapcbvXk+zk9WexBNjZlHFRY4l+Xn+IIWoQOqdja/AUrApGh
BuIo86ZwMA45k0dWararMPVA+FN2p4Dj2PUtTxeANeyUz8Nwd3HJyXcwNOKdDyzt/oYxr4thk0lt
/FOpXB+Lk/FZvFOI0/fyTLPHjGW/hYq6rq/8nG07SCKc7GxgrxIETkIsq1KqByj02W7I2mEOQ3Un
xueVw+I7rUVucxCuAlIxTd7AAJcyc6JOXWItXg9a/402gwQOu9rs6H5LVzMiK1yKnYLcrWoNxw3R
3Uy0tKBdNjbL/DfdAOn8mWoFRlqOklhWX3CQvJCh1VfKnag4ch8yComKs4JA5McBxvVnXyPlF45p
/QBDCvNi17G5LzlPvLQotZSYf2c+yt8X7KYjpHGmHbIiyU2/MTsW+33LimCR5pAJSE3/WG24NtFM
BtcFpOgfyXREmgW6chtlFEXEwgiaQsgVvavyJaytKYtSxCJaYDL5Cb8il3v3OvBaN53Fliy3ZoL4
Zj6LkoFUAfNaGAOGyfWo1VpCb6YQ6KyjjHV4yllRvW0MKbJdY+X4OAOf2QtJ19SBMkSbG62uPNP4
6uwUAj0C+4mn0BhhfGASkSIcxuqi2idzeX/ZyQ/+wwt+1rZh3wB1GDNkUtnS2Oqtn/uIp4PixQJ2
uYQWtnBfjcC5i8HeNTIBeI/slFBcIlvUp7FfBKNvwgVO2mR4P59F+klnvCMcWLJslFp/vDSgMJmm
bCFfZ4Uw6m/eS67lNWh3UYVcv7C0PUx5wPLG8wUPc89gW8ghYbKy+eqc1W1ynmzB3IwnMku2vMe1
ojN9WJNKmnlydYASzOJrxTuKYJftYUjIN1Yuxin5jxeaGsRoCeu+MaqsfGxFHC6ezMJ1QgleQa6D
wcAQyV30DE43usGavA+qVo+u/JJ2x5RHiDVf3JoeVEfb5bbVTENDH5uW8tSrO5KOZWhDRyZMUN+H
oBfdH+TvtBSvYsrnGoYgeS1l+yTnEfuH3LFO58Yyu+zn9+RL8lvP4nhZ1evsgyw0ZKjG+Ng10kLU
1JFOUKrnNk/LRfOTUg/36YYWCKzCYfGOiK3ngNJcFDj6+g1rZnMCYFj5jmp6wKw/AX7i28WVFo6m
VgZRHqdlevbbu1jReso4EENdO2Iyi3IwISf7dXXayeQwIXokslc0YpnNWMBJ7dFCz458evDiWQVy
qQKH2o6fOQg8gtoWYKlWWGQDcum1xVlNubaxrSTK1D6TXxDkAi9xq3HjolTc8yrsdRY0hx1z0BnV
d8EqxJjAYynPuP2hUUCDRGhr0+o1g2q0rff+XhA+09hfP45fIhuFHe6d5wX4VrUF6m8FFpBvSNGj
MmJKuLQrfLFQeolGZovbqdue2CCt7NyclAHWe7PPc/aHc6iRctYH45FX35lPNQejdmZ3yWvFYpGr
SUKGsf3X05Ycj5HpG4gj1KpZ3l2Y+XKoBEN9I0D8sGLoUSKu65y/53399Z0hOJvYl0uabZq+QtOS
T2h7TpsXMPDX0sxyw+Ncm4DnXtMbY2/yUP5wSRIVVRgOFOroVhdPK+IuYvWIP617iNpf3t7nKKs6
hNLMrOW99kS5cZszQdDHS3gFMKH9yS0QrUWijLFD/WHI6FITWjym87nf3E7NVcoOlGThLfwqGPkG
YFl5RJKmbCcCEKKWOYvehytZGzjZs/caeSqRXulvZ9Dyk9LwMZN5iJ7/PW24XMbf8vAvlf5PWsh6
zNkFJViLzVaXRSnXqaZ5Onfs9OnhqMA50Nu2kzdGpaH91ynnnYDVOCgXT81NRZMH+NtJNdMPRYUE
kPbf0Jm/ngWy3UkYg2n3D7vMyXU1VwUonHMng3NyD77vVeDsGUEk8sYJvQXFKPORY/jLLRLqBkbK
UqCr2ISJ3ssXHCW7vxjdfEaBsEwvke5ro0yAT5brEx4Vxi1S671IImWMGaoiEgHh74yiYmuwNVqu
Y/+s5FN4Sh9mgxs/oDW6/UXAH8scjLXicgpUbPMhoK7p0+h8IwgKhdc4CNHiRamCWL5XK7iN0RID
GTrrf1yERfyEzLDnAu0SprJ+q3SGhJ3+mU/Iag4npL2BaP5xhgIYw23Ov2L8DDfc+MwJGy99uD3m
02dUDwoJR85yx4oGViJJlT/DikbidpIHNcm1N/4RvvMpSI3CxqB9wKTN1Fw7CFTtGYxPruigqtN3
Ni/CZijukqy2Anp7b8ecTyb/Kc6L3q88d7dHjr/Avfr4/sH1eNy/wvXdVF2gP/xIdi/sCdxH/fca
KwRsYw/3eROCnjPY6CYx+9w5m8HExNRW+/JI3kkB0R/bA2ps6FpshrdL7rm7knpDl1lUObYZKkF4
R+vChVKBQ1pRBKJxXHpWtHVvHH1mLO3s31fW9oe5144w6VEEbWGiOP8OoQYMgPnS0rBf8D35Kb3h
6pHzSM/rf5M7sz9m0c/aikntss9kORTDCTvB74deyMNydS89eDyPirR+jnln9i5Jpz27I76tnN1Y
h1ccHkqtBnsH7RoZKbzm/uVxztiOf1pkioLAgWjiiDNxrEgMxjuZLw2GBzuWU+ddbgXiYp0bN4Ei
t2wTCArh1zY1UlkNKLAnsj0k700lTRhSDLoZ7zA7bLsQiD3uldNuWaMU1DrZBDVQfdZ6AGZZHErm
MTJe0BcvreVgcUOzK0JcJe+dSMc1zBbH//CJ2S/jhGHEefsTdY4G4LE5f1BKu2qF0OBo/uU7Pd6b
olkllzTQ5gABZo9gl8B8gtUZ17SV6xUNOP/jzFzMBC6Yw6RU2PCcN1FHi+OJ3/vP/Kssxjr4K70C
YCWRVBSWIn9qbXtN3IUrVzhRdCelSVqXIkMijOdQ8ENF6aDemR5T1cuHQ4F4hvI6BFnWt6IjsdL6
v2DLhHfueTDvXu7zaYSOgTH7ETn4KCc7Weqg2l4th9OLFo9kqjx0HSNjHWf+ZeOHwQ+JPBWRY4Bd
zYZ2cThnjP7gCP8bDq77rH29XXaQodR7HZdYHvthCYnnT0eq0knULszh+CR++Jm1VUb8tyBhZKks
cvFUw3V0WaPZs31WEKnuKBp6cBwrYjyPH5Ua8BprtRP0zaIz1wbzJCA0r8GTFQqPmiuzSeMxmD2r
Bl5tj62FRMJIjBkUiopVQUV2HC/kbNAlg0Ol+PEoZrbP3gdEohx2lctJrvG11YqIsUrSN8tP6R9Y
v5iEjhTFwv98xvBeNCb++IWgolA+9jOXjRkbELdkYEwrN7ROEDx4sWckf/6JtOR+6VmXllw3iNwO
1IQnwn0FKHBpJUuJeMd0FPcrWA3ixNmMJfD284yEegBYkEtnMH8IZQcpEIngYGN5C/TJZlQITBss
e+LBrxMq04ae167U/ZbIiCxay5EuHshaVmU5ORi3t5fywaq5ox+ZLfYxdpCs81rYGA5xvgRkM1LZ
ev50xgQev+R8XMlykxSPhUWBEUamKc9mMUc71423nCjTzzvFiOl3zMRy5t3ontf7LBbcZXjjSAT3
0fQUdCY7rQDjOe/JybZ/T/0p6PYY/+Ot7TgZsTPTNfJbwGBkRY68Qb6OB3RHytGPu51hSeB+0iW5
pfP5IRgrI0fjavqsYwuiDcHjlqYWJO+Pw4ecV2UDNtryM+q0Cr8LkzxS+4XlMc1gG1R+pvnLJ2+x
akLLdRKeAbBHMN89WZ58YkCbu1Izthixq3DTTelpZMKMBuCaOBaE0hKGQfkgvOfOMKDWlVKo+OUE
DzoIoQ30Sx1QreJ3F++dgm05y1HMGBbTXCJJp5TUmssH2bSaXMhyZJiocq+r31ZYPanjVwXRmOjL
lqKpYm3GgEUaO1Sctb6MY4UnzMwoa+FfJwnHZ5dpnON7iy4MmDGSGL+aYcwP7L93P3NbPsOcyFWW
BfDc7iDdHHPpiMGBOLnjyRjt8XltY6T3VXsuvBzzFmANY9aSzVgwMXfkr8GITJ3sEMoiiVKjeFgX
K3U2H2ujJjZMEUrHNMB2QdpyP1dWqZaRKsoED3VNO3gx14rAiqZ61YlcNBdaE+xDtGi4WsnizVDu
Igd0EBynamdf891PCupborpwXKRf8I5yi+wqwcGDEQbgS3z4Etwd8/8wcQKi03Bbqabzrrv/SHpq
QO2lnaw3yyL0GHWkUSYFmjedigP53zchoNchyT8K0y10O61xy48mO9d2Rp1VVSMWFyAb2lIRiCyA
UkaDf5LO2BOBWlbXBwbHM13L75h7hVc+xOHMmksWCRW27SNWMx9tWy5CBj8tceBSBR0R+wvMn1+5
J79pn8fB6Kx7d6fv4AncfNoirmYZPR5HOKwBx400x5gwpZdev4/Tc/p24xqjCpmCaqTSVAB+LPvy
iLs0fYQrz4IOT9PRVUEcxE1GBjkGuTCPP/9YpJYS0Kzmy2lhDzAl11jaQlYoeiVky1OYm8FZqKsm
dDUdmftFQIuaC7XWMUQuObzAPaj2ya5YECMJrtgId02N2feynQvnMZJDIKaOYa5EjUU/6fPmMsY+
9mvQKgLy+1FKlb1DWSzby1HxIVbcfZJ0RfKqlZy1GwS/QQMQggGjceXOshdCjEHp0ZgSgZngxlt+
MznoBEEWS/8m/PEgTSmxK/L9nt1OTbnYDh2zS2lqqgy0T7DFAaof4xd7nLM7qA0tdGQPCC/IsMmS
UACOqTLogjXTcNQfs8qKI/0qMmtlvodGLFhtKfmPYf6O4oWqec235qZgK5oww+ODX19hw0grNEqv
6wHnOyIjoyLn2HyL6R3N4RLFdTEjNKqWSFcric2Lb0uwxtv8xqvYARtRNsJdUh2fLlVn+UToPm5V
PoMpToK094rNcfF0dyLHTlzW0UpbNJgwl/uYVQ1/JkxJn9jSlvip+5ylnDs55ope7ubF3Xif6GvN
F0Haonqo7EJJzJe/MmWPyRUEtRfa+aX/efI/ZohxNuvM8xHhZ5O3VOeA7C3B886Dqk10ysGG0l3I
2Hmi1kKW+KwBoO9KISrrIh3DGTpQppkHUkN5wdGgF7E1WMWuCHG6omHTiQq3Hiiom6sqpeVdt4+P
aHBSKe8a2IYvLCY2kzGoQCo/4S/c8f+ZknUaeDklwNmQj1nzfqVOwPvOFudZdFbl4RiOh44d0Z9l
/iybzmGUJgx12DPvfL2ghtR4FOTyyaZSrBSIjjQMcqMy3S/5ketoHUgt6DzyCr9Zc4qmvZ6Fu2Vm
7OXaAZ1XuHcuHQfjBuzAjWT/xyKoiV7sdNlaUDx7zQmC+ody77VYiFXFW9QZRuIlbOGVx5SHXeha
YICOQ1RNxwWCe/Y40Xy1xcq1p8/2aAGReIDPZJC3
`protect end_protected
