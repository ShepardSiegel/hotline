`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gXe90db+1HClJ8d1aHd2oYl1FGquoZWp2MXh50OUOgn65wxlea6TDDy5lThX4QjZRJQ4dPRE5UYk
Q0CXGNEgjA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VZOdjyZDsUzfsy8REPaav/3A939amx8ElvsAcyEIsxrKjGqoeMnQMoKbs/+JeSpM6bcBUFbpsmbT
zgKajGIca04ZAJwKzVSCLniWPZLqU6D2xZ51ccdHfS9UwJY0/qZMz4UrBqlQeSDkfKyO6met8Xfc
kTG2BmbwjtC3y+vkVog=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ul1azkXpOgHx+qFSd0TOrL7EznzkedDMeCYDUmlQoJpclsKyWKmhknx+CBXo3oubSpsjoTlHwEA1
spyRZSxmUNqwFJ/0J71jooFA1Q+x97Mog4UNMljxVoO02kXaPdu+JdfkVdApaqQp40oKRtDrw5UX
z2qQZmWJDXqf+VGXze8OykbB+Yaia73ywv5OJ4JRvtlxqNg0LyThKpQi8QlOWnLKawAn7J8JYQ1J
By+Yz17wnacN36KWxQGxEwtt8+YiERCxglZA0l+aExy1+qQMFZPN3AL8B+pN1isWNU0NJxV+o2XE
wt989NX6yO2DtYjyGyqy1+W6MqW5ypZzpU3qPQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4CeL1foOCkhJ+fFpq4rlZB9uC+ZD3/MTZsDN4Me60LWlFZAaiSdiE2jhaSeJcT7HpcoyeP5L7JIX
9QKHJ+SXab/l7VntXRpz7oX3DyyGrJ1JTMxoys7GVy91dpe/zY4541PLlVjaiJ1suWCKrcGjo/tt
xysUAAQ+57zdohdGOQI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hAWV4Uxswv/x6xEwTgm2xw9FdG+AoWEHF1P5pvqk7+Tj0iuB18SMk+YPk7bku4h7mNFEAf/AWrhh
2MA3O51bgcge/gsQ804XFnlL0rqYXhvFHtcK0aHBzovZoA80uy1ueCbo6sKbjsCrtqfj3GcFVCuM
WwcSbEmB57vcFgsj54bBzj8MlJomoCbdKQwEKwpDD4AKz8zcSWKy/s1CZX/PDQYmdMsSQfeidzLv
RkPabAF4uFGp/unOh4JG8mPMzxAKPo0wq8x9wxi4ElJwKvYq9GNv2K6Sv37OjKR3dd+bq+OplcOz
algxcVXB3cEWiPEsse6zvPhUygrghgsOdAl/6Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30608)
`protect data_block
wl/Le5URYUIuxmYV7+D/hslZ7HdutnWNEtTzpo+RxpMGUzza+ZTUOE1rIReJ6EgEFrjQBBI7wIbn
ASskxTf8/MGsvxdO9VoF9G1HtGBZT/NriXtK7E+MY/UTZQVuoUUzfHgdHilUyKLuwINgNXqLSLRb
tfJA7bV1RDsZuk93IA1zjeciafS9MeNe8xy2zyCsryyGPypKHBX4oAs6jlrDSgHa//83BKpVZ9Vo
juQFr/XdulGtQP7fqUhWrKgnbFoU0qgYH+bjWnBWQQqMP3C2rjAOMJi/b54aQEjlDQQFLJcYW7HY
Ao3+h1FAzeGpzyQTbEyfeMaoWuD2wZtgSX9ySFqIOBBkn33gGhEqpkD7JiGbRLxdJjq0qkhBTTc4
PbvBmqggcb7h3h7whbq1Rc+NYsxlJw+zM+/LPMou5CVx4S465ESgLI904k+lsYYQEDytjJiK9Pn/
2RksjHMsqoZyyWtUe8ZCHtuO230Sp7PyVkJJxdLqT/rvU7Std9AJ/BDdW3If/n0WBvfdHskVcpdP
rTia/3JfZ67jO/oRqNLosHEbOgKonBh1gUhD87jhADq8w8d5jDaei32hk5UuucTyBU2Ze/c8jx5t
L0TF851LbSb9VQNdzHH4Nwh8Wsr3scX/TTsOMjyKf+ZvFi3jHZ7eHfEUhc+DwyWrjUp5I2blex9v
VqYLsgs4B9IpboWpU6jBv1yftOD7lBTar+UWuUzpl0kX9JjNEV1qCu78eDvFE+0eex9iQBGErAoy
4rOhghi3fVEaNUKAJeCKSsDVt6AdTExAPXjww9AWFnfyVw2f5Fw8fggJTBxI37cVDTnzlp+87L67
T3jzMFKKZbuv3NAEyWdtPeO3PNXxu6qUszpUz29lYMB/Bu+hMM6r0BsL4d7e36as3q8py2sBF0Mw
W5mylRBiFYo+lmHbBfPMDoCUJW8UPqRpQRefRs++MqTuKkVjT/A7oICEuHUihFdmyVzKeU+nT9j7
HmJSxHFzIgAu+r4T7xNI39kMrwOx08h5ffEQgz5PjtJH+m+EPmXZjiTXdzyyqJc6b+VoEW6swgCT
9cIs5wsvY9LmAlE84kV7BSoya5xQudy6kxQg1OTwNIfsKuQ7iHSDQISXTOvIXLeTKw2c3pL1wTyz
8IYi+f64WrM37NPCJ/gE824cTzkYVD8PbVQNCmFTDMeFz6rh4GL+UFg2sIEZtGA2jdimQppYu+3s
nDsaPLXBIJebzuidOiMoghrIxMUKLhBlaMwd0ayWg4uYiOTAK005y63+MHK/0IOgESKAZvJM76du
lzuOaqhL0kaOdjPTMLGPo346rcIzvMIflwUusmjbvINWok13UuTO/KD7wjpwHD8eFTcJgq7kAiRz
O5A0Xup0m1BI3F5Qjd/cT0T8gd1rBkC0GovqXeK3Zj8vnY3jFRPsj/tznQ1RHW8sJP2tnRF91G0U
y39B//QUo84z4AgZpNFfz7MqE5fzluJjYt0BdIK17vKxfKU/YkJAmZvmZGCIceWX6wzbj+ucmSA6
if+VTVXc03N9l4jDQ9JINlMsaBOaR2MKAJX/zkPbZ1kbt+Ax5bDCwEkL14XvqUj+uv1ge3MKOj9H
KFWFzv9WjTGUtJN9ytsa/9uENN3LyKO408iir7eGQp4jzvK1RTIcvwUwJnqUJmL2oawneoZF8mQb
UTylrq/IP0IT99einDg/y6Dd0K6s5NnjxOf81VSCiOzYdHI9p6wmsrlYd2pYV+h7329dgWIsM97y
Mz3SS1IyyagDhtie4Hph24gMVA+ToJIbQLYj2IcTsMDzjlmeV8Xaw/gUTxM5EBR5l6nCHIZxhk/B
5WVb1o8ILlmg+jSUZsf7+JB7HiIEN4FtIEeTaoO/4vnRoWgHLes4OBFc1TOI4cIQrvhvwGbQZoPR
koOIabZgYFgrEWpoUo8xH3KDlXC6Hhi2/rTzbUX4HbOMhT4bKn5spohvV5QBvfx7CyEfWK0SBfSK
2VE6T8oWUQZFvsBbLpdKR4UqqocFf/ZuqG8ZmcJtavhX8Ejb6cZwsZkRDizpFEGASoQFo/vc3b0k
B+1y1wlOsPzCIlN3oCk+6f9Vj+fAUWK1Zlvw55XX93GiMl16jBVMEEsRVuBg+m3tcp9OY47XmUCj
nydk1H4odh7BGsja48lLHFVbskUEB5dKtY5r5I0IdNqX2rkVoC6NxAij7/ocC9A3zl/xo5qESii2
tZpoqGLNJP8vzgWTjdSjApRpKGxdw1t2JtcuK+qYIeSF+cC4qMQoz3aGUQUz9g8LdBFCc5+9FkW0
F2Q0yyvqV09/i+swAUSC0cBSxz40yxjdQ+JN2gWt9KOobxHZqd19ReSSR+N9ddx/CbuHPiOFatAQ
7w0EWm+jeMAwRbOTzgJP/PV8l1fs658lZYB6KkM4zdlLcHpbqaOCimZsOTT6rFC0FWLMjWUEpZSn
KXPREBx8ANTCmsIa0vgvjdHok7+3EFNyERxfgPKh/2of8X6xYa8SmCU9Wc0XUrI4RLmKalB48TLR
wg+INoU2q+YHvXjVN+vaIWHjdGal4aFmFUf+a1iU/tPjROQNJNE+BDpMFjCGSAFCaQub3xD80PAZ
95s2qvcbUF88O9fQD5Ihl1gmhAGvgiOSf/qLqflj36CU5K/u/fH9r60/TOF6IDJoqYxeeRNPXj2I
X/Q2Y3LooU3qBhSw5jIwh3p6dx55Mpoh0/LlWjfwmMqdL4IELD8FJ+I8Fte4rZyBCRtYXZ7fes5M
GDARJD3hDzcmw+GIf05m4PwMCOqLnpmLDk6M/SUdmnKVw/y7EzAWvLw33WHhoRJ0dyO2DcHDtW0F
4hiuCb+8uAw4t0Ie07WNnGDUxNsN16iNNsLKXNrGXsucCyKcq6rhOeeKhoDeQG0gI93Ka57+UHYf
fctu1nVzE3MUswvxT8Nr6ktVp+Qffw31SdjFDwvw8ULptFs1WTd8C7oR6heevISGAEbmCloQDQCg
7kXIIfzayAWJkLy1M6q5zVe7i3K2DciAIG2q1XrH/CcMIJ3e+9OQahPj7tG0UM5O1sxUn+zlbeUC
4wRh1aCTZTGKdjYXtWnXsk+AtRCSHlo3izNjaPZQwK/kAVP0xXekdssZ9Xi0rGZ7Nfq1XsLnit90
yP4uQ8191GepJ25URx7LZxsIIOMftiEV9X/bxfsMDgU/l2rn5wz9dLYH1ttDTcbud9db7Bl3szfz
EGkrJZXXBvZYPAgCYLzWh9fK7FRb5vG9FEDKK58yLMBHobySPrpwFpjO0ATK+t3+s0PenPzWbreG
WKZDDXfojtBuS5zYZD9OCWhlHQ05d5zjKmhaU3njoIqBfHGkjw+rhWT2Gwx6DVslX1ZksyZrFYjV
6Is8L/sP2eI3pkgNB6nWzkkpl/kdwGN5+9BA7KDPbPPFxS2m0RX1CND4WDjucZDoKk/3TMv1OQCF
HpQ/XBb9W63f+weKL7o/FVSpztJDSbq1F+Kq+mrT/M2yX3DhDN7uw+m0PHI9n5D0BAYTCg2++zss
hpT2zQQBEW0vYnj+eTz6Z0zPAvmskIXaIpw02HT0JqNEL99UJZmE3FWzJhNZ7E2CuZ1K7IEYifYE
svVDbnKu26EysIP0HT8/nBzFVyGzQH7R+Li2IHXuY0MnBE+o7qf+QQPYdXCIC7nYoXI5apYEpP9n
eGZRQXSl8oPYL/W6SC0a0y5++UII8iu0iXrIRbeFj0CzDGZ3vbizG6e1HsavPx2p/c9+oucjaOSj
iRymsdicnCxFRTB59cmKDX5hTXtuVXEDtSt7+MFFamC14tHsZ66s/3qDU3Ci2+9TUrbdG59L2YwV
VEwvS/vIYqtKY43lSZe/cWmro3CO4HaW20MUvQdRZ525AWcVtQjbi5xfvG+c1mZdX73QEbiBSEC1
zrqUCqC98B3edGdT7GEeagmW65LjRCX1ZaJaepsEI/5DPWgZlFPRRWm2N6AqydxPyF1GKVOkOsRN
5yBgl5unnnw9cU9NxOUE9STxr8NoxYqRWl5WxaZEl2mFPOAjWFc0HU/Yy/94aZvQVA/h+ckrm0jg
wX85bzBwTsagc0A0hQ6brzPuxEazduSrhMVdmJaBd9pK4vOFHOzKyT3NA2BiLHS05wVpBgKve+Mt
IfwJU8Ul6YjQGFxmhQ0YN3BQ2PSq0IMCxwyWCJ71lIlO/wRxs5L4V82BtoIMIIg+meQ4hgGpO0HA
z2aP8dGLp5IQKcw/ougRHC8kJrLzX42FQm9PvXWM5eh7BRC8L4bX0xFnuXvf7XYN7OqGwNN857Nj
pWB03PaT4PBNf1gLzC21hnUiliq4j61BovxZpG5idiBX4aTudXuyuldIo4nAxFqAM2DK218RDqva
CCGYirkyb/OjYzES/P268v8FNnaAznGSXZ81XQo422fX7DKLPNfAlmtvEKYE2XN9D3EM5DV5r+vu
0bsvz7M7EgaK+Lf75zOh91nYEXJuo7wyMfJtOGMe02VTDkqj/A+43FQBojYfDby/tbgp6IaoxwkR
eaE2JuH+96ivyRVWi0yXagvEBxjF/CB3MR015SN9TdOGoBywiWOiY/AyPgWoIus8UscITJKfSWmi
m/ERZYOjOZ0MOTEUZqKfEDHSdpLMIkbbsfbwYNgA/XQDPBHErGZ3WYWxgjEtJgmAMQkq6gFO99gQ
05L34Fc2LfKU/no0Ry8eduNulJOdNSVn19mvJanWS2/9ZJLxC5/AJx9c3eOZ/XWWarnkFD6+De6s
s7RAUJh+kquLJ6PSLYWK4P6yMJcsccrAe4Vo7aoBT3nTvNylA5HONOirVNESiHohXl8rRdzCi6Fa
F/zoEENzhNlJejHMtvrWdWtGjXetqwAEcObfgNrfZ4CYy2tPk6X+5rVmezIwWrhUJwy6yCapgTf7
dhaPSWPKFT24RW9CY9KFRl9tRJ5eMfP965Ls0E/3F43oxmdDpnyM8kBdF1YPCyDoeeKhI3G63Qqn
laRfs/H3m4hpHUfqtaW+/Pr6MJFNpFZL94Sb6yAjlM+3I3QBStySg9FYaw7oTHcbyN8uSDnp0AsU
IcROttDcRhXwFKhWxshzDX+qv0nnZMiyXrGCq6FHnBWobCnd5Dr7u53wRIs+ikaw0UY9hOJjw6wY
2A1req0H8rdS4k8hfkK4sX/9QHpx2S42TpII/y49BM/jvNMcLmfCByyI+h+r0g2yg6CRsBeZhjyn
NB2p5sphz5qqpAk2zCw2uUiA2sYP+eySu6H4Rj9JK6x0LN/b4gpNxRvHrcXriR2gz44h2HbaZigj
7JB0H05KTmKh4fuTmQuECwjmQFXsingfyZATWLRSkYw8ovZXwJByb8ntsCRs6KPNxsNmJkP5Evtd
BSzIVKqsoDvr+MgU5j+iOFLbcn1WMF8B2RFioQXKnzW8oAauTlAjFodKwBcmHTh0blpi9FPAbuex
VaZYbBOEtp4wLfR6OeXrN6zHabDIvP+sZIQ7wTfhEu86qRtN2Y4jvcWvqVEiO45MMfG2Q+4Y/T1V
Zz8ZCK1n32Pya5ON5Y0ip+PDfZpOxQxNjNQVIFNAhTisDPhEnkZ1ImZYkGxr/mFWtxGEOg8Rk1Yw
CKIV4sU5hxszUX/Ayt7BFFfKAOjCAcd8BsGPgaks0UrBRQKlDgz7q52vilYfEhe73m6xshipAqrk
P7K/dNz3VRxehvWi2Lds/Ds0EG1683ErtHsDFDRISD5U0SslNsYExAvHl4rwkobU12dEhjXsIbQt
3IJb4LhRRJpj9QiVdSprmQJJ0fb3K3KU1sDYmufe/wvHgaFDU3+yIpZSICnzEW0GRwjMgArjYals
LeQlBpaIVtiTH6y555Vj5yMyGNT69T9CqH8YW1NavWgJd4+yYnKLYNszUQVkJMRMbHittDQea3JN
BsW7DipzU5F5shT3cT/vzASwy9yNhuBeBuq54A+K7zDYgQz01AKnOPotBjMuW2MMPzPQGo1F4wWm
rm5etfXi0Ub9/ZhObQthJZfjoV0LA8zfO03l57TT8P/QVma209yj3sFrQqyp5y8qjGE8Ig4cqSMF
01u5+3xViUD1wLqaw1ZTaM7zK/rTWXLTsXGI5W5Wwkekln2uIrsa2iKmdxDut5dpjTuIBWl63hLI
de+HpTCUYjcCXhToICgJ28aQD0Vxp3of4P2SwkBtOHlfvwlcL6IxBPmZRZXGlBFrdvlWj+YmcLsN
bWO0K9Vek7Vd3ret8CNfeYu1GzpqJsOZ2aXKfluQN8xk/G3Tp+P8hylNVzqWOqVNaeMq7a17NuaH
UM+mJQ1xavB6T3DkAy/lKuCWG0gz2vFxdEzql19fmUc8azD5Y3TXnjrvr27zlwG4n1Z8nFF2jdhV
XKBJXSrdZqJqKhT94aIOJDTEmvHTa/1l1jqPyPUWvdXeSklu537bx/T1BhNJVKpRQjpfP7c0f9Sm
O4mmCnXTOw5bejkb24TeVhIT6YkyjkPLCxDlQzEBZQ1trMcCPBSbqC0/vVOVphdYYtrGzAhq+Qvt
x35sKsL4oi45TNxTvTtJGFokatlkGtZYOSGxap3oPLJFtOUNc83dHafwYw419l3RgLC+wIMyTDjf
o3PZ+Tfv/BmN3LbFVMJ8UMa6vLF1U2cVOqMcDVYfjSYxL7vEHg7YOjtPbgLVsjp5zF3EsMGDjvHW
zBwIv+F091dZ3bM21tRC/T0VH/TimIgphrWjMhaqUwqxXs29ROJvwmn4zCoqqjVtbHGxjuv3VzWx
UlGNAsGhCEidqy9S8pymSvLon0GOVNc0lVRzYE0/IQGPHkgy9xbRVS/UUeGuHFod9tWzwhi1fnhr
IinyXGoedz5HGlctjtAOHSx3+Yn+vjeCbwj9W6mXGUrD0jV1giZsc4iF13QPjIX2QkpiESKhxb0n
kVVDeTAlNI8q9tirXMiyJamoTgNZy0SGAz8Q3F9bOO8QJ/fCpADTvSws7Qm4N0UK+NU43cAz2ZEa
IpsEdqmcPKMJ9gQIdpGDQsqtEn0R17DObIYe1So7llnW6qn1wlTHciTkUgztgof1cyACTCbN82Je
bF1Ci/oK2mwLOuVhgTRq7YIQSjMWb2WHF9QHWd7ultz9RcKRxU2VbtS9fIOBZoYHviNc4B+ytzHZ
gVpuqv/3PoTXNUvTK/nCAXQvYI886BWOeboFjVPYscfau7yfpQOcqZq06C0tAxrJs1mSt5+OBwB9
cmFP1UqT6IUiVtrantJL67IXa6IkCk3lh+euLI00Qg5xfxH07bEyU2kZzVMKR/CWwmkP7yhbwuiO
fOCIN3COfKbMZfOD1lGStWxUrB+PtnYu6YRThyLqnhB2vlX10dALvX+lMWwrE+Fiu9yrqPRLO8M8
Hsoh4rYxM6PXUvYYqYMawi15PLr8JBGYC8vH2tggLr0i7rQU55H03uhXUDdBYQITVCJwvFJkeCWd
ncPYgMdQ0pI0rH3V2sgURcetE0u4bJNMwz+nWwsVC/1Fjyw7LkV/yFVVFmXLYHog3hPMgr5fsTzx
B8N9Y1bctjvIOyN0IA8FnSkxOJ4mJ/1n0WHvhYXsuQw9VlRI3hWQYjDb9NHk4e3wWyq+UHqRgEnq
HL44a4XqAvzw3/2t1x/2WzpZWSEG5F7mZKuCDBgVy1XN5RTXaqtxc8RMhW3Tw//pGfzj8+5kqYUJ
OVur0qeKk9oRT6Mib489e21WTZ/eeZZJfcbTRgY35PdWT7aoDmttKiLVn+TEwj4gc8ZdS6i+wStB
earj2Y5AlpR7z2zfnW9ExESeGZZJtxqNCdNr1EX5WLSKLcGqbgQHVwT8nMsSCyvug4T2IlwPiORZ
6770jwzcem5nhuCx2N8BO4a4jIRdGmD5LRn3PEsOzmrt9e2+oydpAdxsGm/8AjKg+kK9oDVqEY+l
HjPqftxm5MyQ3nrfYwpik8gWSVB98b5QJHZZFBcv+st52N3p/lHyAE70HL2qnCPxLpvQJsc3sNwt
xx5G+NippMqO19fxWnmU8kHKkGiNjWbw+13PPo7hllXWiWlxcZ1IarfFhzSQAbJjCLRwpiErIbmq
hvMVXecxMG9aypqqqCxGCB/vBBVMX0tC973v1yzIc+DZqLvmvy7BKz8kT+h5TOdIaqr7k5aAjggd
hE5YDxoStWcGv0q3mmRh6FDvGlxNukt61i3JBtdaAnbl9f0uR/5dkWT3rZ4ftSNDi4Z7yMuIe/Is
jIYlCn13jHR23xJf5/sAsdrtOMhyd8f+b7sKeRW52b/R3DBxq9O6pqAeln4XtcTfIKk9tAM7w1cz
//P8RLLeAww6D7XlRBewCW8atEPN9z0QgR9PpCm9+8FSyRKQc5jO6pMZ1/M2dzHGdb6ozmfVK6ha
9TeH4L01YZ5ftjFdzl2Asv089oVJcApWsTkCsOrMjUbiEdkefjprvkLYri5OjbLwSSrX5px1WyAD
hNilLmIgTaGmjlPC3sZYC/8qHwtdd3JLolEIoguUz9pjgOLa7aCwGKf++obS1+JSnmeaJEvkO19K
92Ydpe/lOU+ZSLs+nUN/JTJ1S8yKSMTEM7r3LlbDVpsCr1b3xeqnSBNL9HplakAl6/9yWLXwumuI
oOnbiyX6BAXNhETX+5+Pj2TbpQHqqkD0Dk0a/lGRBbZ4ZhTfxSnTrky76KFiVtjVriWk6KwhxMeD
Ixsrpf0oe0C5o8uP/HJpFZ65rNledyuIxPFujQTtz5NXWyDLzNX17DgaMQlE6Ai72XvgixkBhWrw
6eWRy0Y9dLQBW0XZRT/J2HAhbQsnAp56swGJZ3zpfa3nHmK28Tdk6jPyViYLxl9EW5spi1CFumEF
s/0zVVyQzAKxOyx7ER3P0256STDbxTsfO5kfUykeTc56wcVPwc9jbUoDpv5Hu1VAaq3ciWUMgnrC
YqjKntG6WO9IH0kiIaLpBQAgwgsjrPQ2wKWUkuijDQJYunRZi1B1BrbOXMA7flkH+Etwceg8juTO
fPoHVjMl8lL2v3le0qtpyJT1RHUdfq8hCiV+6gDTYfSCr0hPP2c1NJk9m5jGqdhCq53P8GIymrIz
6UA3sV4MQKTrU+0v/8uoT6NTsu5wgVdBzx22nt3m/nJx55AAmoPns7kPEMGKxPfAXuXVnUQBv+Yt
cOvQTOSbxmPW6KNLHZGTUdj8zNfM5phCX+5pgnydhqFs6nP0KN1rW16CXAEWNT+7CpRH0msy7Ee0
Y/BHJxj8Z+Td4ZqvToY/Yg5Y7LbumZAWBEfO0WMt+OFZ12fnh5wkvTuhkx1kd6enGwC0I3mKDpXE
MI7Pc46Zeymja2bU1AqyWnQb+qOYTvCOpIkhNYUGB0957zlk4EbzNJFGLBmPypl8myc+xHeYWIAQ
bHkZ1sd4gTklx68+5Zdv1tRGk8I7GDQ/7Zyf9+dzdX7+QvkwDX+NqV6Aw+7LGmLN9LEzOPDVZC6g
RhiUDHrs53LiA3EBctAljz1UePCT8+ykrAoZXvL9/815YgNgRvaMIcu20pLftQX+CjyEDql7s51O
4Zj3LEX4Fz71S7Sha5O9Ztg2HtY1Lwifa+vaif++KYUYZMaXqGGCONnf9tHopCL6YQsS1Ct5IfHo
oxTBn+2KVYVp4KTlV4RHB2CC6u8ric1r++V4eODaea15Rv061GCUhVk3VVS8QI5ZyuaT6qqMIjuR
eeVmyPsmi5Ufujrs006BvQR+3SWol1SsvaSOS0f2pr+XZvDAI6QtsW5SO6ymYVdq1SKR83j28ZT1
FPmFHVrygwMtDBQvp0dsSuX300AXe1DolHqmKDjgAu6Tibl5yPW9ONrpxR6glqnYMDqXXdjic+we
OwsLZMeoQcfqAzBaAXgTccoyZZhPyiUdVMSiHzyOxw37nW1OxzRtdOq7tGVsiYfUpJCn/xtFB4XX
GMtrcs/4lTZXdZOyFslxTWGun0H6IOpAWfrsBGSKeS8N26Hc3MSoXVeG5+NptXdOHv62drrCAHtK
XiM0Jvg+YCbgBj8nQ0B19Fc9Ri1aoELFSNeY60zr2dBemvGbK55wowS4LChuEfNQVLT9fMq2yy+K
uLxyXt/+/2AbNBnP8S+DUp7aKhgUgXNw7MZvWHLj/h9lULCwrmK0YrQYHCQp+Ql5zAr+UAFR9RMn
ydpnlOTf7DXTjb6jEpRRnogJhQR+nPiB3+h6oYtbfiCdfw72mRTxFJJci4BBQjbCzPfFXPv6PTZ6
50GR2Qhmfn39hhHsaZpsbwZ0VGas8y/rFcOkAWGvdyhRPueqlGjxS7MFhyjLEJC3s5BT9qEJVvzO
AA/DjQCmT7VsYT3miby8sNmtH+FKqGMO/dqHsUOIlv3mQW00azZx/EehL9vi0KyxqbSpJxXD+g7S
TkvmJ0k+Xw+1fwbk75SJlvZJZezq8TTigp8jIrW+sgoNH2bHiek83sdvhKej5l3E0KD/BYLSL+2f
npgCO9cmU4qZbAvTaUPxxIJMWUTo922Ac44PCftlyhWrKpEG5GOAa6qpzXipLSoOqR/v2jmX0IxA
QrgfZM8vOXnvdEtxXfsH6PeqmUXs0xqTjxOWJw/POIPPm6cQv5QMKUK7P4kb3AfaLFVkbYxOfogo
vIGR2etxfH0SZsCzPjUgcGmGdomwm6xrmWocFWh3wh3YgK/RV9eJ0D01EhOn2VU7PP+RLto2j7Cb
tDHUcLgut5WzG2DqLyHSak34CjKzBT93T2GdGRB8moq3ekQQzs2VtiAY3T4PHdQGdGCfGw7jhTDK
mXNxJBSzJYlVfzYyXIm8GoJYvjlcHfZ+zUYsq4muLEZZvzhB5pDA5Tgh8A42YDOZ1GgPnCjFxhVs
oBnkBDNJTz3sdlkyxp9uCFUDWCzQBJqzNgONWtJqGApRTaD5f427V+co9ApU4O0dAplTy13UxT1u
jA8xSTAGo8iXLwis6vJvpSxf01MtBKrKil9m4aEbwKbV92A5/Q/I6Q5nKP3aDJvQlXIfo1CYjyrT
ideS+ymAPj/uz6Nz/cVrKImVoAEfYawnnDIcHMwpijELntoSl/F75vBzn+k4Gen7wHUotBwmTp+N
q2NjADWgf+5TrdlFk+DFs6z2GWA+bM172qWNzH6w90h85W9fsrRgLYrOSSqrbeZFP8DqO29q2Inl
8GVLHm1w+HpRVCgS+CrgDCmWk5T476sn29JpuDqb1Us7NL2ld2Suc0lN0KL2PVD6HbBFeGscmbOz
rFVbRx8j3Ks6glPBdt2pBYAXZX71ByCshzhKNXZ1njZ/F9hA9xEtMLCYyh3en2B2wUGOif87kgyi
bSg2KL9K+DoYiTggd/O5xba1kx9ICcQ4aknApN4PlLDOpCVG4LzRIBd0Zc71lQgnqhcLo12aQxgj
Yie6kPLbizFnuGdH7tDoFyCoBt3hS6gEYQv4ngaM1yQCPSclG62nH44/F6v6bmv+65B9LVYHHQjk
uraTSMrYV41eDAdeM4GlKH0l7peB5aO0Jwv1Aqw0GQQZ1P5jmrkytugo0swoTYnHdlX+AEET6Fn3
6MfeN1rbRKV0w72WUXR5uIjAj7dp7At7Uf3Yq4Z/NpIuSAa3jEu7MRzn7o9zwuSpX7WZI8RqfsRp
BZoARvrmGc+yaV154eTx0uW4WFTlEZJ3oJHGSeS+B6MqWKfugQfWDa5BMIUPbRXXwx96SX8HRxrb
TbQMcVYrLBG2qaT2fdS78c64bH7YY6dhQBF2kSbVPqYfy69vLzIL0plPEhhcnvQd6ahQ1OdSBseE
MYTgyhTjF38zjMoBbRcaUdw+x2dm7+r5podE4tXcYA3LUOVHm5L+XYdLwO7CopCjc7c6jrsR18Ff
k/BvKmG6MYV048JkCQX4TB890U9WOHeqXHEYRcylyKbeD5dZLlmW8mERF5QO4knR0+AkNp0YClqY
C9pqtRNPdnpC6GLMkLkufIP+mt3RpCVwQW9S0ozsR3maNjr5mSp5LCnsHqj/ic9xiAwmzoynEqFR
nS0LXP4GDLRkBUbb5r8IH5MPeQa89cqVlTdmApA/CIVNmesiRjwAix+WEC9E3wBnlQidVsk/W19O
8cMgldXlMWBcM1bY501RaiprktXwrxW3txkfgQytkRwlNHdhbtkiv/46SLfVF0e9O6tAuSSKdhQm
dRFx2mR+WsGqOirec4sl7vkk9tPBV7oXx2g0vVXHlaedOpSIwEkdX8pp/tTzsUegg7e0tIqKuRcI
HIqoH2g6vbJj+jM6TcDo5wg6zFOGvK7qfhN7uhkt6Fe71CtmZSbKt7bUsVY6dZqjY5sToF/LkQJd
CQu0qXg5XYEUneUBn94iPcMXXlA4T7zxrjBw1Km/aodt/rhJF59dR5zTeIYTbxYMWBORvXoHjQZc
1u4KfyMGUBRfzhEP+Ud/ac/zAbjKN4JP0ojhILDiyuyvSXWM1Mr+AA+7tMamBWL6a1/k9vjeIXCZ
C2p1MrdQCIE55jigZ3NB5EshK/xWDYob84lCcThgdQAZSjXXEcPY3sifqomlVtW64o0Ppx9O4Vx7
Dp5wJ0h/j1qGDf+dLNFoFDVvgjXlh5QZAlHvYgNaeXw+n6+LbSTCtec3whMQZcg6/UjlGn8UAyKr
26QHRy9A1VyXidIQ6jaCX6fOwIH8hJRJhUwbpD0Y5vPmEJGIbmbzsYJRD9E/Y2Zhpz2bxoaL8/ca
M+gR1WW3wDRKxvlom54LrX8InhEzfKFdBksZt5N7co2p+TfNUcwk3lFU26xyWM2n8uH0CiQtpk9T
452EzZ2GkjDk1aA5DiHbW2qk3j2Sziq3tIEVIr+m50t84/4F5kzuoFUdKPclkKoZaa70odx/Q+t6
7WrkjUClfeQKDHNa0Z8yRNzDyI621DnO/LzWQcrk5KnKOUZydos405rNiNL5KOsG5OawPJ574O5k
f20VO+ra8l4RKnlZNPJIiWxy93cEbLVVT5eHBVJnQlYO3HCcyfSh5CnXfqaNJS/wRD3Xa+2xy0ug
9h56jNdg63odiXAV56swBCaPASH2z+AkQIF6DVARh5cksyT+thDdlDdDkskvJrqiJ95KL10mXUVJ
iem1YZCUqrTW4dcanscYFgu055nN4uH243ZgP4esygiCm4it22PoqoomIsRsliRuTax5eZuxCnSZ
hI1IWrWen7vTazkpIHI+y5KwTf3GQe6lM+R5e8+6XxbDnuGk7FiJ3Rzb04pRiMmGCOYawjGorCMh
vu2Syz45P8e543JNsI6jW/obo8oHG5iUrI1xFmGOv8MGWaHkr87MW/TBPT/Gm98YZ0rKFlKc/Eei
5QOU67Q8/F5x8ii6ReQ86CKjnTNVYjvZZ0qLoywXuWYliEi2Bg4FpDZ2Cfn5XVMZfuIuELttgyFE
nN2RJYIcvX5hqh++Hrje5IJI4XoqhYHrySd49Gb6YfEmA3NhBj9reV55hCPVA7XKHLnOs+sapgMT
eHxBCRnDkWhnC/q/ceEiOavF8iDpQUE3I3qsCL5hifWCWAHHbKmAQL7rSkOqlLYpcH8Y22zuMt3H
iANADtOoCngXMYqH8bHUT6PkG97mZNhpUEaABR7HZdTHE5tuCdVaHGBuK2Tj7HrgInLtLC+QL8F0
rfZmmFcxiwZh95oE6KqOlENENf1J6VWTy8IIdzgLA08ws8c7NRkvkIjlp5Z4bwaomZ9dPGEG8tNr
70ygabk/xHMiT9wCHWgTZ6LaqkKAFvz5g1yRdZ4tkVwkFnx1x8TxwnBmdUnb/5zQ1UIgKwVM/IbY
ucyFkowEYDvctXs5iDEn6KZ6hIUgA6MvsHPEfW6lobZw/UcdjQ63lQyS98+NJsi4y0oKa6Th7d5A
MnXA2SKH1flIZ5D3Fd523Lltv/lS4uR9/h37CcNfCCrcymRLs+N/nsMImjLMjySh7a4Nc70gPx8M
cRJe6Ea+qAHRNcjQoF4KdP5IGNq5RO79bPAGLDlN+utNVXS/+yDBPdqfLM85ls0U5ZvKFHkjFfZH
9RCH1MRPAjEFvjoFgQVmZR29J9EYmEYj+h2qoQF+sUB58XOUmIETRAnji6FhqjnHnVgIHIpBge3y
qR3IJwHXuef9Ond1AnUQHOkHSLMkDBNwf1ZgBDHRyZmOHJSd8qllx9RDV7KftVlIEEsufk/hrtxL
cJJ8fFp4AfGCK2Y4+jYMjZQAlQrh2/XXvd5SLn41v2Xf0Xh4qTf6MT1cSIIUZohDpyOLnOqTRi7Y
F+7RfvhnUKgV67s+gV8fAhTDNNjElwzrIR6xpDuOypqxTEt2/wy1/t7oBEFYaUFQ5a3EEYgomBKI
UOnD5GAUx3G5ukJ4OoGBF2VhUiRoB9UYaCkei4plpsn5u96vrVnCLGOcsjlWl6MGSiJnzdTGjEdw
gifDij7iBV3rMcovI/K6BawtSMrvW0cTAtV4FJN/b0tCwNJRwyWHL5ZtH470tdJ3IsjBNnI2XSIi
otAFFnSm8XllptWGgfNhbGPQviHUBNv0Xzb31wn45gKcXhLsiMkAxSPhsYT++wWJAzKAWNfACYeH
X8IrBdxnpqXAqvtEPxs1RjnYgmajJ1qXC0Z9J+cPhTMNckGqh6Yq/nGmjnGQiQuxx9X5g1T5KWYa
jUOmMSnniLHyNu8Y9jzh/cIbbOcZ0AVwKBl/FPEfBtX7QAv0Pc/DkoDUEBaOxGmxEKheez5279u/
HJ1YbF8Pvt3u6Y3pqbpMgv8X51c/juRnfOE9riKLDwQ7AHc2PRE4OrH4hZJteHGKhbgCXQoQvtyZ
4Unw38F4p9fbc9L1aXfFzj9WlNtxUeaGgz3fbnw4gYLQRqtDbdxQCTUd1aMD7EwTlyRH2ydNe3Mt
dk/YcRKO3jeZ2z2CDWXtXa8feeRvquEsrwl9qA6K4xwiNCX9YwsXk+zWMR5u6aYD8TDl5TvUWLxm
YPC3337WZtJE0VICb5Qldi37X3YuLkL3S2ZuS1OYMPGSEVnzbRJFKxjLmI9G8XCvD2jSVXSxWJ/L
BXvO3zcuMKpr6Jc82nd/FVi5nn5MhZthxAIAsaPvZiM7jabVwQLZ32sr1eGZ18qu4mSnp0MOMfje
cxUWL9lCIR6v6pGXWyVGyj9ma5JAk4qDjaeKww40gvaj4o44Q5jaxmN2T1aD4W3Foaj5CFJRkx/n
PEiBSwn4DEnMdRzNbcEC4ngAAE385MwGB+UvTbWv+4KIl7+IXaH0Gma0hWg4XxKlrdBld7op7BBz
AjBepp3HKxnMg319UdE6cFVhMgYBND97+3X9nqclFLG/e5arZ0hpM4NmNjuIO8FEAKSSVqGnP+D+
/UnLdNG8nNVlnRxVx/z57MhosdIdA5OZHfqUUhAcmt69bZOq1tGIMVnP5/qBpLPn6juQV5mN2I1D
/iQyzpyTcTYQN4OHPOcg6pLhu9YDrSojTBVksofjDhwBI2gguTuffKErPv3b0Th4v//y9jMBS50G
w2tVGEfJKBk5gewGXns8e0GQSb2o3VadGNZuBlm5DAviBOuFqYmklj0OTzuj88yI8L7gXfWOdM8H
t6wYBdQPBDiuDs1bLC2DArCV+VK4U/L5uUqmnaCk6j9/FCZwn+uDmpt4OOiy0i9tZhRWWqmk+IiQ
6Q0s5Mdf+2uHlxz+5R6/kJaa9ChgqMmvjhE41pvqvfKIAU3bXxWOTrp3plN9R+PruSh8FZ1yd/FC
ua9JigeAZAfH2oBM1fe0qb1rLljPOULEasUw5rgtvj58eMwFCYllkLs39Alzz+QDdXWJDHAIKv1d
oStxh3zdQwXuhyCwdCw5sFwXx0GOywdEXuCu6LOQNFTGDsU+nwS9jmwaQJ5BK5tMvvY8vKqyZua9
OZuqyPm+G1LEOm68nMrc1jfijZ/SGViFNryDDddgy1jjcX1gcEinEF6ao0FKis9SDGmUWegh9qag
fkVj8f25zG9D8nVKp2qqLVcuTmtKfgt3Nf1qsm1wlxhWErCOGQgxwqMRZgf+dhuKJBENZo5FPLeT
VXPGxWok6UEGYT+kn7r89//z48GPPd6XjF4owbaxu9yWWkSXkM6Qp1oE/CeerI4a+hPvwk0VLe2U
ThX0QINzUD+vNSBegoWqmrBcL10ZmmpWQLtsY+4afF8fcOgp5wa2OmzXqGmg1R0CM//IsE3TDUu1
7FZsPAL0W/ievy3D8fNFy1T/bWvQmM7qwZjo+i4GyZCeQzHR+CbmblUcubQCErFVvQA6rgjG+q0S
wzhieQxmIKZcPYJm4/axaomHK4nH9nwrVoukLCa+TrXTJVXKB6oTSOwVIMQwGMJACwYC9TUdWtdT
PIP2+fEExr499dr5D6YdFZB0GxGNvlbzmTRobWnB1BAJKFOGy+23wq7sg544bRoYVbXV0QRfE7Zb
v9BgMJethvxaRvoJ4QDPu7xm4HmYTGjrSZeMl6S9c3KkyqVw47gym0mOsAcBV7Vyekh8Vnd5gFB4
9JELZzZF5uxTrE6HseDth3C+h7Z3FM8n4/MAaYqQe8s9x5FCCDmrEjWeu+1CLyhcnwtCHe5duAoZ
ii2Zbv3oqqxpr7SrTuanJmzqkAgo63Ui00zMESiahCziEyV+jtnFERO4LynHUK24T1LftPZbSP+K
NcAzpIHmz6d6HQAsuN0MNrqqIl+EfahZpJuMvoZl1JftPouUIy7UhqZmOrY1ex454yhmqnM/rW/Y
NhG2mO+5N/Y4BmuVDwEzmD+wB0i0lq5P8MgUPbiWe4BGzs6KA5INSyxhhpQTfaw6obNHYMPaTL/F
iYud9a69QPGtnfwA9lExrT05NgO/P/HkubKm7goYDk7MUWBK+/Y8eNZBAf65sslrvaQ4syDyLm81
Lpy77Ao77Te8n7HBzZZQLlG+JRY7h6QY+sMrwTZFkgdNV+DVMtPrLNin+1O47wTi5oTjWyfpOcvP
u8JJTet+tz3d5lZPkkj3x6z8ymkMhUnpHLU6JqYR+NQlwpguc5JFp5T3LqqM3uUMtJOr/+iayx4D
wZbhIrmKz+GJErKxsYFnXq6TrVVLmslUt356567iFru9luTws5rJdzCiT01QsApta7sSLR+VBSDT
NDa7JblMh0jkfyhYzhOCjeaGXn2dhQUPuTsl0LkOMNKbaTpIZaUk4CbbgR4LKNacwG6qdKi+oW2q
9DGutpvuqM3kR+ca2trRYaH+C89E5/7zS6S9HJlxGJYYH0qeLKJXg7YPL7zUuxGmfxXjuAFwP3LY
Zehl1R/LGlIMSlQg2QB34JIg+QfemUxEFvh2HjZzNUUHY+f6BKs9ulx65cCqoonRfGa4Y+heNPaK
Ckvj+M1snihkeLY2eq2eURHrin+cjB8HQEIdBwolVUyQSua9SmjBJehxp/9C2g4t1Mrauc28RmFi
YvqWWQmfdiZYHLn+Mn48kIRhkR9A3OJr2T0cyK65RWTwVvSVWbDfMWsk0cuUBB7cJcbG8c3jetGQ
qW5f1gIUBxNp0bXInqxgPESbGuPTCvFANOy+Ryy7FHiP8gz7YqiIKm3ZwYsXA/DApWXiBD5YreVD
1Gm0XP2IwqU+UCNBQ4uVyIrLwOfl5ub5+JlXjCO7pU7k52TaiCztzuvsbgexc5sZTP22gJ74yJ3q
RhFZnH7A48HWJSdAOj+UX+79sRGSFZG942NGDtGuG3WxaGyuEt86MKjUgFeX4x6xjwKfOB90MJgE
PmoKlUnvpvFgJxhVAvYCk7lBQ/5vQLWJ2Ve2SrPe0Jhr8lBONxkeZXkHH0gFbsVbOspPZTjeoKwX
jLecAcK4AeI91qOFVPDIj4IayLuEkKmJLMeoRXzfQuxMTtZ9IVtGAx/Clam9E4gqmCwJSw3v2Mwx
Wbap11BGRpOa1jiW59EGFzTGVOU9Xp4RYYKpt6V4COXU1UZqiTcYn3J+KXsiXXbjuo5DAviOEbJk
1bDwDsEKn1TNtDXtR9lPMI7vrA4e1pEEJk4sXobzASvvdqbdyvmmGd+zwmq7iSrn/Ec1u3CnK9Ur
OrVLYl444OI1KYqxVhRqK8tz1N3h12BU03pgJU4vVU83O5y2X9fe+msnWN1uGiu9//rPiwW7dkqm
QJVOaz33jUaUn3SBXiqRWQx9GEU9gZBwie10UA4DTN9WqxIgDyuO4FtPU8/YH68+YFJdtQxajF0e
tFlea/La6VcAfR6NO4rLk6hqPNuYoJLLBIW6AydUADf8XdFszteKc1w2aISCQ0hOdcIXMA9+BjUx
M2gVMM6bQifpjno7iFesDEKiCO/IugKmSZHYmFSKyootyteGw2aoKTlMvZKtMuyBHKi4KLgsApEd
ldKepBFzlwqewGzhZQPIuLNbonGXSFyrLY6/quU0gpWZrOxGKbO2ahuUQmBuM9WCJ3wiuky7Xr8w
ZRoiK+cHt8Wti6ADPRQrl4UG99ovbEZbFtZkYhyRleuKjUGGGIvlCZs0488aWj7ee5DCsa2KvOOq
1LFEq7I/5p6oWNlDXPJHGd4RRMw1e2QeA6SbCx4ZiVIzzHvF5Rul/cCFqeWMXmT14F4kGraYmRf1
bd6YfoKtf9ORW+BIPUP4Iu7nuqVDycDnHmv7P8cPJZ5tlCCVyVBv9cHPr7lkIFCgYAMCzFrfm2c0
cdWlc3uvkCV62Evmb4cwB+x7eWFb/mQ6WolzqzWaRfCQ+a1YF5FVSgLDeik8JKT26BYwzZ+5f59T
oaZ2gLPS2p4eWiAVzOnNo+4VpxSo7MNWIo2RUi5Hck/3QxxRYogFL8hzPOjQ2Ev3/IxOY+3y+KKu
NCAh9O1AHfm2wG+tu2W2id1fIgFcWjz2t/x7ygHmReRN/br/L+U/zdvjrR7dz3uKOxsmI5Ga3u7a
UTnpj7zMI4FiZr4E5KYHwGTakZC2rE2ZqbBh02GSGZEByVaYpcrNQh92jNDi7TYIeKXtyKq0bCNP
bOHBR3VpeKepUs/AN043xRcK0T3qhGCQuFQvgPqLLR9idL/nb3rg2kW6kfA2Wt2cJxtZbXQvEFqQ
Jaheb3pvvPDiAwi7l2t4OnHWAA8oTw7CHm1BmAJ+bjq2h4EqwNYUNp3RxklGabUxHPryNgyFxXxz
uRZxvt3oz3IE7H9jiAm3lQFl2xYNab2Ez/HLTxe3EgDVspVo8rbyiu0SjosnPpUBmWhzA8jBTMn9
v861rTQETWREuzHX/F0nzXJVoHtSiv1xw9uL3OXAPM25FFA5yJ2jnTFiC4ijKYt7YpwL4xGkJT3F
ZpnctHfKMEAbQOPXhnALLZZvaDHcHEqabOby312QK5N6YS0BzZfP4HZ4SUZNX2DjWX7Tvd9KRICa
/wL7nIuL3WLliURGEOMsoA/nFQqgX+G1HbnkYvnlvi5br1ClVdAdSd6Y8vKUwEj7Q37f4sZs/9J8
pXk25+l/tVynW260Tx16vM7ZJtP+sfxGopNqzU3DsB9PrPYPwD9LxztSQSViaJfg08Z1X1YAs9Xh
GLz1PgNRitE74xlytD3DeuQ2buZ/aVefiC0FOCpGXOkKa6o5KHFuRfCNwp6ABtPonGyMeliqn4dw
CypRnw6h3bNlj6R6OS/IRe9fNmF+AO6GUfkA3VgmTpdXPaod0gCDf/mw9qv1q6HYeFwc7kxaPbE4
+MpZAGRZST+r+xYhYSiSLIqUp9Hmr1zAkZRGZ5m7yMIOzW367CZKQ3RwesOr1NkQoIg2dF3EiCCT
6uNmNI0FTWUWPByTlWRNMNOOeTw2qGETgBdTsXTOq+59cvGFzf8sYnwDYZChxhnU+ZzteWdnOOPK
6+o5RUwlykiXXF19VtCaOXMEoICflOng0dS35kztaCAwEFFiCmpBSUmllcMwU9W7J11htbcAqgeW
/s+wZTgVjGfy86ajiRz4ZmLfEoiNDmThkAqmf5Hxksp0xTy9zt1700vqbJmhcsZvydqnfePYC7xr
Y0M2Wp+UrX+ujKReS+JwV5J62snkWXZdn77OJeICSoDdfbLBK8DqgrA//mUlpdHBzBjjQYecFemB
8LA8frNCcMwUiihdtFMacH307wYsvWeIJDv0ItfuN05RhdCYpOs43abvwOvzs80YDJmCnguJRJcJ
g228AeV/biXCZJeszmygz6IdRsBGtu+iH0vtHSZ0o2tAz6sguuA8S3iVBTcmUGdLfz6exMI1MgjG
jCHh182a3qDoW2lFMlbnqeJSlumaG3aeImztaat93rcfDUXRnLD5Hq1f30anVXMr1OveeL/9sAUA
AOypbEiZZ4vIII1enE5Bk5koJEDskyUpOBwNZ7jwKBcR5W5sxzQ3qZbQakJy69acWUCyqXVgtmAM
nlpJ61zUvYVtXnU28RUtgxil+l1wCJhrGBjDeeS0s83ovTXkVf5HMpqIaqbVPKl7Y7XQhrcOPNCW
7EAW5Ed3KrxjqUCS96PDtfVlUlgFOPBnfsgd6N/nk12I6N8NDJiqWCe18NKILo+ni9wyecZKErfE
2Ang3IUJ/bB2CviiGikRnvnGxySvfLMui9k2wnHQPPDPl95BsOBW1mF67eY9fbXsM0bnxbpaAXaQ
uoLP5ahza8v3kLdRvrbh+x5pYlCYjo77czSAAh8HBH1oCyCDvBiKCCrpWQsjuHit9q/rP9yeq8Uu
wiwZ9X6wghWr+aYty8MMYaDunci24UzKQdkrflZ/wFOLbELh4OOvOGB+lu8btbMnLLgz5kwipWVl
pmCFMYFL2IQN9utBpyZW+hPOVnRLwb3Pvb6lVmAEZFme6NBgCtuLkscqIxZ+Ale/qa733dK6yWrV
AFqB3IUx8MycKaueOrlzRj/YLkvFMdzeIOimCe0MuP6rh2+iUW5NDlam1qMM0hjuAthVFZFEu81U
7HdKXuRVbf7B0Fwz6tYG4tsCq14mbuvhvDh4fKCv/ExRzwxSrWYLuMHWcPJFUfTpeHuF2CGO3pZU
6sfw/CmqS96YTfqAwHVQjZMirXJtSAswTw5E79JWbpV4ohSyI8hQSCb/7grje5XBgHlOMZaNxytB
lKhEkiuiifOBnsVa/CISbed7fSS5651iXUiL8Zr5v4AWh3CHGteEiS5ubr8TCisnAN37xcJhEjSQ
SRmPm6hM9anwOfH06wo48QCmcSfnOy4rqEK+NSE9UnOUQKgPIGTgdQTN00xg7m6YkpD05/YHpMuv
IFHG8+DZ3T4BuaeRPleWOc/Dz6hksIIYX+H3Za4rZbtsFXd4y+sNyPlTszvx4ads5pd/ArbO4b0U
TG1L8g/yoKoXZ/G/f+qSA2f+Ga2b3Z3eN4ymjA2Mk8NOPGrub9zUhkNSIhOzuYxuZgeXNZAy2Wyp
ALcr1VJFSnSUPWFDtEwbgwIuquD6Az2Z89XWw08QP87fc2Jf7ITlEiFWC87aNxGhK05y6CVX/Abr
OaFJW6uM2Z7jcQEeWHnSXumTGU2az06n12Tw0dEria25I8ykUDaBuwkQUJjLyS6e/B6lBavLiQqK
PaVomoz8F321H6NPA5/XcHZaViqTLHhTfymVW00rhphqxw/cj3J8z6OEzWSeOWOBbqv2trD3PbTg
nak4FH6lp4iQXMuL5AiulSe8ptJnr+nDg7bdSfE3BRAo0s6LWXC8242oUwX8TRmlG+2E8Q/NNGzY
LGFbO3ocC4HAB6llJqNejZmC0r1yuUpKe0tg7CQsVZAr6xQ+4Eo1A/Ri5j2MU1aV5casQ4a8sk+L
GbQTdqPleVQoAoNZVTDLhaCTVVb3fG+C6tLSgXf8BhuMNQV/WcDMgMdLYRDgP6g056FNo/MCdGoF
1SsXmJ1iwS0CwiYNGPycK18aG16CjSQJXzoxaZbhvDL8mLxrPAfulnboy3ZkmiMUEMcWs3ffHgqb
yrPAtDjIhOeTJ95sXY4Cm9MsyPzPV+sBwqtUEOESeVCJweoteAJ+7fHUNlnaZDR+gDMpP8csY6B4
ArKyxBYzaMaBPkq6UciRGEpogJpDBf+Kxvgdl+lYcYNnakDozlRKSY9QU9k6wBmx0jOJaQbZhvqf
JpkaV2RMQXb+kmPv4YQhIS7lV1CtEYIPHv9l6dwFDyTgfBC9Xdn2zIImIjRqhqoLVQWlFhFxvWWy
8FK3vLa86/P/6/nZ6YLak9J9fqvu+TlpKe2uBiBpS+E5fwvTq5sydZFeZHuvoirhs0dsB3gjDlW1
l5nSHDfhGvyr6uoiLo7EadjqalvDNnA2rAtQCZB0cJbJQN9XiL0t2puWUftpgo29RpoxC/6rmmE9
erxF5ilqt9ZWgTng3O12Pl0MGIolK04mQui32OIYp8+s5KPeZmCunR7drdvtsv7qOn9nWlRXiJkp
bddR5daruNkv+JmGTscmUR/IrSc42hmoh81W4p8oWYMxerYzNqoLnxxV+0GPtrv5gPBk9tPN03i8
aPs7K/DackIs28DR705r6C01GD7IpT3wTYUcggSOmGbvKxKgD1oozsUcwiTCG0QOyu9hc/NWxBhZ
KJ3vgAytfbhBpDhLRZNLMT0SAn10i9Yg/nyT+yLPRjaOMuojOrE2iP/0ega7ECqpYO3ahh7EDPaT
H2ec+mLbpgri+ozcH9QDW42GWIPDEeD4CZ3r1Lc7zw9lwkCT9Zlob+S8CCPtgOgf2OZpdXxhoyWL
6oN7YrsfHPAbXFvsZrS31dlB+OCwFQZyUnqQIfdGQybjl+hOpERhqEsgasWtdZYZDysqveUWk7+I
6/LsU6QUjmsLvpSOjabupC690n4cwHkc8z0Fl6M8CkLwVjTZ+nwXsLiiWU5FLjlsKPEhKUm18Lnu
D6uny1PYmVeVuXLZO/EY8pTRlBc6gAp8n1FwwJp14vs9p+z5hNsEMn2q09ICS4IGCCnvQjpRtqoW
v1cEvGUx3wqJ+pA9juVPk4Cc2Al2saxSAT3LNHQufWI+IggdnhsMd6jMPbJpV//sNQZfBmTQp4e2
DboS9Y0Deeom1VyXTxnfAHX8CFUqjeSxsrL712XrxYxruovoZqAohpiUFy5vyV95/p1fI2HVh5Rq
4K1LRdszFn6ACpgMzsstgg0dHNR/gSQdlRuHIbBpdp9LW+fjfhC3xsoRYr31IHNXz/UzDgLsZtkn
yOe1vCWiYfwfYO2Di97HglQJXTTQAeZfCpQTbRiBZUSXnLuOUw5mRlbaLLyuKQMgUM2Dp2DlORso
2WfHbMjAGPty7n4TIEqQGVQS05ACQhHk2ZR2Ot/q+pKIMA0/q5qJ+FO+B6q0c+kQwLW5Y6fHjL0x
BSS7MkYZii0z3+Ik9ZPTZJS3PDEhTW7G1qXljqhbmtMOtTus3NeIa64IjsOGFKfajP61Gzyg9MFP
qPh+9T8o/iMy6eJSj7+aUF4dnoeP7Ba6CJpV7PrANVF1AC2rqpJ6c1cOlKdsAM3fB7/mViIk+ij+
AyKd9juBl8ZnTQhVjK6HG/BeaI1rymu5B2/IcHBd5VGapEc6Z/awsa663UndFc7VQhpMT6cXdcTd
rpnVRMv/SdhOEvIgig6uP8c+MpdKkzL8R4/wYWPgQNc1MVMHyFWGdY9YHDcdlGFb9uDf7RPPc0qD
yYVn1ZZYjzLRkl6kL26d6TcTcV6YcHU0bTAJ+TiNmYTVzfi/rU2oya9csiZ31Rf8B5OkSYHP09dE
ET33FzT6VPj8VWieyv59lJ2eFP9VTvQPG9r0v21yzjGtdcK5BOYrh1kspMFGjSwW9dxxbehpXc53
oKQaAMi16LD+wd0KxHYZDC7bu/LZf/x70E84561ULiIFocttN03ftZakMj1WUFmkQ+mnOVY380eH
Z5SUpb8eyPBFcxlj5TNCofbbOZ3t2hEUxkW07ySIvs3gDbMnvAJar3m6BTs32jbsEjuDimITpGaM
By+r8gP1Mt2bE20yC1KkXMqsKtnKS+nOIhckLDYjfgsxe3YZKCjyw4KxwuSy9sampEKO8PjdW73U
3wwdg1bX2Bi4fjiF0RtVgmAbEj67UtILIntV2W3HPXRiEJeofZB9BJIQrfGaHA1nZRnavYSWWarA
pgdzxwlL3EDp0cRSZ+JOYgyufq2BJJzOO2YvQb6y9orxDBm3URbcUgUHEzVzTHDDD6xBJWkIOaWq
NKUERKj3sJZLkvxB8M6E3hg1JNLvl+b4ntNN9KVYebBG12FUUxZenGpnR/AlclnVkOzaNBEs92z7
Q4bQCm+AxI2hSbbo0wXZCSGz22qluwoyfyCkut8jJzBSVFy/EJNwJ2elhuz1+gBce5FdoSq98SIM
t1pfO+kXTUp1sXLCBXsKhD0Fp2COwrRgexUPvgE+bjLlztrgHNNKeLdH2CW6MPotWAhv82ZzuWPt
INxEFEOFcArKlCWoeqiYjrbFiiGmvz+tKmlmEUoE34ljJNrkRevba38Vm7lEGts2BLOSZiPeDBNZ
+DkMGoFX4FHy7G0jXTQdI3Qixyls1Q1NiMZkYRklQ5tcwKy24OWC+OvgoW5BpRYlmIE145b/W48f
fbBJvJn5+tiUoTN+WCM74nb+gF/McwPqBDdXSj6VldWmCT+v0QbKgBsvwZuq6PRO/4Le1eTFUHb8
HEio9bnUGcA/zbn9h/uDIdMVtOHOTtEkHzQSDNvvbDfrMncP7yMnLG3JA+F0lGgx7Nlvl5/SsMSV
aSUngejpQOvZYuMGwtRd85YbaqVHxn6490dccP9rgRCUMjhh0fRFrlopaol3GCJ3PwVmcc0OfX3X
tlvmo1hRquuwecoBYwxx9o6p4ZVZL8qygEDAPHCMU2eUdmOm6B5ThM87HCB65kkykc/ffGYWuq4f
MF777pHt4qghUJwRQIHzvGM3yuBImogm+TuYM2etQTvZwy3gEIwYEVm4zxNBtQJt1Fz0Op1sEVPN
k1V2ZnVttFiCuE2aR5/Fkge93QMy6Mruh53OF9/sqTZdMKrjTBHCUxEj6yKTrcaiYEhKdDvNbP1b
0KWS9v2w6P84R7bLUT7m/KI1HTUompxm1cRH1M2vAJRF13f8dj1z6rm56Hn7s5gKL8ePu06zMrnG
oTLsVywjZtwOyoliuxOf9ELjzoEoMldLLZYyqXCwZ4WtX2JimEelJgudKi04TDo7kIIpuYnAH2kY
YiGPmd5twvBnT0EsK3QsXKhhfYmzLW3yK1tu0aXeGeJQRogqwnlkWshCSb+ZMGIP86mYbfRMEo3j
5JMXmWsBf59J+dJsyVQgWh/vjhczE6JhHpvrzr0k+nDMTRztbWVwYD9O7wavYJ1xLLEGVE6qO/Qf
al53sRMqN0aP7YOEHMzpKiPVIcX/CYkAFYTBAl4LwMLwx1baRHtD3qaNh4jgzIDerzMGRwNV2I40
YARMIL608VPQzn1O2t0W+8DgHJ+raGFLoiLLx4gtIMF1dFYNkZY2ssb9Rg34WnuHehm7SjdKwFQv
Mxwky40vo8aJU+HxlIXS4WU6NtyGvos6HJeUAr/PM6vtXfhaGVXxwZTP2kgQzLGstaG4hVbAF3fQ
H3k/vsm9gsnGrz/EDYCu0YYGdv0K3QoZRDPdOlctGSqeM9jId9gT9f7ZYNhEhzEgtTVigBg79Igs
xkArYxlvGvye8rcAUfKc3m3q9H6vU08iFZO01P9FBrMfPu2eWfMgbO4AkL61BMhiK6pwPXj2GQh0
SbVYSm5ButoaFAq4OepjQZEDAZ9ZoPwFqr0ZtslAwrtmhleAPnyjr6dJsES63YXvzptTUTwQL6LU
nc3K00muAgG5viUcJqSpJH3uhp+/OJQFA05D+jNECQIZ+Ad13E8c7w+bfEvV3qb50nePmM6VOcQQ
ivmSP+laE5nk15KnGO7hPWfqu4s6gTeN6bUHU6hTpYPBg82PNmi2FnAvYHHyb1OMJ5uiFAO+sZPc
gArJvfg0mxrGsbEdEpRt0gvOU7ltRHk1q6WGJQvXDDetnMoB2OBozJrHoFd9r0kQgr9+Hcd6svSl
Nmx377byrTRRg3JxP3h2Auhv/P7CMa79sbXA+zVLOpYq7vP9SAkOiLT0/pWExXHAyPe2Hjsf544r
sHfCy/PtZeA7hBjk+fS1JC4u25Q+C0M5MwtxHR3sfc0VWtbYIUZBhqA694Z1AFnVDAMyL5SvqRAD
TTaWlESz81GIoqbcfOt2uTb4iD/KDJrx+O8APoy+KGryMXwySmbL7K+shncU/GvLzFQyrVuUrG/A
gSC/4E2WD3mS3cTUEMr6xjm9Aiok3D/pbGX7fXEsP4KZUKiLbAqeeShbtQCODew2ujjc2Hcd0I3A
/5LEbx0lYQPyUViYUzlM1+e68JpkiaNxBLyWg4VD+M6LUB9p6LZS9+kVuBg71+cxMHH1UMnf/mBb
3Ojtq2ambZy0/DDptdMP4CKAZuteKgz9c9ezh9HKD3AVlE0BcvoQbP7SMFzvlKb2fgmbEvu4Yf6/
Rv5x1N47Ndhdd9haPUSB8ORYVtsX1wmD93heNMeahjAJjgkB1f/U3oyr0pE1UDQnn4KVhq94CJxK
pWdIwFJPnHPA9kjGSAg8sbpw97eGP1Ou5bb6V4++2ah9oboa16O/EYb+2oZFZQRdTjVLHNp0kNc6
jDZKIzmK8p5zgnkH+bLCYvxBpd0nOlD+0fUHXTbl95g9V+qFJOB9vbvjkHccEhjvDM5VJF4rwLz9
hNBrqtVAP/cpaCXJCTCXgpjmwzDQWvGBypDhqW4Ul7fx5vFewyZxbsftB2UCrXi00+aXPWu9d6If
cvJUmrCiov8X99s2JNLhSu+en+/I2sjM+lqVdHrE2GYEY++gc/LXztFScsTVfQvrBq6W3F3zJXZQ
kTzIk/Pyji5eQkzQjghupZDMNzBTyImWJXMxnqUS0/bg0DqqEyqxtswFTuxrbHs1CLH0jRJtZpDS
TbtJaEpdhn92cveLmb4HO4eIFX80+IjR8sYQLqxqL7qYMOlNYIzMU3C/VLOG4z2A5eAy2JXUc4rd
WXt2/pkVm1iKGOFrezzjNMxSZpDJFVP60RTEyUEf+hOt5/srARx1SNMoxd3iVtkR8ytYk3k48Qut
CMe2ceEaXqwVxBoUCz737IH5TjVuDrj+1YLnuLUx/avyGS7iBbmJ1oxLDro5LMynCdnxclAFmevK
NHwHdm2GlL1/+7wlsAFzGxDOqwaMabwMhhVAlQQzsy4zICMQc/33iqm3HUrEj96blrpWMS7bbWWf
81Tq5CSfTr/YoO0r1kpsD37+zEDrNii4Sa4bvzwszThQHK4bD6Ox369iA0DNQJLs4JW+gtqH+tyc
x0T5D9klBHE5uOCCxNFVzNrDw67SIlsgeUeP9Uc3u3Kku6DLSt9vyEYb7CfPNKSZjG8c3GRT23Jw
DZZlM2yj7eTe3noubwcbIKDLLuPCJZXTJV3iEDEFTzOVnLfi755ZgT71o4JXQ1aGVJaVnCWCAuvY
TQO+pWRSVLLURmXp8K+Idz3HV1vu0RPwKVo2FyO+kzSvKgteu7Gl4qAeTWcyC8RSCEq8ZUR/XqUh
pAy7N7/Wp/F9AL94mi+LIH0rnq5/Ro+5r2e2jhubG1CFAG14EEiyIrCQvcrkaeaENZvLb15jmqFr
3Edbfh6YI+Wo/Ja4TEcYc9RqioFIk8hmYYEsHoekR3r0sfGBkkJixLC1nTrejHBAjEyKfxd4vW5h
GPKXZfNVDUdp59pOn7sMB4m2n+JC10tTSjKJ7uJH1PMa8on6xJvtMuVI4GmBRsKkR48Kk2RgijiQ
SSAIwsIKPWpimlL979+jUlkGTeDn3Hdci/xpX8VIiAb5vuZowRcS4P5eWaCD22IZXwcksUIP74/y
q3gIn10589wEC9/LLcv3kPdc/GwDyf5oxqypQW0R1U05YesctwZI4krV6eaK2+qpVQEM3z+J2xa5
rgMgpRgJkpvQ/GEfQhKHqKKhMci6eLQuILVaPnbZFq/MijUNTlV39Yyh5/ma4eugmVFZ1eRmLZIU
FRKR2jvggVLn5NaTEDzM4SqGuTlnFMIRQCVscuhp/nyb8KqzBAz43SJbGr0t8o3o8xfYShEKzKAH
YRJ4PlXSBnap6CpiOBq++NCOyV2v442jcNv87rkN+ihaYGqT7Z8kjVEGFRcMUQ0bWp9EIDOsI9iD
wY43aADsdo4BnUv7HRW1pD4g9ODC406ScaVCTNd8MVtSikV/10dnkQFoFQ+Y6QmhEIFwI8wNPjaj
DKTIoyRVefpmWJVP++VmJ8P2HWEvBxANKiaeZp1DYlZ8U0V7k8VXmODk+DFWnPuUxvISZtrvVQZO
SSgN3FUZZz4Sm9XvfbWdtkMVg6HSJ0fydsL2fpIGn+UlYDqvV3eXb7B9aeu8uqWKu1yJjon+BlAB
O/EvIUNSPEA9WH6/xLqlqHy4l5aBIyKrhBIQ9Bvn6RALaTSmpV9vMm+BxLBLD2SU5Hevo0jVgJ3b
tUoue9Co3UADk1e/AEAh5nntnhCGdOfOYCAUyFUAICnvpdlX+SBArDDnPSPzEXfUKukkeEUZJUfc
tY8VIxHrG3UCqLog9LOyb1gbGgPSWFgb+cLn5GG/TyKa6Tu2V9PVctCdHIzxYAAgz1bNQEtEm6eK
o33DiYY8xzgZJ9xvxMXa2rHPezVWqLsIQ3nvbdITvyngboxqZ6xXfKvzchM6BLMMFLd1IEBLtVG+
QAYNXMcSPvLUyWWCZXEgh1rbG/03FHhnpNWmEmC0AKZZiiAxeUPm3FdDVevAuPoIAEqVVkzcUBGF
JGpvOomDVVkoONh+xmLqDoLCtfo/kl4oz2hBBXjnlAwO9mv+I5rC2eK1kQ2KchpROYv5uyr1DGsg
nXW2kbGNgn8wAZgFqdDSCZYa4dN1q4z6vO/+jEkX6u90lUk83UUNmQd593ELUuzckT7kI8g6Q65z
Yb/uPZdTw3o35bj4meWFlULfGaIy5n3wp4s3exUGmeA6RzMttp3nas/NRaA7SBXS0huiA7e9Ko3g
xIVDIZwwASRuDnLb0cC3Db362jsGi/Vo2DW+1Fh35JeDyz0S2oRVJArzQgDb4aCWCPLnwXtWP7NY
hqsSfKb0n+hLtzkF9zkoWxZBVeRjocgWKxsOouBqYkLt+HtIH3nptIAOf7fY9TjRDLsUjyAkuZv+
CbvjzwOBGilIyqqrzFWX6CiqNBSZ+Nzgy/IRnkIW4ZaL/Be0KlqwlWLq5oLM1YTpsD2TEi1egf7Q
VYgeyOjBJY/0zXMTtZ35vr7JyY3v7E47J+bWGjFKIXqa3LfMntuJbE16e64XI7ek1HSsavYVR0NY
HkWJz5hSKo1WQSOb+jB8nmxoFM3eeuFDBCs3j01SXVsr237ZHXhy6HHjyTzBTffulHByUqEkICrH
KBSvgw8RJ8tkuvhjF4VSshEbK01cKLPS9yhANwfKjXUuq+/KJA+iI8qiY2bl8+UdCDfdIg3BXNli
ZU7lHHgEfMhCeDQaFddPzp2xw5yx2oo4bNpc4SfM0HqyGrLV5DdRqQDcKKyxLfIG1AYLbP52EHkz
VcSbiHfPFDPcYmrwMjr5sru++nnNUCOldACt/z/eYI3Y7Z72cKqglUUUedbwfIu9nxVJEowMzTr7
Z9EKs5juwqpk3XC2E7blu8Z1Tmvbb1kmlGP9njOAJ68uqDyJdm+gB/nxnPYFdaW8rvC092uhKTqp
vBpXY0YJJMgtFlNmYt4TGLruQGt4NgfLNEbetkZ720VMHuN6bh8c7F7Iwhw7dTHRzY5gVyJsh/Ja
993ibg5PtHDYtyqX+UeCufQpZl23FqZZ7wYTY8To17wlY+lEGSi50Hh9RiwC7CvqIBVsIApmKiMv
llKU/CpMX300aD0wmIACHdU62aM0e8bzurQ/Mwj03xpIDEszHqgtMvFWjdNFsftK/WvAlQDQ0qOm
dd8ZZGNTzvsLkukj93gOGaV/c34miWSF8oy08xlqvKTjCtd87x80NDtH7leb+L3WY/lIALxXOeOZ
+dKAcBkw8u9O14WmqN/e20J4rBo55WCj526RVYDnV/Sp3pTeS+FxdZ5SfelNm2wChiRpvvjVHdHr
Pl7qtNulbKHtHjGRlmWPolLEzA3v6fEDGQRpi9vdBX/zGBr71dK1NLPIIAJ9rr4SloQDPCq2mup9
4FklAwx3gPbsM/fopBCaUzrirp3+qpox9QKgMOuLV/hxDovHZkrHA6YBvl2UTL1ezybm4sJ9aAnr
OmdJieHX9pq4zJQNvnV0OZEy2TODSF6UjbjNOhp9oxAMs5NAsLxsdb5A8lJ3TIuK3inZ8cHfojJT
mHg0fXexAGy0/NdOIbWgp+CymqDYwK1tHCMsUT1FhJYk+QHv2zCHqqqtAzLnpiwlmiMkwBSFA1jz
uKKi87PYZapYbzkqnjADY+JJViKE3w5JChjN15QizlfEk6DvYiCwxc12zd9fQ9jZ5JJNh4FmVkLb
ZPKWGINIx6CEVJWZGJFD77WYKG2+9cKhws+PQmg433ubD/KhNDc0Pye3prIEgGuQOPICqlmrkCTI
K2rIN8g39Eqk1vGwMgk0zG5msM8ZVB67UslUkTcrb+zpNSog/pbebl5ngk+WR0BBNrf4eM0TRqHI
ApmIrlxyy9yhK1QFo9Tk3MGiS6bwmG4hw14Sm02hHJdm8+kHdMpfala1w1hdBMh0JybYdN8noiQN
9KAFV4y8DfL69VqGaKfD9suNxoOn/DNw/yfyr/vBQzlx0gCco/LmY8U0mexdgwUvmwKXd/3KHnwq
2AlQ9Gd2VBGNwhzICJPwp9B8TTiQpc3HnBzjEJ6xtnMTFrXD5YH3tPz5reJH1W5VnGejqSivKwvc
6UJ3yMX0XOXAVd0zzR2aZWdAASgkyT+txr/B3o/BndPSjWJDKwfHQhR/nmScn3hyT2+Mjg0lV/hm
219zpPvff+SUMJ8AxYRezCv8xj3zP31pQFQ52t1TRJugM2qKYVXWEOoxQmPWaQrWknWJiOKkC8Jq
pDaVPPEaaKi+Ub4fKjtTE8kjtTQqng/lEDzwaeeCUMwcirS3uSW93Cw46VLG0Dfjdzcl/hsEYqOT
NPN78yAcGgmFueTA+Kiqtv8IOsqPJg1hIic3l3eFqqT7YjysjDJv/cZe7ZM1TCuIwMokN3ehxPyn
ShpsT4zNPU+A7famiMuY3Do2KmQsgprGFlmgD3iZw5mPLWWfBweMS76fgXhLMXJ48F666KQUuZ6Y
e5Dy6dTc6g8lq84zmEtpPq00XSslW2IPfVUy9TeLLE3HrnMheqw9pxBuafvznaVNkasyxFIaV6PF
ZnDl5AgH5H2h8FjsmL9qpjBY3vVAkOMsHVwv4YV1DtBBUv/aqIvA+TsvoABQbQLWHLI52e2XaMI7
Hcde1axT0BRl6GUF+M7rWRlSN5N1ZFrsT2vrB02i/OhaiLSBJSLSzi+/jSYVVG0uuxtvssiPT3rW
yJ7MM2H3e23d+ucBvKVn9ks+O9XBT0yOU00vhmsdtfbTeBan+G+tDch81RuGae2WYbaIxq7LrLCy
m/HRSm7Akch1yqesG7BWCMc0q0IAmbvbAeqaTq1tw3cJUxbja4E7oDC79gvcMHkfY0CpD1sr8x4u
4cSi3HTypJJHZykeDx3d7eUlRPrVNWjSYijycdBnvEP6NjIHq5DPI2Ew5/GIL423TOgV/yWTDmoV
dHriljopyjkLA3NfIRUFhwB78k1Pf/5UIGc2OXrTNvVdKE7vhbPfPj4w5VzwZhhwUwbTGxxlSisy
1fbW8FC4/vXgj8/WHJlwxrtozzoH3AqYu5HqqKXDkFtsNqRt7+HITHIqqryfRcM9FdvZ1JgVu4yX
7D+ZBeTRZQ3+tYn03NkjbEeFd6CWnJD2qtfXT6Mn/dAjUgPyPqPca6XdfwtH5SH2Xw7VC/IXbGyv
gRFXJvB2HqDGUwjavlMddnS5p1F1d9/X2QlDFx4doMoXqDn98xL6fVXUgFZ3n2tjteKX0/VqJbvq
R6X2+YFy2SkX18UyLnonEot6yljmDKRQHM+L61Vl1JGU6DfuOVsCfyjSTihHszlAKsqzHbueEu91
3oQKGBEJoVtro4j3FQSOPTAj2YZ5acPa/ApKD5FVGbKhYfeFecL6vE3zT598NCUY8kgs7tqm9K77
tk4Pp5Y3E77WGbFLM5nxF8ybetS/HltltHL7v9s+XhOvJqTF64gid6zogE56+KyoGzGLllfA0lNq
buP00U8Phi7GInkN3wOhTvQy3w5nW0ouE02hqLgondl0L99SsIODbWAZZdJlwlVsdKHYA3yW33Q+
B+pAfq9fW7CUi+FALyQJPZt50D1FRFGGLFgvO3CmMJml6QEiLWf5a9zjqDkK+hcsfl710qQ/Ze4i
rRdb3IZGiYcmRfNUdNKXvhBrsrHzz1Tk1KQZAmnbWUstCrRYlfIkcH8lMLVl4EuNDyDg6UkiL628
qu8y1FFRTBNf/3YWyNiAGr+wMLrAX1Sr6m+F2fyY3BTEsCxY93U/syr89F71mIMBiddwqUblSYhl
wbjjpFyP1DCn96Rfacaf1x7x8PolBeCV2YQ/znl37Nf+rd+J/++GkXiqqA4agH0hsv86I2eAown0
cp84soVsYjMogDXeRcxaqFc6tWPKzXzHL3FRVbin4Z6tBFZNtpcV0AxxSywmUZ/9fAvJ/d21gaoo
VX5I6cxbm2gdNp6YKJ9q1lUprVOnH2GdhODLg+EWp1RChjSsNC8AbRUVredwFnpbseU5hwOznk2i
XVYeo+ppsMb3c0CIQrVWGkjdH64ujz6EeP8cLzUGHaj6tv/gSmdyXAxCDz2dkAAYzAGybkvKNf4K
uWoTtgrZySQ5ml3Rv1n5l3CPyxpt9fKuyPAYTAbrNNe4QZWqnIDXoTl/wyyGuCz5oijoo/Wnpo0g
W/7gFLIuB2x/HRRVSh5Cm7O+9SfB44WjzqJKcTCok/Bk6jNRgqT6KvxQMWrRApJTuCDx96oJBRKh
PrRXQ0RG115djsFD+8JrM5jz2n5JKkznPmybl/tPeIGmneEyyzLoSF/VEXEx8J/f15z/yMhwvGN0
Oakjg57MaJm5NvOaCfJz/fzhG8yuzrOU7Fur+1CcKpASiomSKxYJSrjmLbW3hqPJFsscTub0hlpe
5Er9Za2S/w/LRTp4DVunTvjnucew6UtRL4//qqPWdd1irwXkivSpr7mR/EZNc/HlTWaDjEBoiPPJ
s8eqJau1wvokU8mP2OvW4XrlPxuEgq4UoMIUWPjI1eJaL4qrNDQMpw9RU3QdIZ7hXi6xDaenoFKo
35+QycOhfe/za9ZinrtDBkqqcZRzDTeGzVGt2w9xZ6MuYkPkL8BxE+5Ypw6UEU8iJYMHx9J6wiix
ObqybHVTF/y1T3UvTFYKtvdO1fPMCFXe8ZKSLQZh5LA1KewKvZ9uuAn0+nua3w5eiDkuhdNLkOB+
O12i4LWhjpcwZWcjb/Tj9x7mvRni81dQSTOUIrhgeZIYqXcd0aHTWuo7RP9kQijFeACPaq6G+5TD
g0xbjq/VjLWx01uETQR3qspSCMzjAgebcS3z+i8MvKdYuzsyOYmX38o9Gc/qihcWDUtyAz9HJyBx
xJEPPLKnTvsAM1kMbh2rFiXFMXrJmC2+rEvpiTQzXIac2lj3sTSJUbneh6Ud7gGuI4BMHK+cZ/2j
Xb41CNqHHaJduox3gCEpeAZt8RMkrwKxHWu80GRyYXD8ad1tNX/XwN4MbiVEawEoBiZGmkqV1XOG
aAfycwRBTDljdJGHfAa0sJP9GztPDm3R1dlfXKr47vxxl8Vk5MxUH98t8W3Z7fOAP9tSTzGRmOOr
dvkXz5AIsE0A7cQVel2mJgslY8qHUQnLkqLNfIV0XvOU155EYo7SqyKs8uEVUZVqvP2w/wljpLq2
3kr/sjX8TVdLe373ELlnz2qSQzKki+F+ECsa7m+af2n2EbDKQftVFUCizscfebxU3HtsG6cHm1CX
yGJTLaYfftPpHZrHA4Ph2Z/fZzdGlbVNw+OpDpI8af8YWO783HEfRtrGEcCovzsr9S81UTLMZMYr
/eYOAeoIrG7cQTNrbS5vSg1E/UAfJyN/G8fbW3GW02zgUAWTGS84d9ukGmxZzLhYJKk84t1FrI0D
ni5kNGztOKIbUfwhDTNQmhFfFyZYgfw1+Km89Dy9ISZmapNdZojbpiZsER5WsA8SY2V06lJyMhuV
182Ks4lrCaib+H6P9oAdvbRZUvb8WK8gXVR7IcseLdPrsI9LYwscNBxMcA3qkGe1C7dpCUhRbron
BsoL1EfmRydhHCFNSRk9VANZy8bJo9iYVFLwC4amGElqArHY+IJgeFNXjQiL09UlCO8QBTorP9sl
nkNzzVoG1uy+aUPDDvCkjM1EjTdYp9XiVw5p1VhCTqujh9UNn9xMhJlDqMffDwg9F8bVuB4vHFgS
T/1HbG+6AROsNuZPnyvx/cg9eKDQ3wec5yqPU6xGEU070vqkUi8UKcmtWgT2UNoqj4t8D+OYh/Jh
Sh96aVzoEPjROzfYwi6MdM8uMQwAamkx9o753DlJkRcPKUpiVyRIOTm/PDxbU3P6TCC0DjUU5QPe
Op192o47L+ttn21DtHCLGHLyVbodoWNwhoMExDgn049pOyrFejPMHFWyn160l0dCFvOFoIL6Flbm
rBsbqd6Uw0nQLXRSd9XLlJ/nw5QKeNAhU4bl4EdIIjWzx1G9qy3eZjaJV4EpmDxhTQ/PiPFN4Q+F
Syga4d52grp4vPaynJmJCOELNhFdEwX7W+G+bxRiw2JiCT2xS5v4AwOOr1gGVbLkZ2QWWDOmYThk
3NbWWeU8/8rhIJWG5JrlHk1VOK4mpLfDAl/ADgw+4aEH8ifc3ZWXduRnujC1SIAARKACHdbnG9IB
mZFZEIH7C4FPpcS2cWumG5v75iUarMCuT/BZD+UVi4ptHFR5iqVHbwM4woNElMRwB49U+IAdPP3X
NiEEgv+GAisYlRc5w9zF7CEYtlZU4j5AALGG8RflapUzD+fuKzxXfIYfPSYFFWkWPplDdhB/rrxY
ZHh4ll+AnEh0MvV/o8xmJ90XJ7FwI7Qpk7zQf9CJKlfJzWA3l8KgV9iqqVfT7GOO+zWNpjCDlpZj
+EetDBi05vDbbSnHGVM3rKzfkD1ezf01IdXbNmBNxC5siPQYqSZGeo8VxTWlMSqNUpGLftqGG8OH
YyL/r8LEskWqTWnnqdx/1aEBQiK2uU207vYUvHXEdnp+Tmb2bQiOO0AJ4JQg3MJofbSmomLfJPhU
yc6O/7CcqoUVQGlhitZ2Yj6K2D/tlfDjRwEKHlM/85qVdpxVNP5YvYluLFBRVCf0jVC4mOmU2685
se/Gie0+QH4526sqk2/AR6N4xRn5SKNeQTqrouVNVu/6Ixay6XA6TU5FT362NQfMGt5jokqkHjmo
LBKTyMTx8MZbKD5/sFAntAjAbgEgDMaYBwqsP+qO3EmcHb3Mso1XYqOoRyH3a15jdqq1D7Yy4TM2
jnR8tmuIKEK5+PzQmgvkCJg6T6GeHiF+Hq9G5pQGFB5w10zH9i7uGe5NawX8R9ixOAFvKOHf9isT
JCm6h7TtuXVCnRpfWD7myTPt6+yF9wUx0cuIOrNtsOhWuO51Km3lrI/56CFoQ3Rt0il8XZ8BWWVF
eaZorQAKedqmd96aPDhjnpTutaBz9U18jUNjrUW9Ypi0Cwpwa6sY4YScAsPOnvc4KRCWAvsDu4eR
k1Ou+qOVqrAFHMLM94bul7nk/gPG3U14A2k8mDMJVfHmI1ZB+05w8GT1ryd8pgbtQV9VF8MTUH9z
DVUw6eK/T1unu8MwUzdvTFwRaStXRdTuMKHmNfHUEO8WXq3CRRkkqSUQqjzbY7FRAqvz5VomYeJ6
rPe0Ar+qalxV8V2oHwARQr9sUOtb82f8pS+9KzVGSyqGMSGpaQzC+5XXx5ye8x/XV1MDXqQfHIPS
SYdcUzzI3Q/3tF0fgUhPq4AP7ybQVoksIEfdG2Lt/VBItFSUgEhZlhHKs0pwiTKsPHh1Q9+wFjE5
rKb1q2P+ZKphxgA0I/17r3V8kA/TFn8ilC7LWGtDnu99VNaK/sup00oBhzfFFc6J8cO4SCEgwMqI
0e7l+GvNESSL2qdgUawcOTtchY6nJ3iWhxWZP4zI8zZmEc07C8G1CRNpBbEAKIyqZNSo+7/9qd7g
uRy72UfwL0ksT+e4vVmx5PTRDlUuhYrijIrD3ia1Ma5ywQbbm+bgbhQlzVPluAZL4PFpuXczUBQ6
uVOx9bJPqTI7j3ByYpdc4iscWxhfAqR4np12JmqyExQVfsUA8EjoRTZRJ9B2V6n1csUZp3QyZceX
5GA69mxGvEBKLm6lvhkdYmIL+mZdWARWAMxJSxeLkQ57StTz3rFlfR1m0gT2wUYdeaovaL0yiMIl
5AYWsLAAS6j/QRJl+KiujnseOUaJDawLM9Opw46OGLj2iDRymQ66DWR29HqCht/FfhUBX4xOyqTU
NkYaL37XdgFmIJjKB30ZnEKX/0yHCS5Nyl1cCY10gA6Ii4rUnVYk6uqJk7Zb4uHbYZUBTggC0TtR
Z3jmERHyXIBxXL1Cd5YdzT2eIoXfHJJLG4DtpUPWMC2qWNmrZLDd+Z/7YhDXQ+UsR18UAKNuRSRj
nVnHryXL0cYqpIkfWWP1m03iYdiEjzgFSIcOOeA9WraHvCo7J0NxPSq/kLkhhVWvBLuA8+VQGJuV
acQDisIlsNDTFosK9sTbmZ3eAYOcvIFmodOlkBbf6BsK1hU6tuyrYKqxhi7vGJt4yZjJ3n/kRnpz
0il7CJBUvbSQJ2oSkjRLqZ4ixG7kbRddJBLTmAdtfpEPydSfcIDcI3jS7caXu7bC8CWmQZPBrn6y
ENepsJejWPKiZngGmWpWvxR62v/I1atcbJvbvSKXT0jm4meuCAj6xxZ2HBHa4LzDbjZv9/ub989+
UCuxErEcauhIDAbOrddpPdDnhOGQBpNyCX63Dr1wGtU0Ab3dtyoWy39l1j/G++/tIYCMCSVRVVyF
gWoKdl/0H/qqlZzaVmGMLzhQZ9KwvmbZrtLy3oLB7US7QNyRg8IuXK2OBNwUyacVo3w2+txhvoYW
2NxgL7OjR9u0IwCgfmN6iyE5v5kfvkfCGrkECxVN/QyuJYOrzZ7LQzB2h7bm+FsQ7iscCUii0Zhs
Pew/gML0lg4jWvPnUPzVv56frZplDQzeO+Yx1Nvnq1/G60SqrAuBHcBPVPAjziaRbIgib4++0XtU
z8/WSwQa2CpT9WugR+y89iYlIAdYIlRSkfgssuhaUuvgYcKKDbkPmZwViwnCsXbuHgKFDr79+WNH
wnut9QP8v4NudavlLqnQqgZ24Ujoh4SkNHbG8KtsNCf1uquokNy6IgbOKQ1WbUfhfrclJJi6z6tJ
EeJdpxq7BZV7CDiHnolWqBzpsyF9YiQctqHT6ids6gTIO4wW4ryE6XevlqpNwLxLL6Bjowa05+QD
kiVVkjydGJO3JlbXWL93njtOKSKzAIgO043Vh2wI4avgOKqU2Z0eP16JmsgQ0PZ4d35/tL5uZoqa
gOU2/dPdFGSvd0892cYWczW4CejdnXtVlZ67YpIC1QhE3Y/xaZnOYJB/Gik4mmavLcpCRz2yJh+N
/kFe6rTcPuqWfRqqG4WVLG6m0MrRIUDEIn3eXQ1FZzSTWUCFcb/7fViMDeIZP1JjJNAvmNavOjwd
eNvKU8j9uqkIbS0QqUFC+peBPB86pNCHh8FTJnvTGVSAIgdyRgaWyuGKo42zKZ4MWvZCBY3U9dun
tOV24v2O6CsZyBXbFG2gvaEhzGd736zwzEYciSixMt3rBPNGx8e0txEHZEFiYDov57IjL9wsjuGT
LQVa1PJ5/jLcNzZjbiGn+2FISau3GntRJv2thGviqNJgJ5PUmjwpEhDVNwt/jxPwnoUdRjB3sqJA
wWxVD8M3hvlzydjn6yfsemAdEPKJmfhVp7zOfjFzqMDO3OrEaWtXLstf/ED+CaQP1CTp8Ks0i+Bm
SShwmJ3N9ePJDwzycNMkNEhoji1BDsjAqivqIejD4QDoLAH2oYSojzXOn7TKg8BeEfEoJEBoRhVd
BTkHXTpY/hQNpTtzDMc87nYlpR5J7rFXJWZ3z0yd24TU/TqFjtS5WVwqj3t0zQ+cJbg4xzp8StXx
mTLQsMK0hJY6HYcz54TejllltflWEEvRoYuaOfdSPtXRjaR2Hz9SsKkpQA9AccjoHU9yHpnkl9Rh
SWf+1BhoNqOQesrQZHDC07BVY2p1HMqZL0QY54F5FceRBub+AvYDRp1ereAK/kVoIhtRFxl5Dr17
0omNpWjJu+iYJXNevvj8xDU7lPoVZjYveIyLVcdNQnusRAT3UgdwTlr4wShuaE0Ic8dbMentfF72
L6Xk/sXvJCvi+A4wJcB2aH1OTfoaXnYjjgpggmcF17I1rkAg4GMS8TcckfQSjELr2GEnoAMRESQc
sLiv8/LoXw7C6lyHfPL7Fmr7N+CCeX8qW5w91RyC9ujvKH0KllRXVYlydeGXgFR/y4pd5BB4lGns
9RBtSLGiqSRifftnhxttjQPj2Nihf7o8VZZFJitxnxEJj5gA06HZqfetK6KfjNp95gcwm/Z4BWeu
AW398XF1xtmeQ6LVsGeTG7CVZTOBWWkG9oSFbI1aDRL7Ii17/HuJUWbKTUdefML2/O18Vr8TXJaf
JQpsODgIlqPmpy/A/k92/H85qeUnaPrtrluT9/d3nIzf7W6Ef8Q2ZuyISc7wDJxshEqvvgdqu0kE
MIueISRjlcOe8hW1eiZHeT097KB9zY+0DDJ4x6pEAqm7b3LTQUSCwtEXXu/iwIxv3nUNgIUIzrV9
HSHCqndm1YG8yrShQ2JcckMhcd0drfoG/tEDEeoki+XrVogQ6kXohnCjUsmIESYzWCGnJqEC7cuA
YRa0dFdwus9miB0XI+sA68qzsA2A5criHJcDbgk8f4olGsf7zCXWdCN1+NbnQnZBmRIIRP+guNW/
o+tugNEDat7sCJAqnWnfaaJTgFrS5tBl77mKB/mjEH83PxXGF85gfFn3ZMvEcGBx91PNlw8EqFtC
x/DG3DCvgEQM6boX/+PiVGS4qg/VqrOO1jc3qNjmeT8YfjlPmgAbjq18PQb/tdhx8emX00NvLc96
tOGb70XjP6PVLTX2NNiWs6kM9S/CWbVvXHJszQq20Dimh3EUHdrAHUuUhBgLhzdXVWHwd3P7Gk+3
rPXTpicG2Mi82cFGz+fXQLqMomenrKV1PENXwjsdETv6/XrG0M/imbx6pbcA5H60YXmxqCNmKfZH
VHijTsF+9+a2U3jgpoqU5xj5Gxx0BIJ/uHrWkpTPO5Jcg4VPQwbMCQ8qco/8QpjueEednyOkF35v
EMNzZ5IFZ72cprIbKcIcTz4hSbTpi7CjJ5ThBZGHQppJA4BSGXBb1cQBGa8SzhHPI9jikFdTO+8U
5nD5ruNYxOSqyha5n5dAutjj5PjVB2Ihm55HfVZlk7xkhFnDTqm+IjiMFbrsrjIM9Z+DHUGV66XH
56hkSy6UXTJw1/UPvP1NnmfjDPbHbZ0C/zV3HItXH0JVEPM4E+XtgRbvNcbP90e93ISEP5hZLof9
EIvevL45Fm0aCwqvomHdXaMyYMYSMMs3tQcLjwXUqlzqZNyq1d4WE3WuTr2SEQTfSIp0tiHADs1S
Fzpn8Ykmf7C4v/8o0ATZk34OuMXaITMqO9quMZS/B9LmSOjQkvBVN/KlZondUHY0Sfc/BRY4CAzl
qyZAMkg8i6E8vph8iyQ8Ox1w8xDvIgxBzHoRV5fnCDjiCLP+LCRFXFqSyqJBsr3bgOp7x9R4Qjgw
nbpXExNxq2cOIJsrHMRq6MCWzxy3kMvS1YzxMhniv4yJC/wmOT2UfPCuYLqgiFCU0nAy/uQAmKYa
PajUDkMMm42vYrXpJDnyWlgz2NGDbcndsMRr85111jl/EdNm+kxFeb0elr9Uy6fjsk0CwsTtiMCF
KV5VTUElkE88gH9aPM/waIMUrcaSDKmSdF1FL6n/9EfnER+FTIq6vqvLKpo8jfZTNK8JcjFweYOb
kkmUdrgejymlAAXiRN1s4I4zchtfjBkafjvApUQY+r80BKLU5AtzDcj3DdL4hcKpks160390npZ4
llf2wc3ormLirprRtIg5Rgqkl9IH0JBNqHJH1qWcZEB81Nz0Dx6V85/1MkELqp8y3q/IHAUM81/w
hq10EUavBCm9UhrKRaSno6O68WRRQNlJG8mAupzce+4N8cu8W6ueIC+Rqg4z+QZoFzc9QN0GBjNI
wfur73SNF++1s76goNB8SeqSJNm8SxUTNq/C4y0xFOgst8+lUVtePUjUwNn/B3VAivoqzgIT66Y6
NYMgUFL9dtobuX31RLWFzFkYuKCpl5JxpC8nR6ITEV4aIJP9XSkzmcPCfSdfG46LnCqwwUr3fetE
u85zbffoxwb/dT9DmnqcHfNqeLhQHUvZ4bqXtQyEzusSP/4c/jPXFSAmKwouV2XDRvdV/2FE8oqD
JwihZZQCQySq4YT+b4evkwi4LzZeyLx18zzTGay9BZSdzdp1qrvT418Dfgiz+S66xta6Vs1VHrJX
2llMqL1wwZNCI6SRtVPPuzJw0/duKU5Q1wXQtNvrBJaL59tosCPlZWWlk+tD36qBUhYHQ7U87hgA
WVjumAYpO2OC4cWnMiBjMXbqMoECJolMB3nU5TsNTWh+4/rAuMPuw+5B20qSEfPJRxqxCtMd5Pvr
x6X6bgB1NBuiOXv3Jj3JivEymU5baQBaOC+ADDyCNNYG4ICNTSdkT1EbSC6cTagkr4XE+jszNJ8N
4LccTWSDKbEf5cE3Dzi1uTLFMtEFhe0YL54wAQKPJlDoQZqWacq9wBOVdQDIBrGzrAXs8JbzQ3VD
1JwBOOBmaYpY1YlRfm3jp313K0l8caZUpN/XpQunxzZ4zF9BUTQwRyTZFEwehFNMP8fnTQ/0OjC9
h5eblTYirG0y330uHbcHhdZvPX4UU6bHugdvA6KNGUDF9FD3s9l+n8s80Rzdjxz9JvYkb5Pzli9p
jsu87GYj+tdQz2dd5cJ4hZfBcirHp5hnHup/4PhnBQrmZp5qTSGGmN86i5qtDtps59apqQn41Uh+
+UCDaipOQyTDVBpmXEn4lksbOKjGM0LoGK6LTEDYtd/6085urF6/A8xAHaiU4APEp5BCLEN4nDjP
TXA/O/demBu6oYXHu9+YK5Nss8Evy31GBoLYow7ILojdvkGy+X6+rJAMRUcgoI8IaHKR9qG75zs=
`protect end_protected
