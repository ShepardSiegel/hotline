`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DppNp8NRNvqV4iOWT0JvxEwgZo+qeqqOaoOwbgCkp9hNMYFrKkHmfyu8hFaXo5/plHHkgbxxv6T4
z845yds46g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B2GlU1n0NSukbD0lNtdjUcHcy5A/JyxJ6w9HVAeH0r456H8JNIbOn62TPo60P+apV6GeqqXzurt4
JbP6/sAI1bBf4DhXo+WLHetD9q7mnwcG5aiNLYfbkEWnjhSW6sQUIhuDGn39jos19SovbkBJVhUF
Cs5omhdChepA61Sxx2Q=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MZmVheqHSz2CczHKxTzJ+sQLpV7Ek5nB3041WowOFDChIPIkksRWR8925JVoK/yc1Sbx2mIAXhOc
DzxuvE6532pSVv0Vzqa8X+cwfidrZJjQBYeTe0R/Q309fUxzc6vw2EsuXbViqvo1KbvglUX6Xr6G
EjFbn7VF1W0bmEy/9h6PAigNy4rDmOIUEC1ucJAftjcG4glWIoR1X6II0wvo2Sve7sAAMQfonJtk
ZBBQdtVIcQ3gDg5pztnxxL3HhtTeTBkePjmY92UNp/36ZNpmGvi5HP+374TIV2VgEIkq533ao24D
O2KynBuzJWpaGBQVkABcIb2wgec19aAGUcmbBw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Nr9qBSuNqLR585uQc6G6PaiGDftRxB1yvIxWFA7SgH5SETVCeB52SBOf359urRoDRYaDTGATSO/S
N4nWQ9FsuAojOG3qEo6FvtMW76hK2lnZi6Dv2pwanJsik9/VhcdQImjRa2+huERaLiArTWeO00mh
tudt1HEdRmMTY5B7ECQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EkSUwWmRRf95kaGQaWPEJz1YLv8p4zAXxI1h3hVcbl5GRDfyo3D1lOVyP4mYZnoXxbWMnBGae1Gu
UwJfLWXv1K8dL3bkArIwiqdifSnyRBLe9LdtTG+u4qNipjAZCqQJHDZVwjox3uxLvCTABZMqk8ku
nX8pLd5ohr3agCaF0uyo3oDwtPJ88MZFy63RznX5FfdsEl9Q0MgON6dmcy1+S6qsMk21TTG6+Os8
eLv4+nF2wz5/QqNuB4QulQv4t+E1iwukD5OwtfEUdcS1T5GYafBmDw62oMvTP1Q4ksYvbxMoHzeF
9HIb/1j+0/MM9XuY9js0txeNubEtTGe/FLATwg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12560)
`protect data_block
J/Q+yUsewiKez/NlAgf97UQROvZnMCvEZMmw3iG75mGoFv3qmAlZbjwIdkHyRSDxPapzRgk9WZHb
L1vP//dLd9HKypFOWHm/qfdamrEyLDvqt/3a10/sQsPVoqYBt91clhFCru8eYU3uPmEHzlTat4HA
efgGArigXT3butst47MCTEYQtM5feXRrcVYbsqIqFZKoVFpsJqVIpUlP8Si+cYfshkt1QpfLPtXX
6G/tl4BGwepQCVVDLckTh/qAlR52IPsprv5HW0mtg7pT2vdYxfrDQWZeJOAMzUmG2/SjJgFSMr1g
XWcB3JGenwTelHi4y+LzdQqgjLeKNH4nH0g4CtwV4sMFjUgW3kb0aFdd231l2wtEZLTrRZfS3GUW
9vjDzKl77PrwZBA4PeFH2clj8FDuVn7y6POSnDRlAuH9LX0KUuK32D1ArU4KpE2H+lsCq8RFNMA4
sN41WPk+q3j1Mk9wgytj6M0OOR6uvhLxYWg2mZKRJE2r5hPBD1UdKyVZQnx65kcjA7EMME/3fgaQ
cd9AF7CNmibg/wWWS62oLOdh1RsNWLSkRluPhX5q1SInPHIciMW33GPz1c6sr6rGZ5amycNAvJYx
Q4Gm9eUjnX1SBUiQ4zsMtaE0/9DoSYmi2X4NPZdMHp3CwfF9xuPtoWpMLte1Bjf4ST5kWstcNrWW
CK9WEw3FEtXxyBG2GllJS9Ue0ijOfHs6mKY/p+78Vf/v/D3vOMUggKYrj5RoAWZ9/HTglXcKFpaJ
o228rGqenJtQ7IhHNvANM3qZfBn2tW1tOZv3XYta/v2IPS8xNxCYxeS7qRnj51gy92J0mSGVqrWX
M9MEXAftet+4GBXg/ouWfy89jebHg/PJG0WvvaqOpX7YlPNA8NQBXbSGLLH8zaR9Al7jhJWPpM4d
7csWCZhQWIV73i0Wc8UbBI0NwfxWY5zI38Bi/kILpMj6E8gT48dyAF/GWPMoZTYXMV9PcWr6gF+8
Xq06+LM+wly4qUZg734kTCqKvWJrzrr6bjsMZONCnQu+8Mz/gYQxCAce03VpaLlcHTRbSOaYFpHc
ZTsZse2HoFLabN5h6NuXjXNSWhcBhAbesmceUdaCK/UKaC6pKTrEsoR5PubU744+eppRBHV+z+3/
w+gpz5IvoWOeg5JrPZWxfBDxolOt55jvvPu3fZET4EOYK7FLRDytMWyeDud2hYuWjcv5wJ2+Xu2J
dWUJzjpa7Kg2pnzBv7VZwkUXUgD7U14b7qOaL2AYCsPIbMa2MaGTOwKWOYOK3QFf/rXdURkZwxRT
/7qPaa+CKQgCJS86fthnYrklJSVa+6uhEcX2UcPBiGEuixJuVZM5fHqjD0/2BymLJt5L8TNgDHIP
L0r4dRkP1cOqi0bO41ME+ypFbvYXC6Ajuh9buyhdv19iST2znIzPEHomU/hf2hSO6veaZWfqYl2h
hKLnt36S3ilNWzdNlDLSQWZO+LMsWeNNnPDMwhV2I/w/b/xkcPjM/IuWTO4bsR8mRQjrxI8hmB6+
KyTIOWPP0eUyU/wQeRHJmDl/7YIScpOuTAV3feQ6pi1I3ElYEtMlQj4DLx/xV6hRB6wGnms0LduZ
8BsZO/gmDDQLUo+0Om3v01hhS9NOxdP5X5MY1wZjPMmKsx1I6KGJXRxHNFIUVfuS9HTOUV4rrRXc
wt7WOdAi15dvES8JzhbcCL7v4WjfjqP/Al05oHI6KaDBYov+jl+hGnxY3vZafGiJJtHwmZNw741h
B7LouepgAadxWA2yzB+M6I86z44acqgeuDKO+XwfBo/jqXsHG2urcHsMDMdgl1e8uRd6YQ+l+/dY
srg8ev7pSmcl3lr7dYZYEzBBtXSSxjT5HHkqmcLX/zTWYJw/16YOOg4VDXpEr4YmssM4iTcqHvp9
BgHZWUlTkvaPoACN6wt4P+k4sMp2FIfaDSB3tR/X9KTOljUBIYchSThlNNnRs0y22jSKu8ua1Rbo
h7gxYOE+wXJRHmKQ6d3CTTwh2javsSDEJUK4wp/j0uDvVWv8RQPR+Tg9FH2iX698MLWqhyrsxYiu
Hk5JG/px7elVA1RnYNt8lqfnqnS2YupwhMlZyD464zYev7Fj/p5Wzxp2Sk/86Zi5amudBqaNaNjb
8/cPgzpjl1qXEO8pmJStD0e9ddqAgszmTMXWtKiIYKXTWZFukppmnQaJZ4Uv9BWGy1QmDtJ9v/ap
fIZaYdUQXo+wFBCXl2toXmI9kR1Zmu8TeKZ97q4hrNkUaTJFmwcuBR9xb1vhNSXosnj5Dx+RMorn
pxkQ/LSTcmDcPtVCgnDtiDwaW0bMpxrLFWXsRLSET/uEBPNX9YU4c6xasnbKqRWrIem5Ub08Op2T
LBmVB8gOOa9jt/lejkYOQlz+wLaoNT0MJbbPk4veraNcthTtl0brHOlbJEvnNJiLHMURdADMTd/I
AHvMTHzTcMRchR5CCh80Wi1F2QONKhcyCNP6UYnn63k0RN+1hGzpZDu5z2ZnhANqQBU35DM7Ojpt
L3Ag1XM9kUEINFHsqpOUUsIxMoRxySo/EH+NX6LDkliL/FBt5+eoSJR2fnT333Too2KRSmKsHsZX
J07lBkK/uKvFxMBntqZIMTYdLJMPocQYjrTas6BRZHXcAo4fBpQw3hMyjwsy/pMIc+Kfr4v2BP+w
he/wL+uCQSlobKDzLvSd0FF2ZOK8roLa2gk4iHafczTZOwMrtadLp/75iYEof3Gagxnirf/Ugm8M
VpKAyQvRrq0XzigjYpLCWa0kdtIY/tpnEe4JtzbMuBdGXGoSoRWDNIzOcboH7+KFhDILjnYq5Z0o
S8M1tDD28WNNWYTwYKRduU+R04koBJwKFljziNj0e6uJuY2IXf4qC7AEDmnFg3SnaUzGJFvNEqLZ
YhM5fob9j868eIjMv/YOHmD1802nhf2l7LnnhPWWbIeymiOfaTXOfUK0Ro/tWY3+/efaHwvQRfwQ
4vcAE4uwwNuRz3tF2ffsISwf6J0pKr7svMgD02E6WIbgF4cqrzlql+n2V9G2nBJ19PjhEtb1Hhjk
5orOdSipCrrLUlHDkZA9yfXBSY+ae1/hYCi54mIuo/cu6bKPvjKTOaG4nG9B864GiEKEIQ7ag20o
DLF3UYrG1ZQj2/owrGHZhKkC/WbCeK+dPNEfMx1xBP8MfwpAsiBdhp3C4qM18qtFbDWYuDy4Dcqz
yQUSbz7NpBPh9EDNE2zcPv+hCWwWmJX8jftDRLuGxG/AMEw+FIuBbMNnoIrvPTyM368BFstqOfh5
H59qfbNMgpyFmlpvsjaJ4Y2/rlBZDhqc/5w0grKxOML7LNHPARSsQ9ek3JEbedqT/r+lLsi5SJ5t
fwJFRk1dfv1YPPBslVBLTTouaOhmENY310SEp2BTvm9oURJgQBcWTXOHIwaLi4UGofMCZsR0hN5+
p7sl6taaktEr7DCVFEVsr2QogE62wQMb8veFHrBzDj8esNqLtv/u+5smgUzy9+BJ3H/LGKCPnJAK
94d9LuakGWlJIpbbmjsMfFRqTRlSSmbKZ0zttg0p4ksBrmcvmib1mUZUKIxN58/GUZ6uQQi9HOU2
G5JhcHPur3TgN3MPERY9GM6QjisxMfTEHPkdUDS+KWlKVulmC6qGmSDnqJRWx/d1E+mp9eII3ErU
MaoeKKbQVYQe1PiSxyKx4BVDrTcuSd3D3ScjDT2h6fsB7++BJ+EGSanQU+VwPhI4gEWNIEutbJ0N
AXoWslaN4VpycRkyuwDX0RjGeXysOKLAurvDlZS+JSrYAzh0fBJMYBPzkguJ8D3QiSZM8Z38Cv3X
uNd1hJpCZ1cp3Vg/m6R3/NcHWH/Zj2Nq3Oy1zoc0LGq9S5/2eHxYXxyDsl+Fr1eMlzX3U/Z1nbq5
A7rfCG7aOvcjRtrlHYqdvHxmZSsYo0s/UBlfGYUnk12Cwk1ArCQ8PFDiu06bs1k2bQRjARyDYC4P
cxfjbU3zDNgZm9ZarXKNSOlXeZdoSV52RhxAwkgh8dpkFrVUwqNJY10Wdw88bAZIvmpd8jrCwYOT
oMfmlnjWQ9RXFmZkws4ouV8p5wiRChAnRGRQtbUIG/QyqUmovKRsUBQKXgjSxdbw7kAHvHV9rqYV
BM/FjMlKhR5qocMen0X8Z1PrsCL0DNU7L4NgPuv8j0rjMqzQguiS8csscPVWHnOvlmXp+ywK6OeH
EeFo6OTdVdoQxs5tZaz0LSGQMDTObo5I3OJk2U/2kzSJ+XliJ07fOXsueldn2HYZe/W06CenuxWB
zFfUEk1oI+9Ec6/vPSSBJfZwKOPsEccuR9uM9MvGkV6Q/0zUolKQVIg02BvqoVAPh+Zdvokr6+sp
St+jXmUF2BEfLrRAfVf77dTQDy4ptNn5rRAlXA5ER+qLPjTeo/D7LZaCzB1h0DI/egijP4ocS0Z8
o8+0nGJaX+MDRjV5g2RNQwFWXc/JgZmC8rMkhAPoplsX+WbVLXzPJmx6PPxoz7JSFINwjtjzknZc
AQBREdlFn0WP4fNTBJwmmA6tKUYpSA3nX3w66fEIsqaVwHa4+BsCDypKplKclVA6tPyuDtQGcid6
3X45iECFynZ+nDlFpXSUTyxquadgesEdOqeClC8fR/c2wLxvtsP+oUlCz8TnDcUd88MevkEhAGme
kvvnsbU7PGPCSZML9H/gbLdfi9BttlAngpPpjWGnQkMBYgLbbjvWtltyfXl3oNK8m9xD7CwqMHwf
vKBAlYyOrERuU9V2XyKyWACZI6YG6nID5SMjSPEMvmAUrjocXC3Otf70RoU51yXI/SenIufHlYe9
/8o3E/LhUCtZxZO2H6zoHUnso5p5PfyEaXbIW9Ad5zHzNLhH7eynPjvftNgaLOcdpK3X7WlapPpN
VOHQfNkaXNFXdJeK1H7PzrTi35eYhH1u7EommsEm64/nia6W2X3azOclYMYDe03hg1lxBjSFnLc/
SfLGo+HseBlXenVxrVO0djBwzWQF6T22165xvrTeRgABUOXYR6PRSErckzno1yDXpjw5SzZhJkMn
WH1A20/fORwfVb83bFq5TJKjSxWTGEio1uTLuDlgEEXkGfBKOXSwIdUpKDlNTAvjP5udlaZIbzLO
JFVbVnQCn8Jure8aT2VxtON9QPcf1CUzU1Xk2VQxwGiWsbkH5am7Pggxh9S2fEqBIYAFI+0Era/x
+P8f38cLZ9CoVR/Zc1GHrbOOEbpKy98+jdbeMcQ8trzrdLbiP1MnuKuV1rTKYXdr8kMAVF5PtVD2
fipr00P6z3jzQvNu3lMijDr94fBO1ExlcR6Pm+Qp6zUAEqyeTjivhSMyF6Rra/sOYWO6iD/fLk97
xdkGkdzYGdnhYL6+HiGCqLkSNkCKakY1+OZdw2c8uU76Uw7oCx52jPeIahwBAEMV+5gB2HF1QF+b
MrJHEUK3kW5k5ipP6H0RAieKkvPreL01OVWC2U5p3eXmbwYpm2xcWKLL5gLliTb+1/Jzj5F1utU1
jRKO02kA2dYC94NdKUbNdJ3oJSX3MKI1h/EsBrWFt5cIwmKJFL/stG9OVw9x4W16i8aSieZCX+uS
VNN1AX9J8yjwq+mPyS+kOFdc+0EfiuhRUEYVhB4y5+6RPIN5gjr0U1am6xUmGLdViGwH4KaEc14N
RmrfkCiRrJbYqqIoABRj+5vJoBJVeeaRL7rCwdF53zi9tN6ka8OkLcc+5yZwBNDp4MoZZvrIsTOM
/aomAXnj5cC1/F4tJdJlu50y5g6KFoB1dcQJjjlKTmvGRWjOTbZtb9nxyy7LLHWzjT7Ro8N4hcJy
rLEZt/hwN5XRltHYTJBfLEHeG2F4j2oOQBQtuiT8Hbj9678r13oiXlMhjpPSK2QmXaRgHUerPjaR
dfnGOtAtY5zkTPd0DDOnpnMuFoT4cHYF8K9W0GYKAYpL/r9I2d1s4G331hrFF//nUxh/YGkcvZes
wwwZQcQQKGQJrX24neVT2MeBfiJrhF1m0tWbiCfPHw3NhdBnJML7jd+t8YHBBQVj1Xu/GmvyewOs
2jpQjNgXbQiWXWLC8Wxs17lMOvRMIiRuA1EErYFymBO8dQhhOJuXsMCdf/pC1wPlmnGZI/SjfKP6
d5UJCNTvy3UGAEtLcpBf46x2jq1OowQhFPXi4dw1Cneie1bTNREJR2vD5c6IoBjOukIq9phIIPR+
I5Bgnf9r9tvNv6Ow0JLIxLXvOza1DAfWIbHeLWIaLH9P53waA74oxcA76lQyelVe15jXu3IwEKRu
/Nnk1S+9fQVXaWXy1ltjPCtFgaZz6jARn516GM5G3w2jtkprWL6Rp5cNEU57kV7gtmZrVp+X2Xy1
dDktQZasLf1/yz5urgC0feqCe/uOWWWjraXq/5YrCFFaxIZjejgvVNOKVCXzhygPkKt8Mz8bfhk4
JiS3lsdM3oitpTAhgKFqs4vkQLH/2SPZBMU6I+UAdlH651tjOFRjp4M8pGa4EnynVuQyW8JR6+R7
FsQrDUJfJskU3wl1HJDaqof1z4dZksmH8kkgE4kuKpUuP2L/4RyukN/t1sGeNH91dL9d94Ddbf6c
MpNHjbMUMqWpoT8zQobKmEOTnfZWjxHZGH/HyoKLP0DHH1YBjO1wX++kDxbywrmA9wgQrRDvxIzq
/SFH3MXlF+MihaNwl+15uqIuzm4i/9kn1MC2taQKbgFkHSU8+UnEig/G9kHTEzxihgYL7nKGg8mC
S8qEBM+M5IgkHnpcbgPOU5Ud7PEzyOMtYTAux/kKFqG4P0gGzf8O1hTvNT/8zrYwF6mj9rvwY/4p
W0Rra2rC5hAMI/Zm6T++q5+HD+8rdD6tXqUArniIBlOWshdWA3y6lBVqb+gZQaZUd5vOAVadvldS
Ro7WeFPL6/rdCuwaScA+yaM4lwA60c0bcq0cJpeZdJpAvEehcJDrYh3DBsSwBUxfmq3qF87HhOHW
GhG0Uh1xTaAG/KOYqMyjRM0ZPUXeN8ty4q9kN0b59cXSwIT6kZP+nVVPFsUc3+HDtMJWEPKJsfmW
WUKZzz1ujOu+rOGJlo+YFMAiC3SV3pBsbpEvFKDJgWjc7MDtN94saDqLg8/M22UGJL11si+jTTPF
eybHfOXMaXbmZVyPnLbOIYoxmREsDfK55yke1yrHQOMIndYpp0qQlnZWE2aIqRB+fv7AwzwtZiim
1V/+s8VT77ojAkh9YKCWnhPKfbuJU39PoLCAFy2Xp8qvrCZHGIY7teB3csTGescWNTkQPAmSTKpZ
hVIdL4gRMIQyr5n/4RcZL+yi1ZTei1wUuDuwBoDEMxZ7V2zxYcVboeUEM7btuMjPoxGi9w+PI1Wc
rDb+zxJZK1zWZXYziTzs29Fb4LIZBWafhyFEWlrgpkzCXXLfrkz2ZEBz4HyuQBcZuN1ULC7+IvcE
pXEm9PM00UeNs0xdbzvWF7Nr4Hhry3Gy5WAm7laBfsDaNgbh60DLANH7xqOlN9DPLp7zLgFCZ0tN
u08UhV/FoKo3I/xz9Vm1EjOV7HEJqGD2oJ8JH0JNzVu7eRXNtgmZEBgE9DdV+dZ39wkkbEZsatYM
QRH2jKjzfO2WK5Uj55K26jtlJP8go4aPFNeM/jfHL7p3gdGC9a2gbVifv5j4Tof6x1+q9TTRtutl
D+x5cnu2UISTphHDAPJBoJeN07qAHnyr/w7Dm4i9UrUO02YbfjyRhTRkdfnLR/7FmCNVhVzkwrXA
JTOnHfH2RZ9zDeHMWgEZydquaFuKOB8FCqwStzyAJkyokQk5ITzWjobuynx6ZOlOriqDIjJWMptV
lIASOr7bGAn+8GPEWF/zpfyCvC2RuLaBY2vDZY2AUShf+nKnMspdFmMF8MYCE4sNAhTi9AF5osCl
dQ1pWJgleX9/HBKflqcIMnKd0mb0b7vi37oVjS7mdpHuDPiP0UjhoqrdiMeaqKCrO7VU0lkiiN2c
lL6sq6uEN5TNOL57II6IQRQZ0tx+DQqigGQuKdhhuqKt7wkoEJS+KTzEuS/zgCjCxbyHY1h6bKjT
Un6PM4T6hfFOjrXrgWGaL5nPb7ck6k94lKNDSjKdcM4mc2hRcPuq/PqAjfOnJMYcjgUNgBYFS/v/
Euo4Zq446QaP7PToeiNJIgAaZamx1ik/snF4ZV4WXLmqDldeq819oU21ptFEzjc8MONI4vkpvt0x
3IBeWO6rN0XK3Ge0+W9UFBv3AIuLTqd+LrxZd+mMZo3M1bHUQDa4qaWCZJ+bpQJNHkNCcNT2Fb7p
WJ2YuUQ6VrZQEBTH/SJq5/b2o7IAFcvNUpD0aarYU7+BjsxtW3V9b+KKvZP63L0DhlttQo0HmqDb
y1QPJukDM4OyyZyi87nUwER/pwzyM2ZEF7MWychE3sOeqG0pm2gxinNm1b1OkycXEmFP2p7W3G/I
x+1rrl391xNohFFPCJlfRAjmG+32EwRKyrRUU3Hd7dxSwAHYdBChxqwCdRpGFg7jReLxleomPy98
Ox+FooBL2DQ22DLyUtY9C5XaI1uiKQZLFET2ueYFawzNP1kQeo3sm+FWn5Oh1C/EkCL9412JVtyD
5fwyF8o/uTQQz3mv/GEiv7ocd4d5nSrinDoj/g6sV572LOeQY63q0vx3HVhSfYBlQFLeu/8vC6WM
1JZn+KIn8AUUDBizp5GLnQH0APy1jJ/p8yh6wfM8LIrMn8wDgpFmkhHj7jzxuBhBaAninDkm/J4Y
hfIGxYpwd02jJrSAwx2HDTZX/KJJQ5tIMFP0uK/0faAP1sA9ctUQMhZbWMtllxYGiNysc+TImIzI
VDIe7ZdTX4r10lHClM9fDQv6xFhEcWsE2cbo+Hdyqa33yWLx04CFj5uz008Prrrk+GoiGaNXL3Qo
3QX4xUcds+EDujYtreOaJH1Y0r5+Ls3QTlU4GGudcir1qc07WaHs+8S4T+dZhPMjYiLcGAQpOXoB
ClO9OtnXi7fL4pfgT0qOrLiiYmYak6QEQM5pVktXpYe8+xZRROcR2RIPgzpoUI7lXEP090D6P9II
+v9RETbLWBUOUwfi+4aCEXVF1M3PLt4t+GxZtfOH6Ga8e9mSycG6P0pQ7528Sm20pKOfSOa4YCEX
B8/bJduoBa62pxAKzKgpuI9Em7tYHMOnsbm61IE/tPNb72K5cz4+uKnwG+GADmTKaNHN8M4Fll1N
KqT2wXuQ568jwgZ5Ad9Mr311XVUXPY5md5LulM/BOh4NPIwQAGW07OPsPlUPx206gkoSm2R7A6aA
R4E0pqdaENzRsMZb2TXOO54F+GkdsPE1L6PVbG7Oi0mRGBQ0Jy+9B2tpxJRQbF1YmaVgPKbovmyJ
2PzTu/ztD9WxwWwtuFMCNAb1ku5NbpMvZmkiQeP2yRRo3YHb28ojg8h3MjZHzCan55nUwNvASvkU
hImpWeKqDnKq6jELeVfdcNTv3Qq/u0bkWRoRI+TP5a8mOcPVKZ9348WwdV1knRQ9zssS8GKoZpHT
ZwQrGsgLpipQHx3xIN8JOS0C2qzV5QcFk33Suq/r7XkW9cInjk+2ONeBkvf5eReZJutpxI26l5TJ
GhfSc+IMxEUGLwO3R+D2Q0vNPIBXt/5dgE1Vvq/2ronZcLHXHEq4T1q0g1uWIBPgYihi+nNvn82O
5QCAY1/C5Z3z+aKz3YsC+ZmdAYT8thoEyYH5NdAIcLyNTXjmS6e09V/2JHea1sGCwmgvoDKHcYPl
9/2lLDcOEckS5KbEb53OdW2c5F5m8o1xIXariGLlORS4hFwyxR0KJfeK64HrLal1iZS3VBWY4pVL
eGLMgtY2HoAcUVDK/ArRTLs3i7FDqUCakqtYFTr7PPvk63u5tP2HgaGWsMSD2XcBo8H6EMNh7DRN
RO5g6O1FUQwxXcienl/mJrvMBA0pPdyODS7L80HYpgvhVUoYJ8r5lKxS41bFKG4TqKYUNXnZebQo
A4gO4dpm5Jx3vNlQKrnHKxycEiqJysjPCHqCSyVRtipiFuQAPbvdVgVRiiy6b+0ADkmEMRGs6fXY
oeeCzPCFvTB3WtltsST6gAWkjUm9cxM7v+KslQIYeNJICSpxB9FteiMKFW9wZPKkTyUqjKfvU3/C
Dc13uqTFWk9cXYoL1rWQs5GYM+uzgrGfY65VtyTNgk+BqoAQnIw0nxCrIEwNAFlsM86+zTLfuB5e
ht2pPLk7BTZw4o5Z/yQicKlCEi1Z9IjiaQ+6WhuQ8sevcibUV4jZojQB5G6NQgMruaK6czUYNkQZ
RzBRBHjtk40QeJnQZxJpAW6K4Xlrfw6T3U/G2kEv9yLnM719cr9GONBuAFgu9dFKQ9lS4wn/PSku
+PahoS/8pXhxhjBdw4uOim2WasttIqN1oGCU7eR+ZBJkxr2BPC1FStV3Te2y2lTbuBOz3b5iyc7u
ZnJ9c3LW5hPOfNd8q2uc79xKWiH5ysYeGE8kEW7Pzu8Hq5mNlGUTnscJCxxBKeR/cLIlKjbKz8z3
/nCNZhgpdZdtxV25r4AN8GLScg6BXo98JdrIOT2V4Rv4eH8izOvnsr2mXofqE2CIuuDFa14v4+8E
LIDPmv7CefYd13c8Q1MXBonsEXKwQthOgtN58HVcpljg8KZ2qjFlxMBXqrHEISJo7U34jFNPvLte
gAsUNkYVCW3ivr3yvovABFDckWcSsjJXLgmUPVlDjmi4pjG0iA5h/5/NR8+gQNB1Ey8qocp1/TuA
8/JceY+FJC7OT0iRr9rRurn4dBjODl55YZ5GIbR94mjHunEegvC+8MvlVm6nMzGpINJPEa0K4HD1
QXbTI+fkHa3u8AQquTmaEmxxS3jnww/gegW19GwbK/L5oVCffNMAZ14sKFXzhJEWo2HEvQdjqdTc
aVjioCZj+LmhP29xGLlZITPhPPd7YEYIo+u73tb8x/AX9thn1QpXXVIPiWIzW51MW2GYyTWwcEh2
7+AFlrEjl1vdyb+l4Mn9wwtLK5ph9DXBreXdjgfvPvLmG1Oix/KRUHeNJt5Ga81dHQadWmZ9D1GI
k2rPR5SrFjaG8FUxPNc8Zsm8Y+g0IEB0nDlFKorHsYr6cgiX6Qh3kwHcIEoyu4JNzjv1G8byJ/mp
h3gmjCs78htNU18523r8pNN4WIobdheiYu40mNUMeSTIIA5M6qxDBmFu+i/1khzDh89G+tKPSAAE
IIDEpsL6tTivwQ8ElsosGMsBqMw09OA2RliosmkooSnTNOrbySSnNG4PAPK2YiHhC4R5pdGURCw/
w4BNiBrF2cjzKJNC8+EwhxN8z8CFy44tXR3u9fCcAgDLIlFgpiPl42pyIg9rcPhMQtHg+mMUQh4p
r6MXohNccRIJNk8ZMB1d18wBEhhAHYf4BMrzE+Q5nTfhLoabqNcNHpSPIJI0oeQJz1pxGuAliiD2
wwM9oQXeSTlZEnAYWC5FyUacERQSSx/9xTUpzFp7LUOYvDT2LA7y++Yqhed2rlJxe0pWpWgyfZxA
dZjKJF5x7jtmq/MGcnzLQlJKuMHyG9fL2Y/EbMhmX8LL2RfIrOqCclHx0LGsm+tHmfP7VoQCVoil
Zp+LlOBSkMlHEgsOW/66RH8wlAzL7kr9Qsl4oYsQCyV40A5xUkThsR3GxFi7s45QzZzKXH0nCYYp
pEFZtdi5/qrXIEWaYskC1bNRjDt8z1UGmb2NKX/Uvp+i9Y05kRWTrETWxLoECy/bGkJ7WmBkgqMb
T0HDOwuxr/A45K2l9HRKOMl9l27bWhXwkhtASEDp1tQ0Hv4LiAvsJeXxF26uHDssI3OpZvHVKSGo
lJH7y3tobeEWxvzaFcHHnFw/Nr+YhbEt/Xsh37RjKao0/mJDUzdVSa+rM1UJmT+ruJf7eXckZHhk
Ycv4hUJVwU0aEylJET4ZJEiTsF9lwMZZ/UlAYI6Y8+9p4zksQZ8VZ76SSUs6l902XHUZ7Y3LpH00
+1iOPAFszZppKm9Fm6Jgi9gDFJg9kaSxQtfzKmtIffAjfprrGCVsmG+N6SftnHhjtQLJro2LOsXf
+svuKazQ/o0s7WgajTqpON8V3PsY/V6SiY2Sbg3NzpOssCdLol4Kp81O1mnCEdCniWxNWTqBgQU5
nSkCtGWiwBOPS8Zx3FAWt7vBy33Ku+DfwM50Ep0ZcxhVAicsJ20yqRnk4LqkjjqlRBJBry7Z2bEs
PyK9EqTYerNcZrH3WOACP3dpFgfz9kwoCmYf57vsNIEK6qeSjJJfhSXFSbOyMtJop/+SE4PWn45g
DngUPbjDjgqIICnZnBQS8sqnqm4gl12q6k3qajmMPipChUHeE39IKgNX3h1GFR2frzHzfNphQwJ/
OyqGffKFZWGjvu4qMb8sdZtPKduEncIVvFeKuQgoJmC/G7xj1reNdP5YBzeL0k7v0oqYjaTMw53L
0DHTcM7kUSF5UdEwunnJJhraiQFjZKvB1OiB2Bg+kURbFWbfRY66Ujqx0N/i5dBfPI01YIlsENOa
O30RVzFkcfzooQAguiP/PFj0ePf74p5x4zzvmV6s6dR/gCOp3ctp/FJR+LFVAly4qcoTSt1XJjgF
s4s5OjIQDGFXPeCve+NThYzATt7I7FeAJg1K4y0OzITX6KeiBDVC0lgzi96nHpDc7XiiWTlIy6wY
4Z9ithrtKynANTnZyy+diwqYx7zALS8ZYXtsTkyovUxfzN9YyiyvYeeoAQ1nfe4sIc+zi6o38Blp
hI+Y50bWRRpOLY1CMnQnVq4zKj6/ciyo9z64ekmsJ9nYNj/S0Xd3bgbYphoYUPvkz9GU2ZovEnH4
fAiQbBO4daq0Q5HseJIp4M28SkgH1pNnuy5AhO+7lwIz+MltcLK3SIX6HomsCblnK3HdfHEAgPyU
gd7KcBb/nnhqchPkaPjPygQHOOZlk1pAYmSx6AFYA+49lPgKvB8hhDYdUU7d5p+LamA6voJQCuLm
sZFsyzUK0ziWT9ZG2awbYg+BM6PQEq21KOLUVvzWhiky5vEyYIw/HZrHbt1jJyl5uTYnCqjK9Dpa
fUtNGBjUJ0M/0hd7YA4rPFEli43RBSNTpMk+tbeUwqJgUGpP4RL3c07hVbdUIaeTEaKrTRUkc434
Hpbj9HkVH+P0IvaxnikOGHhZTKfqww55krSrWmy/41oksQiuvOPCkg5+0eTvOmpCzdM2mH7vGQzO
2LBKxpNvzUaXYP0sFGxxtBKpE8D37dGM029yO7C4N0f4skkItbkf3FgrAsgjlpiM3OpmLDYJwssF
6XjtCB8QLymg18T7LvXzy0/J/C0Gxp8fcLtBJF5JDUp3aIVPHZqETzilGBTRdEhu1mbmayJEJgSB
YYeg3Xtq4Sh1BQmR9Jp7xSutzmNIWMGK4NEzt6HGvBH5GyEqwEpoWfVZtxlET2zhB1/w+KAZ1jBe
C/sDLtgQ8dhAzsi5hiW1IzX5aOjpBrERI0BW5Z1XYgz54kqE/osQZAA5EJNt04slXeftmxnDgJOJ
Elk7V3UdOmDiMxJkG+8KdSzRbejKaKJuYS2e3RANzcTX6D9NnbqAlzfyZdcuOQh7hBVDq2Jw09Sv
stiDp8+qU1OJWINHqdrhPoLTJTAnw3Mi0oYc2tS4McQw+j/Su05XX3XJEvBHNU2jpVuyKbC5Itt/
4nVSCpbhICojQiozYp7yJ8F9ZXrgRaU0Ly0kBAc9BSTWMizUZ3NZfbKofB8YMo1Xn5v4NlpPI4A6
jGLpoX2P79G5J1vCMyS0ebNIniPvkKgYlwGxqGT8Z6tUNhuCOH949InUM3M+zXEMc3V7gIOMpcHl
M/7DwQrvTli0hbaoDeDk5Q7zU2XZRelpdp4n131OO43nxSS1VkbX8vHYHXodlCsUM7qtzmth59sT
eup80YVRD1JY6atLMOK1T+9upQHSJ/2o7bcH28kTRszqeUgBJx3IEo2Vr5hiAPlb/wTVctys12U/
OYYDviBh6VoUHfEGoo0Fe/hXFATpOF4H1j5lwCoHXHs9Fm+OHuvpWIVoaVcxFBGCq9eBJWSnhMSx
VshNe6knJqKT4pwFnBlmb6nCb2SJS1o5hhPvPzPRfq/3ZTakAMIbKEt0CUGcDucHH9YRdC38k4IM
Z47V44s082RrR1O2R5n0Ezn0AqRloRqfVBjucJBCHKR1xEtgFIBIckGjHFTGZO14U6NPtbi3pSlo
ROMwzhtp7mc/UVvrwf1avmydk0cSjILmVAoLckEHbuqOzGq908Z2CC9zJeNrXrwI3zMVnWD661ue
teKawCKBASmcHLtZmtvS+PHwFoGTGxwz1boP98XGSPSCROPqvfFsrQ6FUzLMOlFmqDDuC9vr7Vg6
Sc5MsHflZMgLHzoJsUBebvsDuJ/W7jHivMXgBWJ44rf8Ba+hTihSN6ptlAqsvAgRS5lEPRoZn4KA
yZiWJEwpm4yUrPYdCtCzFgJjwGaTA1ZDBHINH/LlZ5lOn5WRSxm4N6qCjci9jT54ZRO9E0WD3K6Z
0q1GBzTiuCHvwF6EHydgTPnP2QP6K+Mt0nINOMg93Mnzk2+muL6yAOy7sBIanfaVB+HYAPLHdpJv
ytb/8XQ/fcoWPsuZU99Y6VPbrm/41GZjRZbeNCje6yMErUHFTATygO58CqFIdNfyJbYmPK2WQQo9
+VXDGDujf2rCaHmidclRM1Yk4RIRUJf2oBKCrZbdMaw4s+6WNtHp/p6+XooYJy48aAR63WZxnr32
7VBKlLFuDOVsofwiIsbAq1RRB9NFccYtjzJmTafJREAoDisI504qxg71obuaYYnkxn3uoEU53oxI
GExDrQXyMDIxeMZ/fjN1FCXMLx4o39YG2ZxRnhvDDkPGEoQY33x6MdpRxKLFXncbdk5Fx1Mf5rCQ
66kXoLFroPLsgPGJFcHMRQG0A3QdbiCEsOWeodUqpb0z0Kh+uQXbJrjM8pL5yHyE+laQB2QnBBJs
mj9bzyoq4CiMBfRGZwhdAj8uXxlw6o8IshL0d3bekQwJ+hdtRkcqgFERBaHprVGvyWxT5qISRMfC
cLLO4HsdQJXR3J95WD0nzGHai4KWYWP7Iu2qiIpuk/ybob1GqBmwQRXcArtE4hk6wqaEaDseB+jj
ZbNDcpaKIr8hgE5KaBYOHLRpdlts9GxH0ZxRko3PMhrJ3J7/3PHDyF+omLhWN9QZgyr3sGlhnUBd
6fc8FypoqrD5EFqSS8sSLN8P5QlcdYhG6wGS8o78XoWZ1xLGugTZgz21Xq90hbWI/lEpoRLNcrCT
11lKI38LdMmRLk9Hf+wkIrcxfyvYZbfsP6EYPoMNtqjJkYcrfWr8I+dcRD48kvJRpCynaIXoFXBk
XVpc7kXOlcCbYQ11vIYmalSjjd44lIIEtjwuJ1CmkmWRA50M9SJkVf4cZPo0xL+v60M62i6m0G/1
h1rthtXlplMlDMYfCFQQwE7hbMkEn2ZR4y+rVFEycplEQfqCFVINTy6Uv4HzzrKoWnt8lYDqQOsA
QxMaP4QolcFVkA8T39T7kc3/w1YraBTL1alW28LcFmvrqSjbOIBynY4GBOLXreeziC7ZvTgl+wHk
XpRw+lsdPeO2WKU91ctLdwAxtpog9XT5K/RXgCYF/iskD5B0G29k7bG8MZ8JZZL1uIfdCs0uWFsF
QBjy465HaietJP8i8yr0d2xBHrHIzam9jRqcwgpqrI2qkX85JrWyfBxMcm+S/cm7Qoj0JCuf0hB9
hqk8S8RVFRC9GQ9M0+8Gsmn/bnwFtE9k41zTGQi5JQprnDa0ivD740xveUxE+13tQX9cMyiPvkcE
hYRGloGpSv+oVszbbi7jbMe7n+cLj2OA6NEiE2ndnEODXOLguAkR8/AiTJ+3rkeeDmEhqCpYgSg1
367iwr1rqjbeMB+6wy8aLUbC6ZRiMQTHjK+nPknCh62mLLvVY4bIoL3vVjf7QCmbBRux3t1p6S4P
f5f8BTxOwecyIDbAeX+5KCx5hWRjwWA41WCLZqepdgU8akoTClEesd+rP/Jxjpeh1WA2byjpTc0P
frsu+oFAx6nJ98gX39LMs5IF83rlasQg7tXd/NCFiUebpU2x13JDwytCXjq02ECIzzlIB2PckPYp
yCKb+KB7ZbhtCexjXSUtnHU6XAwiNn5vC4cytU1TK27Uj+qcW6Xxf8D92tT0v27tafjtJU/ruyK5
GtBWWLMzaEioC23t2OAQ5KoFQmzMVyqo4DXWtveNX/xN4vGOFIWZ14xkit+3BaMCw2K2+stHV9KR
lVbPtpgMG+cWtRAqJilMtL5ATN5sY8wziPP5nyvneeKrJVXVO7PXN2p09lFMsYUrgKCLoWvGAtFP
4JHG4ZdTgHNZlw7JX5dipS+eYxry9Gavq3v7q5m+R0tFlkbfQg3jCCvL/Q/R3gso3UuyPTrYjIUh
xDMZxC7pMEeuwVOVrWq3+idGXO7tUkWuEu32LC7ei5cWeryA9ygcnlnqts3Fly3AtiRvIpIxBgGg
ZM/KUZoKbIk82ptFfpElGpK5vGAxb9J29IL+Hzm9eL7KNDZgVbCMlgkzuGu9Ao/7XCSLRYR2i/bG
iiSHN+62SyuuvzfxcYN+6WHQ6COZEr2cVRjJ7Gk8+j+zAdJHZ3zwkzWFqWg0jcHf7SifAaAthvss
yVM9j8fKfRrVEXgldNjxyHai98u0RZohwddTPdlzdBIYmcZ7RBStKsiq6aU7jEEyCgRAE9LGclmV
iSbsLVDYmREnXSuAjevIOfscleMCSYKra4+9utT632YxcqiuWsQsaus6PqJimDbnc6xfitoJpZRD
M8Kk8RP1D4xKgyjXG6OxPfjVDGbJJMxlYk62GYYSE5maIPidwSLzT4tpXad5TNBjfTgYuTVKMInY
mSoO/dH4e3NXdL3F+a/fZR7A1L8=
`protect end_protected
