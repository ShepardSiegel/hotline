`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZpBx8GbvMBGX9hdIIgf/H7tEt5mUQNPbV1wbSJloGY+CK0wJW7i0VgOl9AbdeX2FgXcJ2qzwIKAw
wzGL+AEM7A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
l3z9YAWfccJtsGZbe3mO3omgW5vjtQFJPlIemlVOcLM+FkxIx/LoF9v+sceH0zqLFT6Riq74YQMV
DR6tD0pAthRdx8avY0Apfj3eXKTFu6hrY7pjt/3uu8E3JJW8wBfYmZbXmUUP+9PeWmTZlBLPCc8N
dddNXK+Gz5M4xnNyWUk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UvRtbXXq6rQ+XaV+8S6i7pV/T0b5Q8XXCAFN8a5NJpTdl/UaEoEfn4sbwdyzm+lIQ2FVjl135lD2
WfVGANU30rnBtjYF/+k5VLC7H5QxgYdLV2jGtZKrL8/DXHgFulKTjJZimtue5AHMCh5wKaXebIhx
i0rk6Xsmk77yVpLfiqMNMc8Eir0zDuZ0HHRkG/0qFgilOOG6axCaxRJWeqBwL7oGhwC7GvkKqBaX
OXtjLuCfVR+9/n+qK266WvqAYTLkg5GXkrN0pUdono4x+Vl5SmfMaKP2embd4plIM6YOF+FMB3lN
XsSAhaxPHqWdnr3ndcRvjrmGh7LT/rwlxXb5aA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XTB55km/r7NBeEJOpt0OK5z5pYkkF9kI5noo9cyO2mQJvZ/XtYm/87uIFRFzy7qf6EAvhoFjTNGO
hAU3Sw6Z7+ggkR/LxUauPp952XkTrn418IFOcJzsoHlqY5iuiA4fl0cW6FFPO317EzxTU8jjZrvc
6ypV+Rfw2uuNZvSYJC8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Df/WRXSBwmiK1ucoi6JQHUqJMUrtmhR2pgXbYgsREP9JSJYnbo6mxQbiHlam2cxnnbWK2eO0m1w0
7ogDF9JHmgZT0zgQrp7ykyNPt3Fuy4YYZWBVTV1LP646z+no3B/LxS0/+47LGe1Gx8qeCrxCJqpm
LiYbGcI99v6zIl0MNBTvTTQbgB12vq+MJRVmkQDm4ZRA+/Xk87hwph3qggHGXMsIFhoqHwcDMBqY
nQ3wCm3nJJYr6MP4q427gZIiBNFsi5T8Zo3JOleU8L7oSuorE778yFThymT1iZcrDal2apQtkd4p
jlkh3rcNXGLK7WhdUxMy7/A9BoeM+W0FERSYvQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 42768)
`protect data_block
YC79N75Ti4ajXrr6kVNUxpZJ6L/g59azjpRFaFG3NZ6A3544zrQbMXBtvKJuaBDbUpTYcEJ9Cbpe
sg00YcKN8xF+whfvYmyIzpNW/i/VDV+rit5uqSc2Tbg8qVwZm0l2k0pvANIQTJtbLQnHeQIntETx
7IHDULb1GH3+/9qXo1p8bl1e8VPPOzD3oa7NVeO566a4DQmVn+4BYHwh+7s/PaOifovkfcoqroO+
C2n0WBCw7WRbUDwBWvF6CdjvhfcBql15YKnU84bf8qS5cwhDxpN+lJ3ty6ZvH931uK7bRGlqIJbS
JhPdcyELB/nMiWzKpE1oQz3O2AJ2FyGrsH36Ik1Peg1LnC7iNBypjPMySVl5vHMFtB6mNFnnf9c5
pLBNhubLTSRSH+tZV17BHUDiG5U/XXWasXc2KhocbKg448vS86uNSYVhggWI6I2qcLE2jgXsqVc2
6zk1rvOZJYtn8OVNGFfNg8O6gJnLmMiHwAH3CU9DosrXw/Ux+KAhJFDXhOQdCT45imnLm5YA8+vu
l+iDYmZgueaVAM8ixonlsyat5o1PH4mdM5MGQPltNQb6TgzMeveZ3z7si9yHwhEg/UkJAIIL/xXN
mTCefRDT5JUMsFoBDkUVQdQem8l/UAhyLDGNIGzVy8Vs+h1ZpwEBguJ5ARszWs/TMzQLUIQTjSX5
iUg0VH2aABFLlF2PKutKJzRhYpmTtmQch/v3423km7M4kfz4n40GgmecKbdARVE+NQuU3k69oQ+P
2GJzQ00JrCOEl/jNW+8yTh+jf3xMZRC5b7Wr+WGdrc4siQa9clk2wG36A0GGsyrWRmtzA5kVibRY
SrdIM1Lnat7L14x2yuUZ+VXzt+nPzPCutLFaY6YN4NouBLYZMfFceO8TLGmsjnpZN/+LSrjy2mvD
e2ImVczqThMZwaHV8oqXvZa9l35/4a0b+quvbpbuWiDhb89OCeEQ/K9RKJKWCpBd/g2b8eMx4zhs
zmxwH+blj+0KQo8vkwGgCBAHECbNItTVQJFt6ZWqxgKxev1/uI6TkAMUXp5DSjdVd/mPXl8kHdHn
VnvMPkooT8FzU/bzWj+iALmosR76prdjMS6rIFKmELVkL3YkCm1QZmaHgz9IwA4kfKr5Nge5v5Xt
v416dh7UGtJMwgkmJCwD2gNLKOsvFkuTSxgmyDRVH+W0FDhdtHUM/PrDgm7PoY6u6W/MFNoCR9Dm
hA3ow/3SclouJwUz+Kq+lffpYvvyttq1ylVR2DG9ZoNaEq+KXtewwtgDcYriE1E6tVa3SKJC+Tn6
AOah6PuHoYHhiLLnBQQinemfS6vKO/BmedS4fsvIyWm3197sqhaHTcNcrU6w6g4hjPLp7mleiVFS
OVusq5RijQ5yv98K13TKvt5tvkNFvLd9JLKMhrK2zLZ/60IhE5w2g1peXzHesQJPpT6Kig2sg/1+
zyiVLHTuZSXBRsuQ/Bs7FlYfCwC606FkjljUPiW5JirB6DIw2vm4gL5cZqIGWes6DQdyNrJGALmn
+evEGVYi5O1njOI3r0m/Zgh+qbB31ATLCRVszAYbDl60P+GGCcQVFgDn7B6Q/X0EvfVVCnhigdg3
InkNqPNDH4SW70Cn3F6ln8vnl2VVwgUMYkTAUxWlORU5ROidRrKLjgBSM6kWHXTz/b84KL6HTEq1
OKccC4RiwsPtuO3HSl6MTcT4rSKLyWaD0QMsbEGpmP9g5lxeP4sCYjumtgoO6N7jSu1GVulLtTFi
jqk28y2gs7U0N/OjRNVqeq02eKB8CeNi6GNzYT2isXkuocgWqjOs2Fg1lbkGIb03oELRno6Z/EGS
5FdaeQ5Hjii/9APhG3KNSPirIcqsLaQy1S/zc/lZptHNgrIbdcgYk7Z51BGLgUFsTGbCKUQ/Sw1P
16tRA9MRRUJ8tGPwvFlNB9Cikm45V07fh/Vejq+yo2y9ZkInnALHsppq3Ry4hjNU+28Hb9KeRsg/
X0n3wIjSQq9lnbdUkfRc99xe8N3Tc7Hl6EswrO8YhP1/BZwKc2Rzb/FsltLutE/KajSLUeKyyYKF
F36cTBCzG/iJ8t83hUA7tV6+o+nGbB8spiYX+TQ5acixckMGZjJ54tKfmB/vyeKwFlG7RU8u04dL
Pv18vYdCesm6mCm9UmsDgMQ5nAiIrcgx5mxrv8e4IObsMx6kI+YuZZ2P4n2kBZrDc/ZUIyO+qxao
+wWhy5Rn1jTZzjwct1cQRAka6N80g2yxd3oi6hl3h+9qte611BJYd5r+2L4zagQLdkzugKhUSv/X
YoGzH3CtNDa6Ua89dYnd2RjOr81nUUp4Ckl7L2+xHu7KXEk6JZ2rHQRDKJCblp+bFduzAKsgE+wm
ZB4AkDYEYeAgfaqIXJkOccF2a6SmbizGqtTzQ/7kXwDtUxB2n5C5Ktz9LW9IiSWJCKCwjCPnmtSY
/Xu2nG3Kgf/zB8uI1vK1+AmEp+x+7TXZfjXQHGi4+byTFZTnA7cQYXPffXCXqZMJA6cwUkGXCrAt
lz4aJAC0nN5GLXEnlHo0gh9OJVACpsCRIjpHU060OaBljYY8jLlmZH9WpFUEjsHP1A2Qj0QJthjD
DwHz9iHcUYu+pYXVdSC8A8MzU5ustR6IgT2Dt5PXRJSahkfKf9MKaNAj/OZm8by80eIA8AkcBObD
ry7l3I4I5hYx51MqzkJBwXqO/XS3soaVQrpv/8Hb1k4VZBl6xREBcdbHkC9ETiV2Uu9vV/0I77Yc
bmNzqIE8tyy/7tEzRY2ZGz6OTfOnRWwSUiA6fMz+iSd6dERfo6is07pnOwuYmE6NFBllXdGkDhdh
Gy+LeiMFGvpsGoiOfqJXFdj2467Z8h9OUQ2R/jkYbjlRAREcIQrIYfSuDsH2We67V5cSYx9NBHVt
tcJ95PY+kDt8Udy4lA1xWFcDxAnjftFx6CF3iFGIau8B+PslCZ11IAzBMoSK4PdVvoafI0ltnm2M
QZEco7lxqas3uDTPU4KePX1lNYnQr3aoy6qDMxaZ/5af4ODDO2Z3s4oMCZPQpBtW3QrRHM8vZHRK
MdQZgoHCdFQ4rgtjei4gzqQkZOfe1oiV4PQfrH0tJEdcz/aLHwXtH1JbeArRALpgXqpkAkIjQxqz
02b+/uiPw6jyXpuLqfUpNbFUwctkZXRUEA7TdwDpOo4cuiMJJklSFB9XZ7/97hWIkwUxONP/33Zf
5uJjmjyqWhq1NUfaSP6wwaP5NZkxHqPgn/QHOnZZF7/+eL45szznZKhGIkdLr0c7sG5TpBqHokJq
7Hdc4p0zfdIMUi8FeVPz8vpR0nT5ZpGEvpZ0g9CTYHucNX5qAVoNbDSG+AmP1o4nHtsZC3QE9KtA
92qXKETdqG5aOBGta4MB6keLo9fkBFd7EWD/5hM3IPFJySvsF5FZiiSTA6K+6ToFCVb++L0qgrbB
ncAN/MNZqqwRBRmrniYWET0yqChRZpEQWNfHrZwdldev+bg9ecaV2iPI5AZOPHiZfLnRnQGGxAkm
A7SgjVrLlN8RJrlTS9sVMCgVok/lrlkZ4VNDw30t80XWhxTMXINKHUas4BzmDNX0GUdle0SgqXeb
m4pAPhQ4CIO6W1JxCVu6mW2JbojEWsDyEsQlPiDjMD0tCZenHLn0VnrQxnvKF8Rukrx8uLZjt8Pt
kkW3Uw0zdb6v78qOBY41GJq9UymwOpgTRDeLuaXuDaVBxR+U4Je+kln1JMiswwKITf0l2DukLbxY
277/vSo23UW7jV2C9NJJKjfih5siRIDGqhZhAYmqjQqBdWfyXUv0yV4iQg5a1gQ8XWfY5L0Ha847
MfnSjlkJaD58kJcMvyrCEPl7w7yu8iy4ociIROKbYrT5aY8lXq1yM1R8m/g2nBld/9uW06XvbzkS
cgVt+HLbuEgEIO8yCIdQljV8oebne3VgKld2uVMVH+nba5pdB+H3vfhz05wxwN90cqt/p45ZrXym
MbIH8KRrTvmb1JRnkJClh6XVy7CLgY83mTLEPlX3erOLLaIsZ7SlnyqPknkcRTXvs8Y65DyjBAr1
AX4XGAdlJz6FsHd+Go0AWjP9r3yOtkATHi4K6Bo3DT2afWCGnTbqjnY7DaiyFM1Gg+IJ/Lx7SB2d
B1JbbJe/3q5ji9m/WHY5kCvY0VZDAndthiOE0p8uW5LyIEhab9ghRCIECMZbXQqh4mscg2yUfyZp
S6eqx9ACN/ja5QFu18HSZU7LUEEycy9r/y/9A4UM0ycwInTKQa3mamtsXr7DvzUANInlpRV+NB9q
wNPcX1bxrbHaDfwnHbMmX5urEdIUAvrNkFfDi9WptWBeuxjqb4Hyo6Ff5XkbgyICd19vmM0kLyxG
eG/byEcTv1jILxRKy3ddL/AzV9Rfkvou98Du4cezjPIxzOesHAN+qW8ISBBqc6SU2WIzQskgzMwQ
5rvsavWhlrof+84nZxyWBjBMHkows/YoeVoe9CLl2NCqzVb+a6/3zC1Wk2Q6YyV2xmwkgGI66fyc
uRUwF5mbGLGS4WhgfzkNw1ANuYa9x8qk/jbt6e82TFmc5JMVB//FXMynS3h2rVe3S0FPSOkZe+KG
k/ICfFxWQfmXmHOtwlrdSTfJoZsNhzX1fEm5tGIitSWPQDG/ir721YDgIIA6MeTKYby5wO08q4Ew
oysGDkjiQobBRa6C0gKCz/RNJu83Fw66ztwZV3a+LC9j4++2SwRUPvE9wbpFN/Hd8/aDGQK8qtA1
3EHl0Q+BRe373Qm5EocMiIowy94l8zsEVSMPLYhOny3u62/DwvVF69UclGJrfE/vbAcCnXTVFUew
O1geol5mb+JxFMZCe5ZaShYhUiRybs863WIBrJFWtUv+0mtbMYhUqICpd148wrAovFxiZqoOsvM5
y5p5ebC1TKyW8TisxEHF6Fn0L81B3bAucCb2l2ClD55iUp2kjcwmJSHTT7n9kUcyfQI6SmYnTc/M
X8WGuyxp84T5gopLX2I0nGHaRB21lBiXNMV7k0/JKU7PZl+OKwOf5Vk7q5u7acOVc3+f4R2Nk6TL
WFOJrJBLc9oTCWhTE1Zc9j0Cf4rgQZYcBT7bEiMylRa/THLybElbE+xWqAxNMxbAZ3HRTc1iIf3R
BJ+UH+BRGU5aCp8du4aZ2VRbYDpcqQEiwedXj7I1sq2tpJDwsKGqEnFfKmuTKSFWPDk6mWvYS6MN
fMZ5IYK8idiPaRqcZs0GSxZxyiMNT4qpFYcPMDckltfSViYnMtvT5f1/06EleaSRdM+j/NxJ31h2
ZA5/GkEs+qJLX3L6OFch9aV6Oz6xrtutNMmwrnGcZnEgrqEm+jhJdVfcx20pizP5sJYMC4ptG6kr
0U7WbDc3A8JgCKvZehHJrxlGRfyxkxF/9xyoSSpTeH8Id+6TsOwSYxkaIbVVmX0jLr/lv9ojdv/W
kn2TgHasdx5Ov86c4PHf/x1r6Xa/DY5kfN6CVW7C+m6Cez3+D1U8pMlLFL/tKOPK6x371j9HZQOQ
jH3sviUx7xwR6VYVHl2eKLIzxTOQo8BzkTGS6BTl2sOJ2Wa17e9+a4HjltOaHgyt2udRYePlvpl+
sc9KqVTrGWOAI9jnXAnAnnTPos3AF1DqYh6SIlaAYra7v5j0v9t/FtuCx1Dw4JdPSbRDnTZEQEZu
SKGEYP0oUflMU2zBZrg7m8k8PXABXvjXvSdRmNSg+q2YmqXAOuNvf2UFKyj39M58TmZ9eyC8kx8H
Dq2ISgea95lRtSSZ9RjRQZibSw0PdNWXqBE7WbpLQVtWkdqdCOyiIy+PJgZth/1TYMTodtIJ/PNS
yjCethFNAxvGjbFvN02UwaGV8AdPPtGX6jSEDDXu+QJ+8fPbngNpbAHq5ltDNepQdixlRzjCIeoq
qE1qB8vbhWPDcqIDnjdY8ZEFzoBmoZo0/Fp5vU6DoCl+9j84kqyMicGOauM9kfkKBSR20Z8cnZW8
wHAv2R31LduQ0q8OjAhzFA7J9toNYeMQBbGxjcvy0/pEJcO8gF0jH4/GgwMuzKHFXNXDEpJXSjnh
FkWGBsFL/M0eed0Rlmm5xputsmf/2HZcVNbJsWlBAzZI+HWq2/aANPeTTl/bv2bwHSDQTpCAXarQ
yuqJZ01w3FEKaPa7y515y8FH5YN3J9EeaGDaeNEdj2dsNDxvQ47PEcqnbbG9VxoXf4uv/UFlTS6n
4yxwiFD414RwFkU19o+VQ0twWOmp3iDaiUrw1ne3HLqKFDDvgdjbTGmEiXCAFEE5GHiSfofQT8YT
y2EVO1lEU/8cRYYurUxlt/zUIlRaC9CHwDfRUq2DDOmWMpSsywM5YseQpdmcpkMmn0kEoI9c7z9C
oWTUaWnhDE/RWErwt3/HyF7qfA+jWWvAfbSqhLY9TaieuifI0Std9oHOEMgHWmrPb9a88Gs+3gFP
O24DUo4ltSMuk2HGHysSr0SINh/2nxn+hFTVG6MKKX4UaNuC/6Wzm/42yVDAfwWbgIpqtTAVYSmM
HPQ7zZL9gcN5smxgnez/8kHIaWHdUxIigrEfmR3ckCsuDP+F7HQFNtGof2zvYL12/4S4jcbZm8Ym
7QC3yxzTKF7KoDuhilyupEIsoFlqjE6eZMdaF/8kJBvGeGBJIHuJiSmTOj1LECnvWLCoP4IvYUk2
THHcJPKJ9lAsR4hee3tfKJ6wNK8zwuGkztX3YVUsWCK7X4NRrqVfVmLlEY5iV3vAHNJuYkiHtvnI
cxcJ2I9LatVtGV+QU6eJyDNz5TPLqc6BmAbjfJmPfHKysjDPMsIDmw6FSQD2Z7nYP2ikTxuvj/F2
7jxnEll39GOHy5vEh+i4yhbiCwob3hHwnga1mlffrQ4qgGI24/F4NjElpnnD0FtVMGn/BNBPGugn
qfv/cUMO/UYHl7whAC2OMfOM1y375w/cLl6ER1BSVbNknEC+bOPAUPUdrqVSFeZXCv3lrT10De98
uuilGCTq8dd86lxspMVQqa+oRJXKOx/DQpBizmnMsYRngMHckkPh7RD79APufK6jv1JaLK8zDc8d
W3ir76R8OOpQqSYtdvkQg0uK8dr9pFzyhuPdMMJpnZRk0wGoInhCj9xl+616uQCNVUe+qQjAznUA
6Ku4p3jaTp7qLZu1sgf2rrBGpzsMy8mmCp1oL3s0PIdWuRCxnkSTRoYBWXaRQGjPZ8eJ0cq7/NaC
8aqJYxeYL1vvSUSlkP8dWhSdBWWbFxFz6/qWFNQLg7NFSvAyLXxY2n2vbB+T3XgZGF9s4Z2eUOZF
oKFAMy/CLEUiSgCnrGneqp8mzBSEIn1M53S9CYvpvfeg6sLHOHw5/AlijpWj7fg2EQRCps2jMync
yFdPWVk7QYwwBaVZkt7F2irXj+VEni0yey0Mgysl/vmVHvl3nC2tWgWP3imLgYYwBrEKDAWq2Khc
ANFouqrvhuzM8s8U90QHXtAPSBA7FCMrehU0xAKJW+KlJpjN9F2SeeV/TO8efmeUFYpYxuwXjH1h
vsWXGiCjDOOCrB3ijVN/LSzgGwEdqVPlzTZC8TWsLk1F8uqt8N/3GdagCBylC6Y/5O15PK0uC9Dc
xvFqK+OCRY/ozqRUJxto8gqNZsS13xtMoYeiGD6ysGsJFztqxC5XSLicAs4jMVf3W2qWSo31tfSE
u9UX1Rbm7kqjyc8T3KPgROC8URCaAA1MhjBJmug0+BzqPUOZkw/oetRItasECSQHd6jgmqyO9ZWW
c2DcbWMRhF68FfmZuKTFZWui4YKkdSwndalvsObMPG0VNU5klzOEOJS+Sg13T/guLcA8DMipnKN6
sK59jixa8TnnAoJsDcrzDCKEyQTL+VkXgR34szWXE7m9ZlgJBYoGtc7tsfSd0CBghP/+VAU7Cx3J
BHHb3HYrA3GOH5iXvGzLEtnYKQPwf8Ch7zgLVzNaTrrJNialaOLIZoD9Q/z/5JHVX22eoCeOd5g7
UzQa4Oqq1QoTNhppUFgXbJQaU9J1w9Bs7yrdty/dewKlQnbUtlLcAoz6Ls6wsf1miwVZ5HYCgBbK
2HXxhI3/6NtEu+5CtQ93eL8JIzsY621QE0fnx7IPrFN2XOZqSgaFSyM5SZwLsdufX2x7Hq+7t/PU
VIacd4yZzDbBGj/klfKq0POsJTWUjLmckMpQsEFr18hkh3/E8ZpTPpa/1bia8zMGUqrUOVMWTI3g
8U4vhB6vjS5VlFCeC4pFpPiGyzEYYJ5TmoODSlRLuTv3PIL+yqFhKpppwh66RFuEo6/srfjk6kNB
hLSYRgFQw037WflRMIdxOwKcuor1vD2AU6mdFoFGMpMcVoE5qhOlVE6tZ2D5MMquCnQfYBWmIF8S
9x6iBCVsn0QX4X69dmMbIZOvqZZk4pYcOqiAmsyumistQkkoPk5Lg2r/c2uI2Z96Jd9/AHiLM3N3
0YMUuFtwhCxWM0DpXqlRi/+OE6e+r1w2jnrh58852QqLznyFTQh12oKbzxosTO0Ao5LpLMHBJ+wt
GUHs9dh+acxdCqXoXHbNXpgGQdLpCMma9aRGPfbjSG908cwSugo9j42cA1NShavbDe3JWmrLgt32
hPLcH1z8snc2BKHl9AeQZe1aNg2MoZZL/YtmSlP9A9j8MxT827AG8eq+Skg3VZ/fsUVxwAPrO2m+
1aJsqqp/Y5RRObmI03IPxVCWO2RmKdYY1YFqDW7KHRBQcpOwatJo5mCrgJP1CNiwIXSCk4tUymeO
jyiGvWcumZfqj7fNqxCcvdU/PBoOKUFf4c4qDJHvD+HDVaOY1Xy8H3jOBMEp6dUUUnUrP0NxUBIH
4mpB1unclg7LCOGIfKABoHIzrccyzp7dA0KRu3Lz/GJGXmDVzuPZ141IsVZPWJoyarPMmaemtUT9
ZzF9q0bdOb0kwmPblOO6ZytfjuswL8pmkLpWHYpESv7x5rmMjPJMzECeoulJZgX6hKQb+IZWS607
WXQMort2GEvJmz6x6WyYEzhXDRmvdzsrOiR5j08BdKsppz8U/8DZrDabGSrNy+D2Cr1HVOR2TyV8
9F3yPMeeNslNCDLAt7josmqrc8QehSDFbHZnBeaxo1Jj9fAdOB4aG3+W2Bnq2pC9HsFMpAKGb6Id
QtAvCVyN55a08L2ySMJgVx/4uQgTNi2R388T2WJAyebMjllG+IndiG8Iaocsl47mlpQSzXIbca1z
4e1mUkxGV6HAWsb0/UzpYqkgHLfSY5YHiRy2dtDkKkbqdZDLxWHl5FJr4tFJ5xKOf1QkZbliVbzC
5OwW5WEPKlSWwBhYheogtBijKLXOvh9jPtbaRzw1E5m6TAtkM1CraaMXKEo3mB/hUXlJxcG5HpkH
/FR2DoTYL5mSB4ERdHsuThsvR1KcOWcmlSwLuxl97vHbTeHjBcMJAUMBfRgOoDS++hBprsahaV9k
UFU4hF8zbc7ZE26NdWa0m51TQEi5hSsyeprTe1xL67tY4RJM+Zk5M6wT2PgzragDMmuND6CCuMD+
3g2bWlBikex/apwnGM4ZHnoPhQZUZySDkoyYnVlwh9kCJE7pdkWJYJylufZlU/tnbt5e13Ju4aos
if2QXQBSegTeL4igaGz3oZZX/wF7PYnuJPNdX/WIN3yf34tMmqwkEUxztelMFTugjrEu7q/VM3Ud
qYJzFhEAjEu/IGHQGKpQETWggyfIwJQHFBHXe4JkWijD6wj62gXE37XrMsmHl2KuCvLeyXL904JU
0z6z8Bm0c+pv+hS1j4nosF2WnMmai3lRqdWmxAWzjC3VFhrT1LBFKgT8QcOLBH1Hkbrwm6TBlKZj
oQgEaUYm2hZaojWJgAc5Hqmx4QiQxF0mzgQ/KCbRooHvQoH22sSNaFODeaGMMcMPjIb//c4qUXPo
y1hDrdlazjZZNeiznvhC8i8kXTy/2H+NUA63HWspLctXfyoZ117qTzEesPDIew5r53CCNZc3Y70M
XxXgv3w/H/mmjSfmXlrP7TxSJ1lj5+x98YAkLJEVkOUYdaOL5tIMKX8BRSD51bcO3b9Aztxdb2n4
uY0XDay/BMcojrISt7SdDxjQ75H7pE+x1o5Dg1UkrEQTIF6o3OLwy5UxLNhNrNL6tCZu5tLgqADx
sQwICzkJX3CiX0iBDI9OPvjSLLKazcbmYO3k/O+4w1Rrx2vAdkT+T87D4q3ctopesmqnq0fXTWfn
2EGnu/0TWaoZgoVXaLR9VW3PbaFBeQhC5xUressB82gXzlzmG23KKXLOxmEp7ge5dh02b1X3iZXn
ezEDgj5XHRShwm/ar619rBh5XDEo2aIdVfNEoqnvyCtG4QcexTo4H8yDYITUeIyRA7ZKtkwekBfa
cm8pZQopgxrBCa26DgUyFlucpTSviBgGJXR5GGWwH8dfiLtZKFGv/yngY0FSk+wcVWkSIz490pMN
eWypPxkY3AjTeyNwiaTznn2Z4kN9F1C1cbpJkCW1GUhW2gNwcopcR79Wrymd+f/5jet8dkvnMxH5
OdnPhjLXgodCKENMhlIwY3JgkuJ+TJ2aPp8aGXQ+iw1CTJCFdOolaDEnsgAoSaqzU2zh4vw89eDf
PpXNFpuX1U6rVzVbwYKusnAbqLhiqg1pH8VXK3Wh7B29jql8zBaRH0M8JTzWSzcuR37COZ0l2BO+
eX0zbkFhsyld1BZkC1/6A7eAsKbM/+sN7Asix85qCz15CgeDUiSd1Ti79fkxplB53vlNA0m78Zao
/reFAauufVbctOtxNAe+9F1gGjb2rMPSLve/52M+Dzf/OXT1qI9qQ8yS0sdFKa3KLP2BzkFwSZAU
XG2xgBZOzAywYZU2hhAr9/u8GfLsZpjhbNlYDIytzGnZyW4cQilWv4LWz3HELNqIA0EgFOkPm1OL
ozGCyk8ikMdL4+7K9xzR9fgNtEvtJDWbvPmUmeX9PRDfVt4LCv9yUpGDuPMttcpMiyRF8Pr7aouh
QhOdXKKKHfU/uQjqj8aEgpyFnj1gAtHuoiRNUm9ROmahMsfYdBasPjkpQw4mBeP8tNDb8L6OCv5l
51QkdWSf7d45nJeWrlhH9eCRBvX/alpp7NDc4ueui4WLg0IM36SMJA6LCoMNeTwARR0M6foguaf2
i0adizdzF2PwfUsUcH+MRkNLKieqQoZFoEaXp7cNUXx45lZcOa3G12Q6hP8/jhcBZDkJuSmQkrw2
eZLeviJehx3GWP/0AUk7FeewYIKZTEnCNj/Nf0OriqrZY2vVlAKXFK27eqIwI9feHNG2CFE9AYe5
a/V/wnaliKuasWRaVvMB+cBSBc4/PHlVELzePzcobfuN2YDCzxd6Ic5Kn3BypuqW+BSJmdhFpnkB
arYT7/4SmjPKri0XZ3EQqLBt0GkuK37qevb0RN91Wz9N5ot1mHZVJTn6/Db/Wu5oEtH+b0KbQ9ZX
8OV+9+lMPrGRwwtsaQ4o9JM4MSQhgXPl2LCzq4/m3DyfUDkNiySCHdWxvQF85+T10Exr7eYMNEw6
96lg7qGw32LHPE3Z+NF+ixnkxbM7GvAn08YGpMKCqrbph41hZLZX/R7sUu5aCI4I190sdkfYEhg8
v4hFzBI5egu3+jrR0zUc9IklkgEv/2gEzrjjQ2i54fWFOwB5GrF5qiDlv8DuCSNY9MN1ImYmrEoN
EUnEXz5pEYICacINOi1OwxtmCdCWeq/kUVR9PGfszmqsZM7X+qaS8dTp6boKwbW2HiEOdpHwqt81
PERvT5bf3SMmNUl/h1B2YwubuoDItwmketLXeAcbo9xbktE+3F7V8wmF31tdvu9Sz03WgyA2hdF+
gauQKn6xtA2mgpHcptblIlZjkHklrBaZc14/dVN7E6Em/b6l7eqcaX/ynkC9LkQzZDgKxZkqiskd
wpESFUNtnS7oZ2G+sX6nnqEQyIcw+pRaLB81Y0lRBtuo8hROBYO+r9ErMDlcl+EwFymUuVp47n8Y
5A9aXU1VqMFCeHyK4U+LlboYS4eWg8vM85cwcNqver1PWEeY2c9LmOFsEqCaTPb10pECJJIgfJwS
vbErtQ7bfwzSOibW21A/+kXRPUXcnITH+ATd3GDptHAaL3ElwFmQzSH3epcuY7875HUV2MCA7W5H
WHW0qcFJO3SelAIq7nXNAqavZSO6oX0Jesz3nQUTBlJTYRu0FEaeKWgA+gn2KG/ZJCDlhk+969qQ
XLX/TnmpR+NfmZO69hjtafYBEW+BNfuKfRue7WOERoX6olo29y8+FPAkWDBNwMU+IlOjrlaixKmS
fDJPJbbD73tNe2wy+5JId+pJwRvjkotQcjARujWE2UMAmIEPGGG88QMhj6IOkNlWlR3Oq5ZdCJtg
GbxE+bGr2UfM4BW20Pg4pD2ed6YdyFRnvfwgUo8+FbxjSQ8E+EVGZT2UQOKdD1K50XiKj+2f3ouc
HwcAKu7O2yqG6k00aOF5JHcVyyN+TXm+/cLoo6F/5nmWS4UHrpXX7glMc9Vv7e71IfNgCSMlHNAR
QveOIJAjjrU7nFSz7gXo3qsz26oCfG1TQTliXixlM3cAC9Gt0R25+1ndV2ouHS/i+9Hr3CzzGd7e
eUFN/4NxbulRVetgYZvZm9NqBCbJuecA62tl7asMXEXoDmglneCOtjWw5xrizk3pGvlz0s3ISVSN
cw6ubwypH5SfagwBxCAJEt3IYR+90q9BzyWBr+kODsAacuPonA6IMFCFK10VQSslZoqIQmd0NIC+
3PupOone7UFkApLdYnI5/4ui7zY4uF1pAp91Q8jlJqrU7gginzbvR684koGLYsK7nl/ybsxrEKIe
mf2pLd0/5kzKNlUrb50G1pHXXYioAVV6Sql4PN5Q/i9teFG1H0Ic0N8rdXjFpyhozJPqaVUgfP1G
31zQng+/nqhTLpZa9nTyY2nW2rIiBOiOU8GTWoQDtae7Deee8HhENI/pnoKri52Tu3Aj3JcnCI6W
epvgMsbCOV4Q4SVHiSCbKrJNwQIJZFOaudhYwR352vLBG5Ph3daDyNrrZc8lwLv1eI1IBoy2kn5E
xcVju/TSZHA4C39xthsXrOf3l2mq/AzdyOirI2s0Tod2L6HcL7CRPj2ABbUanbnIymci2tYRWRZm
Hvja77qPgPq/IHbxocMiUJW6eMXYk7sxUm7zOOpjc2L0riL0wSv2wnPzbN+xFhvE56nI4xEgi4bC
7i0r3pNmh+PT3zFoESvdMWONkW/tw66QFsxk1ad4HcsCdQnae/AB/6TRVgyya9KIIP/V7XJ6d7Jn
Rrd6bpjbUbse5xHBFbg7PDKt/oGGJfjoW2RztmcQ/Z380VnBYTlcqh2g23s5EKOyGqAELJWMVn4F
CwZpfNI4J3/iQpV3vnVOpVpdgDAfnD9smpfserqgcNuh7uczkD+IUA0Y3MoMDn6RGCgX+5+e/XAF
zohT0uE2ydz43FTu5R1UBUGTrROPp4gK9rM2msCbJixIepKO1cwEFLTlHALLwSSESVIfcSCmfz5T
GA/7g2Cx+kaHHwDUaDzqk+yYt1NWixvMP7B45hHCSFvED3GKMDqFQMszfr8AcQC582mGj+ivSrgT
nS05cCjy/IfNia4Co9L71r7NGlZGlqqGzkCDYgDmqJQgWQK5jhBQrUr/DEuJ620RvBBX8m67uGfg
QXYrJ+yJ8CGDj8CShBx9MmW/4lfY2u4IGHn6u0g00z3LxqaduuOfioGj9oPTdmCL5rGutYhtrw+U
l/jaZRu+tCGhYjLLPruZJL4sK5yAbAJQ/cW3eB60QVO8G+rmkT/f/0291yAAY2B+1EZEnSzlyHlz
0BtuabWQl/BZOaOGQ7rdLsj5vkVmAprlBvxm1Zms/RsWTGUmVmkdB9L7cqbzbQwCP7X53aAUSOBV
abGTXZzQohGr+g+4ZZOkx0lykzaZUNfiNxDPq2B7vZwqVtoZQmUIb2ivApe2fbdkXbhmfX18u/o+
ANp/DNnG0N2Zh4HDbm6loHa0FwUdGQI424svcbaXRVK4U/GXCGZpsv+RoQnU1JgfNNnHO98RafyV
ZCYQBGsNIPLwzs7ojyObkvADVgW63ZaBFWfSrHS5/SN7hYhVWLq/dwxKIAqDNuKT7/RI3FRLfPsG
uJyEuXAmxDUXBsD0BcAtiqS1faeOQ2YqGFOIvjzueWWwQzLsHkY5ZL8Oj3pocwuPTKi1fHKRAmlP
Ayn7Ibf2JGbP6RTNa/ciueKkbVQQdxJ4I3mimniD/dvEQIdR+jJxMdXPw9409WxhsS9bgCmMBoeY
FyrvQvmL/I6uovSOW3dMHyQ+IgZnsi79UXsD8vQf6OQF6fqEok85IiS1oAE0Ww1g5ihppyZQCw98
K1EBkqIIba+7rTJ0ExGXjnBbCpQaU1MPkIZtucG5/r5eevzqO9difgYCul9bK/RDClI13ZmG8Sen
vcKw1ai37K93vrYIv7+e8eTHhvxIQrtv1tTkvXsBYq3DeF0C44zCFnPRp2QYT5XfVj3tLVJmbPjK
dbzBdqTUBZq+2GS2LxnE+gsAlrTeSsEtSlQdYBbcndz/cuz3XQtefUEQvaaIPqZhvpObGkLmjMgI
J5HL56h8aZ3LwZV6VIdCkfChfN/yEjjZDZ2Z6o7h0NJSoX1V49gDSC+c/8yuF+fOavoyheOGGGPv
QjR7NJHnF9qYrvWHTA9NyhJ9CsRZoplyqweXObA8judpEUxorpZerISMSmKUJPLvvlyXXttNMSPT
zO/9wt/CfpuWT89ylK35mU2ZtXL6IsklQ7uCJybAyCrgeKVtQIuEOE5zCSWOB0IDV5akS03wrxwq
GxdpxoThXX8kCzq8/7L3uqzhnAhdmbeLvklIhvy/Bt4PLhwY1c3UdNuXZbcw7HYQFEqxUYU9bw/V
qxRy8GbM97+v+WNq/9hTS5JijH5p8ibsWtB7CEfG6mTB8BUPXKVFfLNqBovEhpJfmvEbjS+kV9PI
O6i0KaOLyo7x7ijZXb6EnWHiaAxWNLyV9YpTbgbrNC4Ivydop6pQ1mk3ANCbNEZyLDl6YgJaC98p
PPLV2Edx1LOCGflUgoVhe+BHXp68ci48RTJRC4ETlBc8UD29j9ixUagTP6LzWwNCcHlXGWdJ3tL9
oaIbQkP3vxI0WAD2NTEfZsgRjphQpk4MVDyZq57mrurSc63/CNMjnWGxz0nv6yAKMdGF3nZNFmU1
Nbp3eETwBSCcV8Hlac60L5sZqAb9oIV5JbH7Xbb4WspqIf+FOyWOJR2CcIBp/Lm5u5O3RSHqtFdS
83KG9RKCXU1uvKsOCvdp/sI11yu7I845bDK+NCUj3ifJ8UzkhHxCx1x+JZ29ZBqI0sTJdUJCC5Oh
3FwUNf8/c6smKGS0E+N1HWovT4KYj9Rori/7NYbrE1OCIddkWtAAHV7iDYl8F0X+aBBHO802TESk
jXUpSrUmIVHt5wMi+lHoAfIMsosqjZhzOUxoBy+bOq+MAvF+7TVLlo2RWWcNRsRTGT2VYAIm/mUm
gVR35iSTRZpNXPuvH819YPJx/4W7P5hi2Cs+37TUYoOLvngIIjk1yZZQMmMceKsbVQ3+s5qG23nR
Qw5IlfyMgae+TmVLBE6iNOebs2t++A6adJOu55KJKPgWkhsQyi6kcwpbOUTyjwhR0ly9W/5hbrer
W4aeG8Hw4QghAzrqKjkiRq2QfnXpd2YdZBOjuiurELYPFif1e54+9lsFQTDe/g5fMqjzdOEE31F4
R29rTfIm9XnZtdW8BaXMJLHCMeHmoV6AhaPUD19VfzPtdTtfrpczCkcoWbNVHb1dI6r/v70S6Gqi
VclkUltJMsz4trKIedaFanUtK0kgoa4JV+rputtQZVMSHUcbreusRZJQQo1U/VtG4afPUACSrkxK
7/pcgISzeuaBf5m0Q6ZHegMVwyYsmFZrOfJf10t5EIuYmNSW56WqRQRq5pF+/t9yCYTHWYsklku0
f+ycFJVXL9RISSFOfjbP4ZhD9csWLA72pOOfZ30Xt/CohvHe9PcVEJGDLPjMNUTPEP8F5O4jcVlk
/OSEcv97wDYUK4y0BdXNU4R9rJeXiZeu4/QEnDgc+kODgg8FNUmB7q3U9gJ/TZKZ7TefDuK40GpX
ou8xyLpYrwBzb0f8yR47OBjZc9KgzMIBLO3nZD0fjwzPaqbkA9VyrHDi9lfmClBTvU5efE+zs8D0
3Xp+0VkD87L2Pu6EMtWIe9dU2dF/5IBvIjERPwRl7TZbSsmK0L0xtevi3er6XLgbKf08plBTKp5w
9Hro540LGGg2SeTkI8tB3DVVdm20lxTyUQAvzQ1HtJ774gian5SCkVi/XKCiU2rC4PmrpgKS2jUt
ZOV4wIqTEPG2lBz+jb+/nqzvaWTj/Gv3alpZgfxQy2uvxgMeZZn6+wDAVnwxRfvUmR9bvJz/72N0
al1dsysLs8zvowhz1Df79Zis5jUeI1eAPMfz7z8laRw6pcWKAMTzRHknnuG9kOgD1wyiQPhQrxvX
qth6inxIRBlXOz8v7smNoMx8huTQpU0vmqwlBKvi8GnXnI4ZKe73N6Wm1/kzll97/vgYscQSnqBr
hJUYaWRKRoR1htI4+JIVtgKuMD2js9zjFNfT15UYXfAd3N1Kc+xQ3vfYA0GgytbLbLSn94YhPsFA
Ju8EVMipnvlxIoGe9eVFjnGb7YrFWwx2nrgnAgWfeO1Hu12UburQ0+Qwq01GBIQKPO9GuDdhjCSl
3/TrShVqtF7IXgqfWr4wH+78GaPUqPPmbUimpztkcRs1ydXFMn79rY/52JApvZPQ3ZTK8gYvsDFi
R1h6DZc4Q/3HmaJjybeVIRV1cfSWg3F51uAPJQy2AjDGZxgWZR3pGedBPnshEVpX5UgsaAIz2Dlu
z0wHTT8FvvUk8oVrDGSCoX3tCPjZS76YV8amFcEfSSkB8ZINwoDvr5pWG8sAl8pVHRyvTHwTmf4w
1HbClYWTK7D7+F27VxnLWctN51LH37Pw8DgS5hUZKGj2AQZ8eHyQeF2u4SecW4jSwLE9luFvdL1s
zUt1E8EdQBeIizTb/fIMOej+hmoKSB51iffJr/zEeR1i6qpqw8zxPGnpwfpfFolMQywI50sbq3cp
z90ULVgFl/lbB2NyYrYp0go399h4J74CBAMCgDGTHY8gjM7eYFItcMBbvs1kHOiPZXaIBK8SUwNC
eKeb8zk6RLuXeJoXTMVMi87BjfR7HEkun0Tn6DTI15ORqOPWIsVTAMxBV6ZgWSogWz9PaWw++v5S
DZompUrsxEOO/J4O8A4y5N/qjzvL0wtlnbgm1b27xySsoU0dhcswuCg2swnAmsQQ9YVnJPnqD1Q+
IeEa1d8LFy1/WGbcIP+U+QfnZmnVttavB3vQTx66sD3PNbY/3of/gJA3Bff8GTbuCVsBqwB+fCJi
Z491+a8YSSW9xco4eFSwOxUKDmA7bL7Akl9gZFp4FnloOd1AFDCRPRDjVgX8H8y0ZSHsSnFTmK5U
1QoJtLFdDQ2aFVdIOk0UoEwxC9Qo3+f5qdbxb65q0VD/+kACz/ze3DPXWzeZXNFXEAHKW1dGk9fI
/iwREd1tjJtqGwMQEDb6LI4HMbh9t4+k+EC9mtob1u1eW80x5Wiuhqx/XCjmBj+aY48sD3e79i8n
ZUuBWuDBpJ59Vuo5+DbXfqG+YaSZFxhV+BFWte53rXYcgVSaHk7GSwf3YRTBO4G6aM9fRyTaU95k
B0dt12U8cUMafhHZ7WTqZSrIwub0sxpzu098ENssGSt2SwUxVamhfPK/XaHcPesoPDVCEyx1i4t8
wMMvpVV7MYXmv/FSmmwmRZER+cZg0n3EVh0yV2lC9p5MpiYPvgHB1/MVcYrSpTaqMW6u/IQi4V8t
pVS+mkHhveSvvP8f0llnexJdqJ4dDHbppHb18ag1an5jWG2xxDxny4p6szHnoRkcBQMbUwVFo4NQ
H2+Ra5Q4i4nPJFD/cJ0i6IqUPVjaINcO0X6wd7XMxPjyEO96pJ8orvuLkxR2Ru+5EkpbE+lsangv
+TwPPpLeV9j6qQc3dagYJKj9wD50FRZAbifsz/SeJpAGjPT04uUQL0hS8kDWjKj8TwPPU3vshi9S
riD62hyzNOsQluBB1PNjonpZlaRRUIVxSrPfe5D2QvBpWDLJLdT7bo0boxr7v+hwOIUlqIubwZE4
s3teO6w+4RJ3exvm4dSz7rt68tWGuYnWBqQJK9fWvyT0iPidnnudRkVq+8aAOAW/0tgWdM1+/C23
TPFVDY4xT4Sr53UQ5VfuZtYGZ/ISKXCkkuSScVDEuRwmV6MA8xSQ3HJcpqeDBZt/+ZJtI1x/B0lQ
ZnKDxO0MlkkRST8IyWHT5UKoCeBqdiIsXT6OZVtD6T4VOtZoH5K4d3GxGpqHmxW6tjPwJ7sbSGMT
l6D1R/2xu4X+ih1dk23908ctvKEZs/BDHPY0x1BEk1kGtI6L6WKVcQQbB3G6VqPD2c9rOiJdgFAj
BBRjZQM8///WXvLxSFpht6L4bF8TUxUocONk9J2GgOo+AL+VlwzhCXlpHq0eG1G0azVOAfJCc/U8
Mpzv4d0VNqcPJ83jx0EvFBvZ11Q0agJSpHVX1hylOBzSlGr+MuXz8XH7fjeM0eCssdOGxN4108f5
1diFM+NFwyZhVoZjhouLSAv2/flqBCZMJAQCm+FUTI58nOXJjMW02u4tG8H7pRiOoWfl3lmr5fqN
lLtnXejilb6BhxL9JojfDltiFyaD/ejut8j9vick3H7kSoswRa2W8wMMOU92Xigt8UsYaWacPd9E
M1ke0j/IXcZFu5rEqFfBy+yJH6dedvSKxAZgg/Mxpx3WL4miCVvHLmG+bdKqr23AOSv4kDJiEexw
cekTo39/waGPildizmqXhsdQnAZQkOGkhe4Ozxbimp/LW2i2kanFryYJcm3MSTMfEe9+Jbv/nFfu
ikX5GT9sTpNXqfhFt2MHzAgyTQk8S/anzW1VN20gWQm81kcPxC6jjKJxuHk+ytLbn3+V1U8rNHj3
9zs1uzFEN20W2A6anRx99BokEZhxpGfgM8Cs7iqcQwd1/pI3B4KszFfFhW++dLjbkoKlIDD7+6lv
1wI3mnuAQguZg/VE3yb29IK6wo+WUO56HMbcpYgu5RiuwPBshnA6CWO4STIldNQ2vc1HDrzohR/u
o1S9zbQorSQhaoK/uAn8MLyv+UIW0Np+SPGH9MuC+4O9A0Q2Mcew9xwrudX1S1I/e78nissEgxGU
DNpPcR98cP1SqfEODQBPZtPpCBZ57pAJhUdV4QkSkxK52PJn+mYLkcMW1tKFoMWHxj0e4pYrGT9a
guICHahoCRDMkeY+Rqx65pStfbqUrJro/FHGkJNh3WmCEXuWMwJrkjaeUA9F56Txb2pIlH/uYCIr
mZe4oUk8/I0NYkKnSjA1IXUQB3F4gFkzA3Eg9h9C5romJ4X+EVOtmmMlo7mdYycCRr7ijLYOKOGA
LputKLCkoSVua7CWsrGtMqbqPjzjffDsiaEAuWsQ+pBaHQYMVZDNUjqc12BG0sJmk9RL4F5VOFYf
XhIHzWS+0FGv2wWKMmkK//0FFT8kI5Ha7K3G5OYTRJtv1r/zHeX5QDdXNFcqQDkq7sXPC9yCUUBi
3csA8HIMIa0TXI6LGV5qxzpAxqb5GJDg1gbL2199iWz/E0wbIyamAg3QTQnnTn4oPIGSz6FTckNp
BWe16K42YsrJ1QYldnDio87gqtm+d83LPoe4FjCVbcoomZX65XdB+JFsnL7BpbK2b8J7B7caQYT2
yy7kstZntrs8QD4YOgu37z5sQAToC3wS6tPY7kaj3w2R6yqpyC4jsUV1g58O23+2l7/o9g7MWaA6
z4+7DgUe/z67sGSerhLYMeUiOS1lgUIJMtFBrCve1JoPky6omeo3Ci0oMlIufuAVm9a3roIRkqpl
QPGPH4cnjeDwawQnsNHsJn6gQBTQFl8BjuT+8ZDTade+mQcgo4pfJPmwT4i1KiTDheJHFQJv4NwX
0Z46AGTZzwa6rAc+WvnGIXAYu8c+9IIvFTVc4LZtWHAcIYtqa9xqX0fEYDQhCxtdHON2hyDqiJtW
xPfgKkerKkoGgMka1Ipa2ZgSaAgp1dvFpe50MHLp24mLZ/QQiBT5dvXmOccGHB2xdk7P9fz5Vh0M
hVmCIgbegYVktJJB+87/HV1+vh/xVWn3BS0Qrhre5TW3HIi6m/6DH1iTxn2mLCDW9HabHUFXEp9+
CeFWLle8RM0RgzqAL2S8gkznOxZVvyCBPbk0LJQI3idXmGtOo59P473eQPPJvX1kAhZtV8dt0Hjo
r9xaK8miJi13tcGFQPIWrmobs0V+uMI1hrvE7DwnaVBBOgVoQrN4t3z4amFVp7dOdDvK43fC6LqZ
lu0KtsqSxg6OGBA9FhmkhtbnKm5NQ+UexDn7g7cr/FsPMoYU5To9uKkJELOg1g5afRIuZPb83L5/
hH8zoRBhOkFcrjAj/bcfpFBH++wXDSTwP4Gy76z+6GzqB4j6mJbvaPEMOJpdc6vEhn+tad6hXs0d
nPHriVFwaeQr8xyVKmjOfRJaJpITcittfcuGRor/Ll4BJG/mVYDd9GTZSWewNVDUwwg6SyIKMB2d
NvPQIMc/T3MvyFEakoQISjotYxLIKPnNRh03I3MSCrDIFUxZ87UcOURvOkK5ipYH/4scSRZGZ8l/
WgNW+VDZkidYQy4xQ6FYidSBYeIz8etyCeEXbFPMXOx+gW42IX/h+SbQ01vTJEHTnFdZAGC7Qddh
4vOm0t5U2Me35vbTSBUVA7IdwBhbJ6u0v8GV5IMIYWBqwTKBoD+JBB1kam2+AMn/Iy2fdQhRZrNd
T3J3Gv5XFLNfURm3U5LTydZ2hIh1Jf5UsQ2WfCjuAXjmg1QPZ/xxix5prHAhXpsEWUoN7U4VVQF6
zVBsjvLvOB7KENXVJC+pPRiBdG3K4yQZZW8zYUS3kp996oMq/VZ02GQgUBq+O3+vJvMEc8tCPeKB
/JpvT20kA36JUieErc2+QoWAIwiEUjSUpgP4443JwGY3LFzbyo0HHFqjP0u7KYcPCRJXnzDntbKp
WMwCkeg7n2fEbGoKAcWBh4VhqFhKEXp3UIoxvubmY+jUQ2pKoMjgTlTKCW7FbD49tBMihLlSEnz5
bbYEbXS1g9bL9SPOtQnJvgDp4GmLy6aq3Z3kYo9h0Pu5RekPTNKgjjUGpI4zfAuO3JyF3uuikweF
c0YnIrbEhNCmgqHrGKR2UM2G7baVoCMFTR2lqDJcuXQcKam4ob+0mcBWZ99REip0aBCk61PeRVzs
Ev+KCSsRDBb06N/TdStsGSoIdywE7/6JtzHGH5hKBsL8QYjipRjrcpXpHo+4uJrpqbZQxa5DlLHE
eGlTX/Z6Run572NYs8rqS3oII7sMvEnURjeOwaiBBDfKGXzIRuNmR8eWxMPrcmizqETjnmVmLtZv
7JmyDEYaDqJ9Rj1TK4M1AESHMRZ+AioJKK2jDOl4K5KEsALyqChI7ESMBNdcLpXF6A6pcdYSdXyt
CoYpuUPRkm9yps38zCRSIfaI2e76A/A95ZXC1Kbaxbgkkem8gjak+FBEaKxvxdUj5sbBO7b859Or
y9AuEbxtKXaTAmBgvnlRW2ad6/RX54lHALxUvcXf8iqJUtWyQkE0FvxvbRsfo/wqXZbHfj4Vk1tO
5twU5FoYSzsMJIhDfRIH5OhcgR4uiDIdtfySPbneNGxacBJGpD6dYEg7cSo/spHsZZTvM3DPZTtB
8O/q27HDlAZRRxPozuaFlMvOjRkt25Efozbw9XYecBi6TLYX+innuvEeGx6hmi8JP+OzmCthQGnP
hoZSUCmxo6sq2BHcgFkBtq1N+c6aKQ2zovAOT5+anQr7iS+mRU32roaot5J1l2zaX8YKEoCxSkvh
1i54JzBGl0N2Rln4ozqn4r0Ax2cp7e9bl3vHpCtAFE6idGuWFAMRDBd++ribcAZyBdANXPZHNDkb
ni+vvrLeSLbH8wSdsyhWwt8wtDjbjA9UaJE6KRwzv5O4CU51HoSZpNhgYLtGuGEkfQJ2VVp7dcW5
m5xbgA7WaoSLsnda+EdmS28hH0YRdGDlenPvAyi/4nr7NA7vs/bA5zCdPfQu+9GqmGm1HHePOqN3
VdFGOMt4HYmH9nOYlle9zg2sC8Jl8FWQxaiWAlazX3utIz27RTCb5QD9g1KVOs5nYWOraISAehgn
ngJqtOdRvYi3fRgZNyzjMnFjBYLpPDuC0h8nZ7hX7BAE1WlKL6qUlwWVyhsrvGcrE3VxT1cTiDB4
I0+Dt0o+ppY7lN/vgOeCWlbzQpqoecTmhgu8qxgRTGAkI7y5VTtexmvJqxn6OATMnWrdTW7z9fMf
P01FmcP0xo94vAeWfkH3JnL0HPalB0MpTnyLxuf9P1Z9rph15rz7ctXhXQj0d7gK2GhqUgO5jcVC
UhL4iTELsdW7LpjOpDps43It+keCOOeyO7oIUXrnvkIv1STlAW4ru544x5RDOvqNto+PmhpiziUn
pyJpgIvOAfHn3C+8EBPDM+N8ecnUJrFCNiT+6WJEsmfbTfdCskXpFpNEw40jx3cahudpoRRuEGdq
doELCX5BEFowz7MbD0CcdN+GiYbgs15kWxHwp+kc0H9WwjuIaQfbaG+i1WbNL6Nnt81jd7/wmFx+
9SXuYZrztoU8zyA0kaCC6igxayeitFumft4n/Kj82t1j4CUdwe5WQKIftL5PXXFm0BfzLx+CV8Nw
mr5vPwB9ATt9pViMrkVLrIiRoOxz70R7T4E3qQ3Qk6+9Mf5KoisiQhaiu/TeubhOe2wQI1bWPvvU
51ik5YTEmNvPhY19zBpWq90d0vK+mlDgLCyIJ9bCBb+TMVo59/gbwpf5s18lR2LZ6I3ngQDwlkUm
qZUg/pZUg6yziT1IJD1Jyg0lDtJbaiCfhB4113N8v45yr5GtAJj0HZQNRW4kYWL7li6grdJolzHh
V1fQoMbN+D5IYV3jIfxxGk7j+LGVeBHXNVg2nBhxRyPH89nGZIn7x3smYtxkHfa8trTnOOqXUUsz
OfrNx2mQ3aJ0Ha/4B3tMtyrZI/umVpKsMbFOfqFq9lKchiZ2L4lwVQPMkFpiP3oAYAJg1KsSQXZs
ZbJomw3pFRnWREri9IBI2B3bGH1BANE+KawYUWrEtDfQRzK6dYTK3Yd8/8NRasf5OlLZVKpkncyh
H00PMv7lCXRHP53N5xWUsJWCNpv5I8j7xOkiILJimpzqR7ssLZfZSvnHy/sc8h4D4Xg4uOb/GEl8
tiOBDTKgFZdul+2sUf1KjMqdYaV17uEjvvmNPkEVDvMgDIb0M3Z8prKPtK6/XRbqZOFdAJRpaBaa
Fwl1yKqe8Eg5RjBSSS4u5zRHdNsQBQn/UVf+R8bTQKXi4d77qyYi9p3uJfGcQkeg0+1r5ydlQImv
CIz4VLxvRT8RXShEZ3KsMjEyvZh+k3dGciVqwqGFj650OGhZS2z5SNSYafXGaIPOAF2nXoRNO5zC
ljhdpEpKXxJkbt0DeRMBVytFdGesSpDNUgc3D2IHvwDPXdUXQTfKLCtF3wA8umUCJToMZCv/XUBK
eI/IrijIfE6s0SBKGV9i5pmM28fWBbHCXlfswQkqi3+Flav4wsVO90V84APhWoMVtNDNiuEp30gc
FWrKerpSfxEQrfVTNRuP0bIgI5twgnjq0TcVz6sosgj7ooPeaBfBxMgU/MWvhHpZuPmcTjoCQme1
m0C51ksNxH8KLth5VUB7zML8c1TWnnYZyKOpBDG5N3MoVLvLze5DD9kAogso1kEjMOBp2mfA8udP
kiECLgN5p9PLFehmFUjwpSOqVnJEwMMm83yt9014o7GFWRull8mb7XuSsg/OVYzJ9kXwm4ZMh5En
RT2F+8pKLciqgonv0QuC1JrhVwXh6XyT4maOTXLjwRSAVevZcRfzW28WnOqihpxvPxtA2HgirnjX
m/ha/NJ9RRDAJsCyROTyW5JCSQpdYiUQfK6QOiOXa+pAfVhuVkDThXWprDU+6ZdO2utrMkhJcd1E
yd6gjqYmp5J9c8A/fo5f/E5U8SHrxhUeFwFSdn6tCNF9ftcUSCQTTjSqiBjz7z/5c3hMHfnPTMWD
hKoJHsHnzxscdLC/GuERDyzxymrC/gzEcQ6H4sLxg+wnkv6blz3MoZe7GPc41ErbHEJQCIm9eMVq
bmaBzSkzSRZcKzvotPjw3zV/X1Z3S2dTbGfOJE93XWNUgsU8aGnXdX3KGi4/tlnhQ2wMnR9WCcmT
esS+Zkvcw04/x8lRLV1Yqb32/+e4btmYXfnJGPbIRx9wIrFKNB82bKGfw6DMqR7GyG1pCB/oi1Or
adFfDqZK2XuhUyy0kmTiXPETWufQ8dMPSGWgVB3NPm3sdD9ounPU78NQh3NhOB0C+31kuhFeLcz+
9kL15HLMATq74rfo0dpe9C6ks9xwGlG0mPgHRIUGEmhbmUcIfDRESyWR/sfrc99CgYxp9hr+ECdv
cKyAcGiEL2qwV7ObGV5ihDUgzaYa6HzAKQPd29E5ofM043BuoDwbRFpDDMJoGLDbOsNOoI+6+ISX
KqVF0L/9o3ivP0TQGlphvu50Bz8njgahseP1g+SyFTzPMjljg0wO5Io1SFtMJEVuMOrGnlTK+YS3
XTZnhhphLMEGzGDiHcXFc52cDXDjDVsjfHVCwKPiBz1ZEp+yDgUMQM21Q5M6Y1PS5yY8ydzpFBER
p4Nv/xZDQiad8s2G5Um84Iyu6Eg/sxADgHnU/k41Kelqv4WZL6HxZg3xLaL5rwWhRNpYs0FNHWhG
HbCsxGuUTFTqONCg6aenW9577P7f+x9qCZN/lXNv1DiZgsSWR+QioXhU79v8MMWBWBZAC/Iag8u+
oOnjmcQxSJtBuOMVnVEcmb3VZhrCRozGrZqH7f3jV0+EzDnRS8MlYMwJb2Fr8Khcg1Uf/JXrqyPq
4jhUrM3B2ACrK4qMmxHcjGbm+TMiZaHoRvVsk+TzrdiGIgJyxlTCgccX4jybCDWQxa4gumsY3xbd
xCaPF6bZLDUFEnx3W9agEbf79camrRWPn038yd3wDfjC4qrpWJcBmgQxUcyqvj0OquxSG6DubCAw
L/YjT1E6Hw4e1InEud45QMgepAZ8dzi0zJBoVt/zWmslpKbtlGapP6aXxFMyOpIW5xylnH6FZFuy
aTzUxeqMTnDLSNbCFN4c2nu9ftwrpxTh/ENsj+S7JMdxY6chm2d+vJuW1X6kmQmS4LgO+3eBH2ja
8ZyIbRJaNKcflPkL1jkpt+/w574tvQ1G9n1n3BzZjrymw10hSwaALtL+QOgw5jiAupkmxdkWfsGD
cg5Lr5jQ+U1/LObPfSVN21mI7SwZhhGkZLFYkz9/epx78JDPLWD+7bF+XC9L7y3pRDfuPwcT+24r
AFZSoggRuagmVTsbr6tt2qGhlZcEXS7ObD+gqTIIsLGhauhFCdeWaQtN4ZemXftTKxgBurtBGs/J
bIsHeqiSSTfy4UXGd/itrXKqHGoYrXsVbzhLHNV9xeBoNkwU3F8rX12v5XMdV9j+U5AVPixqZYJm
16VS7j/VrzwSYF1UAsP5B+HNsLkWiPKt5CIu2WMOF5AaajItIjUtqLm3sUfEg7npGNv1GLQybmyp
g8ruuuZF2s5qPLoAonYzCKTA3OSv403gDkDEtLzkB33FZTrcFirQtyaY7+N+SsCPADvCuIm9Dwqf
Mod7o1stRWvyk0OmDKLqbWluIwPEbLgAV5snw7tKEiQ2pSNN4OqKGWvjTBWrySgbJToiSu3g6ahJ
40bMl1J5UsSM2LQlfW5eO3HzvNi+xx6FeKRa8ax7JyaJj1ogTwS8MqBcUiW/j0eqM4wUhjBEvlRR
IMxi3vcEg/geQRqFZhz6rJ+Cx/pJ35ChwUBaPtbXy6t7Emk+CchQqx0ft0EsK+XDyljvVgScEJqd
wHzzKX9DD8/0t94BcGJ+rddryvZy1J1UjEVrx6s/+uvloABnQ0B3SiZhdEYr9KJpfDGbvm1Qv3F7
KWFvVik2BCLcDrRt9VYQ6khRnlj0o0eaJVJTDYCIFX98hJtdvk7X5mHzZNSCHaMcZ1to8kOYmtia
pA+lB/aWFbJtM2rrdJAT0OgfFvjvXz3bVa9hfI5K09wjGJPerOUtOSoG6QbRIyq/a+CEgjUVjhQI
3+tskm2pgdIB6F8Aqu9bUvzHBTHYct54+GHojWXT+JgxGk6DSS433UBEKWs+K2NLAJaiE/oiujBd
lIH//Lr1gAgcKHAEbLraIbuJNluJBrYU1o/qVqflXe2ltMFpuozFZldvhqA7VnXBRUbpMpuaAwmm
n53ssxvZdVP3t0QH7rZkTBDsWsBQmM8MvnVzCUX25rl691NeNaVg2/StqFnn5orjOHxonJPzGtCe
4F8ZOra/f56LvwagQwSbKXuabluBCc9+U83IDejfmTrjp3KM6DIUPOnUgM+znltQB/3NTEajjHbL
c+V+jpmQQ9Z2QjP97FXclJar89RIP5Opk+PSSaILYa/0hdeREfTOe4hXhTOVwkrQJgqbaXYBcrH2
fXjpI/WlctcdsXUa9LKzcGZYRS44wZg7NcbAQGvbmhSn2DIQjlUfwcOOLN2v7FF132KVmo9do22j
jmSskRlvJlTu6eTZDGpwldH/U3JFqiuRMhZ+YPb5TPxIuiTxFusJbipkfe6mwoFzM6TWB7RDM8HE
snV7E4f0aIdrrN/zdZcAq8POrg8e9oMDKEnTJEG1qUl/LTyz0FKsmswdYBofBOC1mOxSIkENpJtt
zw5atLlG7vKHGEYX1FExbs+o2Djh8LKXPbVs6zWPCRpWgErdCZfgmJNd3zNjLlHGO1dJ5NQYy/mT
XfscdmUMsB4m3Fnc62GNkVkbs3BxtJmWwLR4h7cY6m92gN2v+5wjrfp/SdLbpLk6tY51hcC6rb0Q
znR0GuhyKXdE+D/C8Avc2r3XqAqb8kF5HeKM0HVFIsc/TWW5qaUBBZi8d0hKS3FSJZywqWVds4zR
FLjf6Q1B0GTJ0e+BlWFer+CySGSW8OZf/qr+zolM9zj5QRzVFZj05pqNKGUfA6hGvWpNgGoDu0PN
OyVYe5TNBQgVRm7hlb7SZTAhx1KA/gBjHBwKtNnhP9dq7L6X+pRSsz7euMXFP7WKtXdZJ5ArlRmW
AKFI02PnSHtCQ5r8chkznRUFjej+Scz7c39NG9PnkIoUBcrBpWjnD9WiGlmJ6U8jnNA9/2sRDDtS
pAEdYyrAPpz5AwZ10JWmvVsjlJB+Z9MR0R5/Sr2FCRusFhX1L7QN4GYUk7R5ZCxvmWfXLpVnPPEX
6ijhEctHf68V8Ivr1iLIU9t3PEc2lq4Y0OsmXSvVcBG2Y2CQFL+p4VLPSdpFJwJTd9sHmt2GmKaT
ZlnBwWEfF4GNvP1Zxl44y+zOsAvIHp1HKZ4XJnl7w4hK+t7SjhFhdIqPfJf/kPOBHYY9vrrCXyWw
N0vFaS0s4kxLe+vn0maJ6E6uERdxmO9B4eHdXpa1NtxkGLUuiAF6NoT2FvG772j7GvbqFoeidUyJ
rrwzO+fBvzyXxoPbjXSyqoVue24SV13CW1b5U05yZ+vsLrztQZyDGzGSuPvJ+w9QCfg1uw5K0b6J
fInmVWtq0oAbrhkrXCWR7YIjha6W7jjH+TUX/6XW/uRtCIy5OQbl+ft8oF2gwPk2fW64xNF6wC8A
qKUULoBr5kTawT0vkt+Mn5S6Wh7LnHZor2WjoOIxKs7+jCHqV1dDQdli4vpsrkU8OfHVVbAhEn09
IFyvfrr964OnyXBg/esTMLmG8bCtFzjlOCFE/2ZyMBGgvEevh+qrHuHRUdruAogmjdbG299O2THB
9bulFp3lK4BfaJ9ffpgXSSSCkenLZplcVuuDUxAmmBSb6uQ1f177h8xCkh1rFs9FMoCrwLbZKWPv
9zOAoNGg191wx1+FcjG8L0n6jLon77FQLABxRKFUT888yD+3EO2g9dK7zXUF843uAPz23sPIhjga
3k23ajI3LUIaZ/H4WQlXnfzFJlaY3NPsqKrgBtLMPPQ6sZ0wOGlcQ9MNJALlkQt1q322q9WjMdys
UQ7Gurf4sg8rL/UnGiWPRX9A/feX7NBYsWEHtaBb+WJJ688zLtQZbQdmnQq/2m7GgsR4TIXuAIax
t67ZuLQmjRKLAKR99nvMsG7qmtsTzu2niI7Jvlvo9Kyc51t5G9id8ru1TVRX6+xXNbMZBTEEYAUU
QWEceFRLDcIcUuyoLV8IPaqv50mMFXe0/77h3Hs9himbwQebdu7Sip6vcCVDZn+PogJIZP05eGX1
sA+hvF+6HQsXzzFLg6oeqdZGHEmPceVCxGpaHV2+ylffqlwSaFYxdf65u2xeoCUEPxhyqAujbnqV
V+sFyj4fE33IitV6Q5/SGvHFXqUi2QTwreWtNmEc/OLzsKgNqx1YbAl8Z0gEfkac6+zQxhj0tKao
LZPlZb0iRZE4LBIyh5Ox0eY5uS69TSteyQLsn9hrEu8HdCKmCkqrnA65nL2sWxQq2xNGKHKHn0fV
Krqsm1Sk+3DkRtWEFRS8cYBQpcOqkxTMfsCz7XHGGhxvmJiuwUcsEOJCYm0g9VxndQnfrfYVjM4v
y+dYb6bvvWZo3PbZZ/KLnGVoaNoWeqWrqb+hPgF1T2lcKvVpXchxTI85VKmKVRhJsqqt2LgSa9ob
ZvDDVagHtwQpHmBhBIt57c1ZUk7aAB58LPPPteMMFfn7ZJgXkSvWOpI3g5EZPaJqK9880FzgtlVR
dOW38hCxsgX2NgtJmaBzkUTuoOo6pT9C0lclrUzQMj7v6YsmJnxx4BTl9sGTgqMKRMQyIOl8SiKv
Lyi0xVYh/MjWKurWkncaB638yDkbwRyqsadOpKHWCGDKJ5nbsmHB/ar3rFoJe8Kx0Kv8gBsj0jUK
fQuSFpiF+qd3AFUqmZtO3T3+pnlyhs2Ci3lGh+RCYBzbFC8H7iguLA6pTrq2C6NPFPLVgbeheJJo
vPuSlexMylxVB7m6V5hWHX89/QDRjOjpnQD3yxIB/Wk0oYH4zESmKSHq1GWqKtTpNl4CbrVy09WY
600GE1SzT5Z+jXVYURJ/ejskzTRbEtGz3fyCDYQYESjqYbXYeKeJsDcpl7dPs8T6atgHawG/83TK
zsb2iZhFy0qn1oyzN4dgJfp+yHxL8IV9A6G2onqJNwjmvNFViDmQcPcewZLHKFGXHeEYArczpKtl
QHGgmZFD+jAtBW7GoBVAZFanVJMr3gII4HwE8bDqrEziOZsg75sC3LLpW4/DrU0KaNFhBoO8/EZZ
kuctgNnQMVbeBX4RPajnraGeAKRoy16aK16f/GY40iJF5zGrQkFPSmZnPTpPcQDe1EDJ/OJoUd1l
od2wmUMnHf+ksiUYP8W4IsBZZr+WddzD0a8p82zblUaolaZAbXqawSQBwjnOEoBCqmXuraCQeKsG
pxNsI9vHeDHoftLLCA0ezm1TD2g1XeOXEmF9gVsA/bl2HKYJYh3GcoM1RiqbCoDmO1Dt9pa+sbGd
vCJD77iHju9NMHbuuoLkDHSVkZrjj2dGfrbaWgsth4/8fxlg0ppuFiItVFCW5ntHPdDa6VwFywhY
zF/aNby8C8ZZ6QH/eKKJuwXWMKVkr1UttxLG9bQo3m70vmp8l/X5ljD+7cz0sa981yKT1bnoOgEj
/c7wmj1oN7UZAZ+XE2t11FL3f8e/9sdrICxPdWeurJCIr1qnqqytbxGhGrP8FiFZJ1cJ/zvWPU2O
GWWn2Vm+2L6aZbOcEHhRPXDnBQ52xAWS8dC4hUehoBhKXh4DWn2ELxxFpDwCmXjDeKd8rglGZHtw
9V8PpqWksi0aLOfAGL7fCBTTWij1YGYUndSoKxmmjnOy4Xa4pXga2M/CaoNI0s0Dlp8SnJDhaWT1
VEa6Vg5ao+qN7a2c/meUN2gC0zdQD1rhWqHUN+lAfRCET6B2+Sq2iD7yXWqxoNP1bskAg6WQbPUR
Q1YOcCfzGe2pALxM9AdE5MHDkc7+CIKt8j4rBRG33pZBS0veuFfumSZw74/z09iVLX2HKmq9/z6Y
aVvTecji6Quo2KRvHwfwVkB8h/GcAPSV4PP/lNXBo4TLcuR/2epODnQTJwtCY6igGK3bLVtkTYFa
2kHnZBtZWGFywjMrql1brO97FmHdFGBaO/keQMX+oHN6tIxW/z3vEHwshXvrMvuFUc9OtqlgKyAy
A9ANfkFN5vJFLzenHU8zzsc91qF6jvhwsoN5QFsd0EzF+3JrCa8uck0WNAyPw5H7X8srGLMkDxFP
bOleZB43k5nrI6xjKH4IdU41DfjljNkBtI1F5N/YyWuizi02aRoym0brMy5qOGVhwJBrFKwz1OKp
X42xPVqI8LnYnhjTUqf0FhxVtUTM1cZVNWp7v8uRI5azycGGzoopoob+hmI7uEKBxf7R2JIwKmdf
qT3Xw8wb+nNFWAzDVee3eR5xcpTbprJ8AYDPy6tRNS3fU5A9J9W0f5G/QHqjC7PxY5+OludDCpmx
9PWUB3ckHoHXeQvF3uZmS3BMZ8pQj8OlYUShHtAyQ7vOvVojZ2Pi7vw0fhsDfx3u4J9SUohRvSA2
LCBGmyUKOUwqKGSEl9V3wJxEDzUxvS8XPFKkzw1NiOO3XLffFRExP20R9MV9g8nIAQGqH1renAlS
jL6KLLTzE8AKQ+TQw0cHkIJMw/2Ruo9ymvB08fYQHPxMWjcd0qD/bWPvFvMPvAiJ6sAT5VYVkOtH
lFk00tM5M8ujpRgnYgRNa3l1USXxSYFwMKosJKHVRvcAtcl7mTknABxlTt+nZFc97WQN7Is4U0P2
XtS/Mc6b2tp7U0xaafEXGuX5e5TwR23LAJaWhYnIB98QaCfo2aMULzTgjbhMVKjg4Os2yR/7gv+w
Cy9pPltr3CoU/hAl47gXTkE959TyTdLri5enjqQH96MvNo/+KHaKnEXR45fXQpcMqv86AcFlrsC5
Dw5poByFplBnEc2LU01fSk9q5YTLgwac60ytH8oX3b9krhngSyh9Fq8mh4wdrIK2obYUUTTDCXeG
1IMGuS9Xgu6xWSf9jbUFDgpnhegismpL0emn7X3ohu4cCDc5am3PzykQyzxvEOilx7ylok506Yj8
oOqufrb5TugEpaBvphNs2ElpoyIdGSP55DljTIXIQ703CQcAfCrxwwm7HuHXpRr2S+jx6YFDqbV4
+7qoYxsrdrsKsfHbQvNZvYDvkh8ZjaK+KHksXKnFSFM5EzkOx3FoigV8eYyB93zxSaFAlv2+4gdI
MloOSGl8npxs8HHZ0R5CjI/qoje40hfnNzA4EH8iVAE49aaTqJ1UWcVBluejJWd10m/dui3lHkYF
LzMdgmrZf9Hc0oMsTb0Ufyd2Epc07eO4hLAHe7eJrTjgzX1PM2aPOp7Y055HPAodI2MW25yly5tK
+GLiPlj3S6fRqi3/J7nh2ZHYdTBiAkgf3kgVnvageKyVcgmJ8KHuXPaJSCwzqzaVPg8jborXQIw5
GnZyFP5A0/pRGcBup/RlETreLRjwob8UM5q0ru3rJHZnDFQDqIhctIhGx7AaN6mFL0Q6olboG4hb
TW0n3uMVWkp1RWLkDQWNh8OkD/PNSjWcF7PrdEIJD4BMGYhiRstwaaqAhJExXr4YedJape9fmPf8
jsWMAG7L53vHh+XcEroOXxWHb0bwvAcZLFxGJDFPkxCJ77M4GcRsFEcJBmvLrRI9F37DmTZpq5QJ
4WPU5TEuxbpsNP2ldk71NIDluqgwgyf04s7gKLDcnmzL/djPdfCbrdYd7RdCasGXFjc0fPRhYTWF
mGJrsVhbclWcjuIQB7Cn/9S35I7rvDDl/OfdZjgAvzqw0k+mKQwkVyoy3MMHwbIVa20R1+qtLvTM
lm6W+fyGV8HG2AFV3ZDGrm/9NK862oUgmom2w2RPwo6/tLa0Ctcf/VhZHbt+HTkm7HLcXMv93UlG
bVLv1juTmEiyZag9c6W6LxOCMmr7mEwLdsnObm2+cS15gqG1SgPQqyimvTCGCZwruANq+qYDGjPT
dWMr0vKJnnncfi5V47k3eSvTHcvxxXeMZkTpkSSaM3ziPzzcrbl63QhWxbzfT51eRIX4qDW/WsZr
cM9Iz3z7HYShaLTPBOD6o9dSdIUoP4mdD6p6O5FbU3o2f5dPdRzupDsGiK+VxGoqAK6yFmUD2vDE
lz/YiTnB7i+jf0X6UVn/9K1Z7gYphUgV6cTgYtd6Ju+ioPIYcM/Jkw6wDGA7jaI7cAKtj1pp30Na
0ItHLqo2FeXSGbSeTKFYlF6W6RgU+SIf1FYPk782qrCJbJRn9NkvHvQNt6ob3lS7rr3BWwG252rr
kmJW3jAzBBHBIA7M6u2KQRmBQFmaKBtqA0Ii7S8WMiUbNxPhbAOSozoT5h1DBg6mfntPfEe8myEp
28VykJYsYRJ4D1Z2bjN+06mXL406sea4HAG3Lyico0wuwNboY/7Ml5Utbl6oII7rp6IkHc+48XJh
lZQh9g621AByJo3Ws5oY4+UeIRqoYYrJ5l84rJ07+FBzW9IzEWX69AgNm/VbVMbBkdSqge6y92zo
8nlYgTqumpeCpTPxFw2GmRwa8p7cULidZV3RsGF31wEbeDwrwVhfdfV4aeVCmboDLUSVlGpBwoRz
Pbp1JyUIhObVK9G0e7JFT5FBBgjXxWtwHV79qZ8eUBRd8eNB2BuzzqIhai6PKU0t7TNBMPy0rmsg
252U+KxM10LSpOzKwAt2IZMPWxy87XGuvM+3XmfliNZZWDvGRGcDGK8Hp16yi2Tw9OlZYN+PGQqY
PWxg5/UUtoWof3qaHUh4w6sJQVxsoSnnw4zZm8lBHMxgkEL1ra7A+drtneuItYu3asGTRVl0lwhd
+A93zjsqKWoSdyO97d7F9LNUzWQ1keW333MUuJkeJVUTaULfQ3Yxd/hhYuthozMtcNp2in+OpdPg
FpViht5VruxYTHoFYOollmyxqZI3wMa37Yak7xn04s87tUq3T0wPjncn5h9IB92D31Ul3K/L/Emt
6iMAKSuCRmJBuCoXEwGMkVihOdk5IHiAqWgQ2X4me8M5ZI6Ggvo8QllQ64IT4weqUlC9emT4cRhS
AOerEBpxJCz34ZfJOzT+koQsfRBirjZecQXJXgO1tua+aoHWMCCnNMPkIENyxO1c8mW9MMSNvUA0
uqwNAjunQvvAUeNePCXLMxm2C/oGaj67mKL2QWXlW+vZyMRWaCQDmkjI87PZcz6sJmAgUB+FHy7y
hdLsfzaCoi9GZIWm4BDMGqIhmkPlXHCJBN5UZLFxFRe/5a9Ytld0sD/3ylEi56HWzCF3zEIyKoVW
hFTqjoCuupCauM014aBDon4gMsgcnj7kMBHAJC2XM5+6v1D8mHbqe+9FZ4CPstaN/eliRJbr93yj
+znlo+xLv8T1hO7cUnJyr1HNnD1i79HsVuAFl4iEu/aRvbVG/fEYMepLdZEfIkfnFiIEM74oMtQN
VN/rJ8nWxoRwiatxhuj3psiyPspttybo/WOeD2D7pthA1euZwF0LZTtkVIcciFYtTxjxMWBdgiGJ
ITaJYhdnR55B+VGISMJQiDXXvKfBfYc8FVmjBgWag/H2L4O1b05DkKUSWfRk0oI2mfXmOozzS+Hy
unn5AKLfZlxTjCjN3zB1CHra1wjdug1Pu+cYRKvyFUEl4f4FLL3/M3iTRSq69/Uw7fw8Ys/kKwnC
wlh8OSDeNzMyU8LnIK3uZUSXVh1jNaayMSY+feFR1KaJN5hyyXi6FnoStgcJD/iXVayKAzYY7iwe
pj8re/yAdNsrQaS7/eVo+/FcA6mfnHGX5oV8CJ6crpz57N1Bbe9oQ/6FdlK3AxlvRJTWoM3cI82m
LxXQE4d2YXKhey1MmINMoHGpM4jQxA9JVTN7mSMaMunC3hf44QfUbut0jxjc+X71bszMkpglWvXi
XQZifIgKBvplZ250TGM0Ox9+qaFRA2/6k6lHvCh+9XIE6hfDapjODgCvSf1yPcR+5MYfVDh51t5s
7dUb0w93wtSP2KkSpSQnuuNsx3nrfwxCAuWqwaJOmqemc/DpIHVnYGjHxM4xlfRib5wrfucFKclp
d+ZScxLChLO0rAgQlXwBxJ1nUH2iJoN6t+z+C5q77iBr8Tpsi+muRmWUoIYHVQx7uIvk8Oo+iZ/K
bcAd4XpQBGx315S9tpQjaTMm1qLOPNKQHpWM2pu/xt1KeWvbTtW5GPRazlvhHB7qXMFXLBaB6E4G
SCQwb39q+dIOj9UtPZ2NbzsO9qSfwUJ/udQgaJbdY4T6lMHowCqTFh3aD9jy8O4Sp20o501Lm+ws
rAUNdrtuyLv01uyMOdhYc0sUtZaf5l5kJgouXRUoxxw+/dwAJ/zVoK1lbMA5ZCkeaDT2rJJqIc2U
zaDZckcVTnGZGbdxAq6N8YtOhThRJfSwnTEpe7QcNkQ4bHQOrUKq2tFTAPkfxH1uHAknzwkfBI9P
GMTO0HmOzLdR8f/yJohSWiIx+hNxqbeGC03OfwPoYcOZZhPyl2psfhcooMHdA97BQJuwpw5pPl85
BMiUPbwjYFNrtY/sE2uAGrfE+tGrbumYfk3YdnYOw0LWdMhqUTIvpW0Q05yMSA1+6+xc9g8GQ3D8
yl4z4QzIUdR2h0nGcM6OLek8kVHI6SYN1PLZq8g3Bku//XsxnZHqofrTdrZcigigvKhH/nYI7ToI
aAWrkI0j2hZQ47+LxObg3Y9Gw0d9LFCvh3wrzIYeJ06G+KET23X7TqyDQnEZ+6eLnEciPUpGOaOk
TT+tBvNYwI3Cs2+Lo8j1Rd9r6buggcqgJUHZWk1KDF/Q9HXL4T4c+xekHlJ39YIi7ZqfHC0yo64z
ebNLtv0CsKl3sHKrZG0xYFGA0Lb8ocHVPHAW6f1DRbSWVAv4ummqD74cDuBjUSWpZzSP/RohxQbc
nmI98bpSam3KHbcUYvXtpurrFDaIJhuf258+oy1iZNZoaBANjSGPeo5YQ4eCzvgasTWz/GfcqAGm
l1RgJITUPQo5+6xCuw6UhpB1J36Nacg5w4lEV8Sqek0mv93eBqxwFy3CEDN1ZJZD6ze7xy/zvY2Y
GrXs5O+GAMWwI2GDiSB9heZtlM/xjhId/YMlwKkWUl+lc2UNCt2qM+AQr1WWt37k6zo1u/KvSfiz
xWg+OZFiXVOCEmR0KRY+/iX+7nryqyFk1F9wpRf47pN/zodPZ8VSCralA8J1EpEUBCxfNCW8PZ3C
Qmb/w31ZYowDgmgZmx8BQ5JhTB0fwETbyNfcAPVgHQzjzscOR9qKRpHwKh4ZEZ3w9V+mCiAD0HJA
YwtSRm5goUXGIUy4eX5J+4N1ST9j4nkSJ4JC1rc3dwqfLVP4zl2N9llxR5ytUiMRDHCKs+QXOLYD
/iqlKe48UamFSHNkqujdxQf1AErId7SfgtuG1dlycEm19zba6YTEoMHFy0r0X3Q/pffUZQ6TUFZ4
zSp5HjB+jndMDzoqUrTnatw4UaCtCkuUxT7HrkjpPwHYXDlY9n403uZj/KS9a+oMcHRtGLZQ03cY
6TdaV4lTR9Ypm98EYFdwZpOT1dE+1+IGJqtuHIv057tr43e6PHrgn3Qd6l61zaDL8fhzUHlwbIfg
cuxZRQR5BR4UipnBAy9MyWx8GtLrVMPlN+iRU20SeZhGgQr2L6aqc7r4qcE/avRpnl7kZpyTJNJe
zo+MyeVn/M8BsDUIEMOXcXamtPd0VnQR4Ob6t3OLA7BzAdlGlwWyCcOLqAEXKw81xdRXVEmz6ty+
pzuTOZjZnDGDJ9Q4BBmf9Ak6FnTZNmxz/q9mJFxawBRTukZ1FL0I03tkc9zKWX9TIXuOVEskvkBy
VT4NEZ2hRocFRIlSd9s9u/wfpg274lT+bcj5I3ApH6Lq6D7+7Cj4U8WggMKpi2a8af0Kx5UPBpE7
LQTwfpww9wIOX8e3Tm2w2bYRWbYwtvvMc5cDw1H3U4opFI+UpYu3ZE/Jir5u/u5+HosY9kkL/VKh
2O8/vGpTo/Pbr5gFmc+ZC0lH0ICKKBmgLiie+ImY9loxilmOydDA7AO73fPmaeN3GvYWv3bFL64Y
gXeGHUPMVuBVQsljggDrLGkBPxmVdY1KPtFj3XSo3ABK2/GBVBtC1ukQRbCu1yDVBtszoKBc2N2I
ENiFos/ouB2cs2GZO7ISAzfjAdUboNnKL4jb4glvs3fo/MSjRRbl6l18N10AqFa4NuGprVueK2wm
7PRBGDwLhR6BLYjuEMBMtAZ9WuPmXx2DA78TJfmSmBfRjzc1eJMQSa/DLBQxnZrtMG8ReTe1YaFC
TTdKr34eceO1fp3ke3qHHCebvp3EzqgbmLAp1E7uEtLkWEtfKS94dnZOoShErR5u+ZxlyLTnEiOe
r0cs0K8z2OsaRVKcpEE7LKt23ze1rqFu5IndgD2lNFL0AeYl8bEVgwNXryXOXrii8o8pHD62+Xaa
k7+//nTMbHgjtJJYCIRIBRqlk5dHU0a01iyO0JcG4VFayvqI9KCFGQzTjjUBep4WvILTsmcAwPF2
vZuyxrPmm6u4inyGqYTVfz+CYTfo5dIicbh5KcmPcsLrs+iQdoJrdsY1/FAAU0R6DNAvlJBPNvcY
rp+IG/VRvMykILEIAv93e22h6kjnP4D4Fvok6Jk97/Wx8tAha2T49cDzk9BEs6RssjZJ/+JHTikG
o6Q8P+zirWKKsglytaNhtBLfrX2Z1qCu+MjnUmZYKvP7oRZw0GlRKi21B5rFFrh4IHjwmZf5pBHt
cwNjnu+g3TtoDOm5vZJ880PqjMw9CcoeHb/tEPZ4T/ywY6EgvLqwNjStjMwsmZccX8idoNKW6P9c
dR83iT5Khz0NZLh4TaidHJpPZ9OuQs0up/PcvoCgtmuLcKUYYqjJ3DiyL2bRgKQGuPgDgzJE8qaR
WLZIowDSYP2MlKcrEZutKYb4tnvgckOzVWP2Z72KyyO2ugbcKqR+5YoETyvd6E7rjYRYdmVYfQGf
p4CW1FqD6UvQOnfdWA4mQ05CX6Ttp26/O5+PE+M01KovPmmgqb3DdW2uOYQk3kPEY6GeTJpSkb8n
zH+gmoOzF9EGwhhFx83cr2t5T70QRimMbtYSxyyMEmgydRKuBX3tTNnd2shhuF69usVrsslFHOfC
Yqp2LBvUdY7QVfbEORyWif4n6PN9E2niVRK8nQod3KdlAVxHNpVPLl55WyDgzZR5riKwOKyerlgd
eLxrVLA3AapqLLtMjp3mZhe9XvFvU7TEFSraLd6XpGHpzIHctbq+o8L83Bo9fwSBXVT6rivsuMnX
QDNzlGrTwcwHW3f9DuxJ3xpctSs6sFdrFY3rAfLa79fdYbkEDp6ji1Ac0KQZe1Zg0zDPF1o1mPTk
LhJzDeejuZghICaTCYMVr0YtFLlFCFi2k9S6htL2kO6xV1VE6V8Nti5DszETdUKGWgp0Wvi0M22U
Kl00485NcLVTZZLZ1/Qyyw8uNGI90PKPSJoVA3J7vMoh9YtmMpU3ejloCsjaYE5HtSTMFFO5+8Xd
IxXvmVLJPLb8WGEiDAa+id21gV5B6/HdCY0oQVLMma7f7gaFAICW3Ok5s2a8cENNNN4UHlqwjS/p
Mm57fe0plK9XESQIfBubeOSJu9J8Igy9LibumrYF/GpzTWp+uJP+iKsP21P4NXLxh++Om0zm+0P5
3/dwAS+Ri9DtdXJumOYttba8XX9CnGSsa86vaY0wtQSK5I0FS/kGHv7LSc07rHAbDF7d7yHJt2Hh
TydNlz6eNLUeErJgOXpuxfuDyAL+Wb4jCurRHYQjaR6doAFUe4vM/c0+Bd3ptZAXC8Nici9KlmHA
Rg9r83kUuTuKnT3Y5vOnHngefi3bbtzU2DhwB+z39RRvDMZeN3jgy1jW4b5wq2oRfgYzYUR05JxE
9F1dNrx7/aNX45yt4WaK0AHFT8iW/zxghU533kGTwNXfj7vTJ9xcg6AZqE06+5ddC9TDbGf6wTFR
/hXExPqRgC1FLuqeUDEv1KMrVQGwfIY4Xvx4cltqaFv+AOUeR3c4ZvQjg1VSps3MfilTdGWD/2/J
OIL4HW9Pn1L04A5xCwKKyFotgn1wGd0RZeRKYgfo5uuh6/xQ/wAg+18ynpBz9XUK6fY3AdMla6ab
82PXqyo8WljZUkS026w9UnenoEWgTSZ+3ldDVtKi1bz4OxyAWT3BnWybc3DAlrRwBwoatIQVL4PT
I9RXdf4HHcW2b3xoC9bN7Kjft5g+3N+CLXY+5ArFRxUUl3eNAlpDolmsATkN+myJWfNE0Uu0wFyW
9B9akFql6s8c0P62tLRt47iCEiPUTqftzxbYdXk5O+IbKScWgu/8Y4hhJsZ6Yg/SxjUMDMuAIQkL
ZXS7SCtwLlrsyG5holIVMSucYxUvbsW9wVdnZmqxxfLoe/4qceAVnj4w04eQ46fMVQBvc1/6aE5+
By+aCn9IGWFMHkDI9dfetT0sW0hHMjtTQloXD7whRmWze0+gHfz5UZOJ3Nn4s5M0Ts6J2OhICxI6
R67WR7r93GZtGKL9Kg9BASI3rlUBM/GjwCXtJC0RJRUKx4CzVzh9polARlowzlAhB1RlUd+VJ4eP
+jIRjgtDe+6UemhkF48XK4XsQme2uuokwgyD5bvk7neaK2Q7kuUye2Ybzs1Lut+oxd9JcnvBc9m1
/+PFDdZRWyBR/laEP8D1VpbulMCmgdTxIjE3grvFD9zNmhOgu4WGKnWcvsTlofkf7P/ZyNNPj2Nm
VBK1VfoIGGkGLCtLXqndAHm9/oXS7sUI77jqkrl+/kWob6YgiWGahpYBxq9ny0Bp6Q1H1KsRnT1j
aOE4znVOnPaslWPWYIIccweaNSblnrWiKM4LNhOikoWnLMtOx194gUma9K6ItKYFPq+KGbZexSTQ
sISDncIf1Az/7F5povT28DJCJKwASpUjuaYDYZzvHE0suOILn0IVvZYjSfeU/vKt/CogaeMEnPjd
3BtOH6U+s7yGALWguQIqrNLH4YozCfstNXy0AxaCYFbqDn7T6FGkT0h3f8vxeHbSA4/+8lIKi8uo
XhyUvcGmOsTbuYI1AWM4nuKhpfHOED4HC6e+rih2WRxswpBLKrb2ja8H7dzymfs5r1VX1uOIsgSG
clINle0rXAMZyvDXe8uY9c/P6/U1zbz48BCYyrxVZ5ode7wfUtPIJY1U/DUHw5wj6Rb/+mNtJl5r
ZUgig4scFmb6zNmGEKxfBnstFqtyU303MtYqVBGbkTxEnM1zWv8FQ8nWHVxViZCUcGluQODc59wv
y+CEec/7POg+VZ8kfOcs1Aqnm0Fg22SaZ2NcsYAPKGzkeStq4qf66ht/nsx4hmikvc5u8MJzQ8nU
NjddoYWI7vddcaRyfx3pubfqokprZBcDRohfUf1crX9B8JIRdEu9h3ln7I0xX0tVQG7g4i5LWJQL
Az7Q9er5Xn4d9Wd7/GlbKrby9MemOwc0BuLg4TPIKJtHpfqVRm2ettSQmHGp5E0VwMoJjk/wIo0h
TOKORaR6ywMI5PGjZgfMMs9KNgjoXuC2B+SmRJ7lwKsP+AruZMK8tNqNp7gveKZeybVQgn8f510u
lUpefcSPB+9N48xFr6iW2n2Cq9q8ScujcqVQgVL8kOjUvMOt8vEbDos6zgJCFHWXevlCIWAxfFKY
Ux+EpH3O6p1wDYgq+5PoQgADizpOeVHlR5lPt/VzeKVoiOjJmwmJfhIdDWDG4PH6OdPOFcMxA5xm
ZtTfCDSrON+AeVRk4eadtx+/fHK4s+n149YvH/DBba5syrscBk8lAnR/UETTlST2TStQsc0PpD0n
LJZeA7bs3gPkTkmOnMsqNxqP6qve4VLkZHtDsYSP8+XEAahkpY58M+ohF2fDj1SLOoxRT8i2/G88
AcpMFjM6NFvvWvD0jKtrs47RGwcXtMymabH/mBiAGrKqRddXxDtD6utPhgSAIhkRm3XXvF8uoatb
+jh6SVBBz19SnYkF958YYDr6rCDyzB1yOzRNArGv7ZuN0PW/JF5OzZRSeMJ0gKz+mjp8Aj13LN7R
SLS4FYWo4bIXRkuC06Dp+RSgrHRpbxY1ex0+zeB33WKVDUQThSdb8sKj4nCySlDUaNaVurD2zr5f
bscWgA2MetE/wqfei6Neff4gck35BG8NlsTd0W/6AirHkUy6QgdAtbU3iQcKp2YraH7h/je20Isw
N5+LLp/s5+fd2RFivniy+P2oI1cov157LJKzU+e0MXkJmTEf8NM7bi8wzwSLTwbM1bSGKqgOasvI
xXpteZILEZTfUuoX03tJpUCgWfdEzZeDnF7mlFWdZDJNDoQex6OUCq/9Ruq5NVJ4T9WKuJAl7kiK
Wh2zOdparJy618Bj6R2XpG0OCCeM1q+YFe997QpLe6JNZRYbunLG1VS+t7Y0Yun1ZguCYjEHHgr9
MYJekS6Voh+tTOFNVxcF7Mmh+Rd7EKGG9YilDVWbsL1dnIwTjP8OpwLhI4vJztsoLpDyKu320xH1
MF6Op1q6ahP9hS4cPfrMABebl4ubYggNdE9MjbAPOdyL3f2BWaIzL3pj1V/F/S55L6ctXvjXXTig
bamZRssSIk9uV7ckE3c8FeQbWYFTUR33WuowUddFHLCkVwGPjlbMwqr5CCCRxGBbtyEjCcV6Tt/0
i6UprI8G2z/GBYrELD0+bb9DvMMY/UYA7HTJA7UHo5PRZGG+1dR9YXhO+e1V3F8LgGJrHUkzogi7
Yu6DVABNhL4g3p/nGSZc3cuNJzN3PhLB366nDJTRR02B0vY38yJC5bMUscArjv03HPdavgnTb0JQ
ucYP685Bn2sU6B/yNPpXEf0VyjTz4hcXVhIzMfblBV2mdqNdtJwp4BIt8T8BSrlA/pY2Qp3XOpbX
HUpxQu8BQYA4YPYZuCvK+0bHCJ4dw8X5T7pR6Qq9WfnhtdzCmBuoSRZhBfr7IMSE6hbfhr8kdVTC
zeI+cuj2PfrJu4Myp+ccXjkLlg9MhHuy8UTTHsebJzYHKy3k4n7RBXmTcM8WXB4JHUQT3gE1r9J9
nIHTp2nGmASKEJT9KjBfoDBGx7R3n3Mb59mijeP1sb7Skawf3/ahsHhQoqQa7fH72C9YEumROkS6
VEI5iAjROfyiNKCe4lizrBgQPJm8TVCYi11xJmkLHXFpmD7K5G2fRaU/DukWateFxOLkfh+5YpxV
JvnnrhOYCgFAeBegfEsOp3piHjKuMO8wTMWq5Blb/l9plbqlpq2uq+RS86ZwywUabcMCIU8UKFdt
0s5bl+TPlgoXWSyRX7I2ZaWSuRowG5J2YgsCXQoZFtY/OuSzzv+j81/+SKQm6XW7hn0zxwE/nXLu
Xp5u3RN7FBsqiVbG2cZuFID0eCFSOuZyoGJJYNHWJlht+JO99L7FZ4l0Vs3k5RjCiV6ZsgujrfeX
XQer/nkLTpKyPpXOQyV4WNRp48FmM3e/QriQUEkDYh26JH9Am/APaGhHCXf1gCEH9m62v14El6ng
Ort94LxdB0wP2QTU2xDGJcCNzacqsvlxP2F8hkAEchwu3Y4IkrPAIrawdwJtZRnEhtHqR/kyk0/E
N22P6y2++44igbV68JtSt9SSuxV4VP7qvQiG+vFhPdXBYuwKKUTEVBtTVqBnvEVmxoezGpR8sC+c
lOnrylZ8tLgh5OqWeMICIPF+bdWJcV41PSnUlSQUyDAUHe9xk7NfkUjUZQzXA983c52uNai5ytx2
8ZvFq3DOcjnGP7DY+F00vsq9AIO/iepNxEOCo+S8hGqtDd05jLrRdz1xnZCXjED+uNYbTgbCq9DG
al37mLO3DfdN2tTJ3a9EtagwhwQhv+PfApX81RJu8TR9/v8tWQaHvR9tpKPetq5WN48NUk8gqRDq
oBQCNffy+khbTIN9j20OOjQ13+173h5eSWm1RgGESWS03Ymru7JiIRJCQoFa4X6+UnXhHyX10QuN
/OjLnS+S843YFOg/fM1D+8S4pFLBZ0XvBi2I74355RukvI3UI4vKPactw2eOd9QarHRqHA5ymJlH
EqGGsS+YJ0EJQKZ5u/E92SBiqoll8vrDfi4ZeaECeQbm/DfCn9sgtEiwodr52Yac0yIwC2gVEoPf
Z+0xs8WRHCgmbtiDSKT8umpUjcayPYdipa11eCMWmrg7o29u2Ll8DLNjuqId2MKSMqg9DyrzA/ya
oSPeYEPqLBJMm+0V8ijvyE5mI/PEkaKxxrPbRBP+qxv4kkWmuzE0FxvAt4sl2iMye/sohq4lS2Qq
0kaXwT/5s0XeikcS+eXJ6j/AfPhLo1MZ57KYj4AwOY1UXmTRMEQlQ8amqRWjNLYPU0W5Wrm7HKEw
GsaX3DigcvNGQxF/owUytmz082ONmBV7m28dQFezveJkMvGI/pIiut3D/OniOld5jNHp0w3xdl9v
/iLZS5A51fXV1w7lMsDDGbFvKKp8rMxPR/olPqwVHWUtLMldgvCXpFHtMOS8nwTL1AgrtqhgeZD/
HmmIIZeJLP5EVEXzY6Q9sZ5eDvoOg5P/Fhp6U5r2TZ79ui4CtS4yGVwVGt65dcwRVepGoQw5AadQ
uOMvkhuGtkFwqJ5p83VNTxH99IT37+eycLynF6W9ju5haJsaTP6Ep4BUhoQYH/1/RDtemdqPJIr2
RpXo6U/Yl3GZJwk+dr6ObVoCwFcVdGe1W8PzfjGKpn6HPZqslmUKpkaHuwqrYjdjsDZUxFN/+Nnd
WdEZG4qMKrqRFWSyvOZFMyHVoE8b4G+fZByoDp9i6JJNHJVjPud21DCVYpz4hvCzpzGsDq0a7DYq
bpd+XFmUUxp5Bxqdgvt4f1EyOFBLNNWIZZ+N2uUZdG0XXsOkZItGrzb0+k5G0Q7eWRB6Z328AhZr
8LLsS9rn1bW+Jk5E01FhlAL/CfkUC7FwofL128LdQ9pSY/8tvz+9+3KOA5hReodpcitghFmKmGE/
fc93BoMlm263ig7ndQ/v7leQhW6VUGTbJQVkevsvym99HohtBIxFl1A5621kcFmJV+Any4317Rg0
5hcerqbeEj73sDjKrr4zhVmNCIk/5/e5g6fZrkDHMud11USzWivFJ++PxMa5YN/Y2wnLQfSGdjgF
m9lPedUCiXmVbV/PTlS1INl8gOq0VYxtSOoNquaLesUj0yl6LzHdOOHRIiQ+Vob4rEcS9pWWFSry
oqiUXQ5Hg6gUuLoerRhhmmvPbEQi6NP1WbDjwhFcBdMzHtesyOVQYBWWCLjWIrtfHNdrT160OjzO
7GNkJq53xfjf8gu1rHOfpJ4OSTO3heUnC1oqs3VxbnrSbHCi7S01bcHxVtDJaL5e3HkN6xu7pQZV
VoHUrbWU5H2T3a1QBhiXLb1XFB/FvzCgAzfGzJAkf2TNvS3R/NycBoaOShkEvWEDSB3u06/y+RzN
UOwSt8/Et0GXsIPfPuNKIDHjBR4LZbvO2OgBu14eU2KzG/TNd16fsWpx7xCTZ69WRuGfMWRaoMIV
E2Qe1gsfcxkW7i6j9l9iQsWtS+ZEJ6aNAxlZVd6MyCQH3omYqoqcwACzvY72zJC7g8n622hzQDkC
aMIBOd6iLHRBm7rOiMZChcRdG1EaAqUHJ4YEdtQtuWHY7P2NzKcYPu1VnyPAXvjIYqU2CkdZVrjd
FLGdv0epqcTta25/Hc6DdqvYzRaN7gLHWDbW3Uvfgo6H4RkgX/3UI6jCg8I5AFJ7Rq6h4/4CS6/U
rSvWEJyPLb28rk2IoI/Atig9EuKMo+1UguUZGxIWvn0E8hSqG3jHzq+z9lFboCIPBCatp/xZLSZA
mAfZ/YCgakbUwHndpmgqNCQrtykAjrGo/MnnoKaMr0TGbwBW+f/PIjwz4JsRPeTKU3axVUC8XZ8W
xunxHaq7N3c77NkgtCYgup4AJV3pEWK4x9uZw1+ilKw69Qz7IkpnaZOibzxYh5YBFWI1AfnCupRd
gWqvWR9ZesJIqvIAHDvRRDXXK3OJl4bZZILFQvDSxhwJJOxp3szhVoubFL2Ox2Ez1jJGrq87qOLg
byGI8SSntzYYoZwK53mt1e3ZcnZB9GgrxsVaZvYi3A7O2V4KieomCs1WxaxJqRVNz6zQqO2+npco
mFzqTm/HY8RvzQDOARCGpniqraWL/CrduWLGV73/AT775cqmwm0RAkjIpuGieyAGPFtbySgPLsgU
0Mxiq/g/0pajQ79Ajsyv7CNm937Y/kRV16EEPZNBWSxcKgbGg1RXSaG1fmKWTPJl61DWLikwCx7X
bpqrR8LYrE3IqjKM2RCnuUxIe+9DF8xUz1yAzn+G1X1LU1oKNUqCcUqNM+sKfk6EChZHVNudPmvP
rfznm9FfdGmFDLu0e4ieXdhfPQF0Dq4Uk1GR6hPKhl1qn3bZSDa8LlezuaAZMeWKQd3wkG/hmp90
cUC143cOpPqB+fH70/4AR+L2vau6FJ28QaIgG19W15Ye8bfNIytzB1gM9Dls5VBptFMoqApxK89H
+AoGSLGMgdUQrPc5R2tug2Q7ti3F0/QrINYCZ7rLC6xE+YLMfIZ3B5r5mTp/ZAsmHV1P+/hFm7le
YlVBA1g4eGC61c4oViRH0duXiDh+HvoGEw26El2Om5Z/d6Y9ZcghEWyKadE9LodJjA7N5xmJ/WEv
sbCo5/d7b0EalhEj2xDHdhSJUnhUZR3y49TZUMrwynA5jN4RjnZl7R3IoEvEfXgVwuBOgcx/XZYC
8gB5hnIWrWIaF/NoicjHxj86IXsKSOytOBsHwRf14ThykdY+tNb/LfopIk2uAX+T174FdtQUPQFu
zstO3CAFkX5N3c6f66mkEGFgepPYmnhpFhIxG/ZApQseWI5NWXXT3pC02Y1dtxBlAHMk18LESaw+
dPk0sfNdYzmey9bKwnC2wiMpwCr6rNtpOAo0zP0gPgTnu3Ex14ZsVkHKOFcIfVJ5y2Pd3EPMG28g
9SKlthOh73bQAotoT6dPXifkUe5aUBTU0uUV7PpwkjdUTEnaKoglwBVx1bbX4Pr+Kf7mrZVF9Rh1
dTYTFukcA5IIKBe9+ebWS/qLX8iz/Lx/+6QDvFgT7Hdz/xsRq+hrBaTOyBZ+5ibCgUsOYLEAzAWl
ju/WQRybMlfCEi04d57jFqYF6f+n3h79/Y69qWAJLJl6lDJBAAjGpXJJ7i/i7uLhgL9X2z4Crkxv
ICN15twomWczRoBmdH7aLrFsQ6gRmm1pSkwKxiLrYxEa/XBtgQSROXMFNmdKm2ghTshon5yT/uti
YkISBKEbLjNL8lgoUy/iOgE+0Sb2YW6UoVMSieY0FRMTWt+hbEoMRUvH6qdZy6h69zS2Bdgr+DRv
L0pqtRe4b3JmustQhzNDQXfS822fJIMy2egXfhRqbkN4IZuplnRQRWFo9BOTeSGQWz0TnpnO/dtx
Ovtxl6hQ3thFXK0MrDoF5rVSEuwc/cVywDMipfA1T0cARLLd+XPYoaw0vY5Rj3CFWFzltkPl3gN9
ouqXYBUxqrSESSxY9TEGamOhj23rLWuBMHA7XVLG+nRNkqEMAZ2rx4XpEV3p2FrOv68i7VPEGLsF
+yrmpOG20e7vN+2TYud0LK9GB19rLiPxZCw9Tt+CqHmotjtFcpxEppAdqD4320glrU53PYJ+Tt4Q
xig10Xm4IEOahu+aM4UxLeSDPjhODirMLMpUbvT8P5sBv1A8kg/hVz/tyomuKZmFyQk4mhiJBEr2
DbBK8oWwextGa7UIXPZDjvqrYFZXGWlqYzzkK9HoyCCgW2AhIHFoJmoRie9Y1MYrM9IaciZZKInO
o8Fnm+WRRfldZs/+L/Ov7IweIoBKu0zOD3k3PXQzXfxg4QVUWpR3o7DzZL/RSghgWBxpMfSniCW7
AQz7HPqAp5yuF/PhggiNohuHKYSjCkFhBxvpqIRldjtm5l7Twk/4pF+CEKHgC3BSwyEgFEy14ki9
kFpBjH/ddgiFJXQE7Jz4p5psjXGFBwV/cUM+AWCOedA4xJLvjNmY8IueT+Ncspi6YKunM9lbpsUj
4kpf2j6PIKoBcxVd2v6AMjtsrSv8+ZtM7IzX/IZY3EtR2mnkn/0SUpc8SNz0HLV/Jh0mUUZBJe6O
NMA7laM9mBI6lHaWeRIenmvcG92qVkFdnx8VqSho6O4sjLggJCZ0fvsrbt8G+tC2U9Ej72al08pW
YPGfOXEQkxMEoH2kP1pvYiAgIcI01W/dc3TgfyJ7eyvrUvK8G6AmMg0Fh2pDYsWYoSYtwfhhMTX+
DC40w9uobK1jAoDr9AAJutVFq44M8JJe0j5HK9mWc/ms7Hk6papIQwDQOGA+sd3Dw6dvcsWXEtiD
wVUPAZBv3oxBuqyqjREFYitypQFR2xjtI7bZUiy6PTZzAySP38v4BDn//01xNBNGMjEhdy8afwHi
b0HzI4a8IqB8xlF/DMa9vSCqrgCr6+H0m7TuVG/MmQ4fnBvidnIlTs4tZRs8TUbTHOIhpaXYnfxF
tqbz2SCRtFbQbfn4Vm3bTOMLg08ITFEZQ1f7HNEf/3iP+X65BgtmI3RHTTi45OcwEUjL+klJ6Ldj
zXAxte3ZZPKxvhQr57uyLECZJqcb4MGkxTH36C21YQxLCldG0/7YZPBEqbo/+6C8XJlOei6Hb65K
BQGMfUks/ph8+9UqpQzd1XqWAJTV34f0Y6+7ANuK5/ibBrJqs1i9dKmUG/FQKkM8BCYnE16JNLat
/jOf7N2diQnV/g0JnQxYRmwaKwQVcqgmu/uX4KC1XCJLy1iJzObfGMnCydKWmdeRdvRpnepZREug
ithYATrNbqnkq+T1N0pvomjKbAySP/jn1vTe/+QQer7xc/z1E+yX1cMqivfQ5mTve+/zniTAWM5f
P54E8+GoeBhVsN81D4iwfSEgitVguK4r1ss4cGHXwIwCsuRhDsLZyHco0F+IuQek7q9dFwyxG+oW
7nlZmGhzIfHhznnlQaPms3T0V2M4QYDt31aqCF4maNO9b/HZJ1XhFF7c5yh9Vs6pREvvQg8jga96
rL+xBMCQRwSi9YHnzATEdwTm6onNEbKYmST0uvzlQc+o0jOheX2vWTLT/g2gV8jjpKixzcHLlFt8
fJPhmRqTZiIcJ0NLY08Qw/yruc2Ueo9nDAGpFxpv75PAO3te8gtne3t1TgOtG0SUrNokTISmzPUo
GtXrJuGZD828UqfU73xpel2+x4g9dCrQfBZlavO/2wK9eCwPLWkVkxOFLZ3DRSRx7W78E8InmMqF
svsknB+McnFTKgi+WBG7AFDkM8UeQYynBr+Fye88WZiTBWO9co07UAKZGkBkLAhQoT6m4eO/WtqI
9WoTKmgPz3Rul9enHILLQB9cJTJ3seRImPN9l+8lyXScTGS6o59Zz6ydkN8WLA3f8COLwVDixpqR
aaqAkHq5a/GXORR9lvX5QXqlO/jQXNRND5v0r+Yn2A/VH6Cb+wn9mMot0UuqHokyFdCz56OwjSCz
rkx103gpdg2SATZ6G4fZFLmSTblE0Ble0mLkUnQ3OQ78JCpp8TA0rex4mIV9eoxTNi2XIirgWtr0
EHileRXQ9z0l5uVo7115EKn8qfFk3kXqlry4+82J6tblQnp3SO7Z4vgctyQWa123CMX/ovB5IDLS
Z0Ej5TvUqZIFmB6Rn9WSpWst6qFdYOoxzcKTgSgyHR/CXJgpU59Dy+chGG1tioSQLAQJSd2JwEb+
8SY83LcL4uEuQJo07b33fe79sAglXVe9moqTTBuBTf7rJq1Rle6LLCFa/896gZsScdF0xU92JpbX
RWDA4q7s+po8ehk9vp4H8RDweOi1nR5hECH5XXmGug0mBfKZ4i7Y/V3yqDBA1//J1hAs7J6eLqjn
o6s8tJVbYQTZj4w0MKm20GvD5ezlcaFCht2vh0TVZqAr9IyFVCltYjc+knTonreTvnqiPguq41jx
KhxFOr0JtRU9nUpZMJz1cMQusrR4kvT4FrmOVzNJGjL6CcDW74v18nKZrDmnT87TvmbwljQe6lnV
REymTXisS8VkVW1e++oHwf1NDfAQuSx2M53fQjs2MoWeMe6ADBsxuPjyMpqqwAEQIHD/pP9HTJGU
5CezPLC0ij1WKJloXgxvW1o0O9/BVdBfVhg8U5mU9nCP8D5ZdrOMhzJdrdZLa/BdE58mkwAZMZ6f
nLwnfRdQ5vN9u5bwgqK9RAPnhXMbbdkO0mLJ68/Dsh8WkRr/1YSE7snbO7DAvwoNLsAuGmU70IoW
HegMUePVwQXAWyjtirBhCgmIDUvlqHNDygfxSTWiGegT5Sqn6UWBgX5hianjtBdyQbT6VAucje8G
A/fyB3hEBFZgVMgVNi8pzlNRNSfzkUEQhDCgVYwL91KSUEjdCFrpPgk4NrU3t0Wr3ofHJiswbL4Z
P7VlV2wD+zNWhFXCe6P1/PJzsYt0ibXiPadFsbkDWDlpbKRysBxjS/1yhiaPjpCxgK+dLwEcxLqv
0anzF87bY2AdJUOKL/zI+to9FbvUk8TBN15V/Tl/papvVyGrooVTZRxHB/BQDtTpbYQjSYA1UnL8
vJvfP/j5vrprxNTSWBBE0uEuZQWK0R1n/zOrViw3AqADCamNA0Pm3kt5ZAUuau/xyB6legDpzAez
u5xdaeaKiT7zLozQ7zOiFX2TRmm9T2jq8KPoZP+rTNdjK92K/c6ufxaO+vLe+bCrrj01nZWVnShi
2Oup/M8k/KNKjKa76Isbn9I1L/abE+AtSmloFPn4OpqXLxau5QfOQHcQbd5ptZZwdFXms/DY1ewL
m5luKBqEn9bGJbysqcWRTaBqEftQE4GC+qv8SI7E676fltqlpQSMfojwjt8W8W1YQU5gwAvRdLu6
gEKX2V9V/gvGaYFdlBW9J/sBTzwheLL0dyU9Uy0TSlIPhSaL18mNLYk6fefr0pNRJjJA+3HVov9e
/27QM1Id9P12LpQvnRIAwxa6MOvseePTe12SXIfiak+5wGdMpjvOQvrWcSNo1D7sqw0wFBC689BH
9VUpWFmf1T45bk6DDb+qTw0mY+AilVvplAM3z56mguFD54M7jK5KJGZWNlHv4E4Wnbbln/G1GPe4
8iOSbKTNIirul7NSg6uXYDWYftZKggQ5aTzffYJhU9HlzH/cz55oGiTC/pc+Sp5Py5ij6UpRCOT1
MtQdbboUrSX47TIPubkgeLHCut+5HCZwCv552sbvruROmobVxxuNrwMxmMbBE2FpKGHYzIB0qdXF
uOZI30Dd+IKpiBq6kyZY54dZQhmKvvZ/TqhBZpQ+d1WwnAo2UcNOSfVyCiqoDDr3OVPitNq42x9L
CMRc/kEk+fUqa1nSKelKqLNbUQqTpRkfgEUIqOJMQNTG3fIcEDmGFFhsPEG6YZ2oNCFxtfQAvKDa
E8LIBpgYTW31rWE4F+EcYBNcPdMMI1dF+y9ITWS9u9dwjzh/+nNq4uLD6NmapkK8zBakodUS5Dwp
gNlJ8lS9/ue2c3IeKzrCut1Oiawr1UbyZvgIwR+cHcPBECLSAGpH2chShMk8UlYcz01HWAK4/V4q
l9hhxp/bKY9Rx2c6UnPFBhkQcwIGo4jekSiL87Kp4rZ2keVUhxDKFHQyI11GggTtZ6+xIBDprxgJ
6HYmVipxZS95eE4bDgKeyStrq5YqrWvlq/shE1Kay81KnXqcov98NMpw4v7Gm3P6skSxi7QzEear
H5TMRlo0nXuQcFic1vGh8dWIYRjl3k8Xsyr3x89ks21bg04piSWpWadglTcsWGjxzQLFTKdILuwc
79cAwZP/aN3tzacBym17Fdvoc0uQvrfCpeq96E8Jnxzo52yN7YJZPNuxVsnrqe7rlT4QKzNQZRSD
c16G7nOf5lG5DDBi+QZBG5qL1+SKbkDgcdePLgdoa37w1qPFND7Tag1qzDUjaWNRYv3bcRUZESEi
AdGB/YW3cOCQyn4tduUj4eN5UAG4R4FP+p47XctPdf0BhIkMVNxN81gtWdhYouRezoPaO2HDeUDx
vbNHvUCi1nf8blx5MR3PLrLUL3BlSUUG5wfzP8aSC+GbufgRT+3fBK7osQCjOfzlvB68TMR7w/wB
K71SZbbEM2u+3YCIgt31P27Cr4MGhyuiuAijiq5gPJvq3ijVbyBZ7bbP8A7U+76Wbu06eoPQ8xrZ
xLqbaDY3PNwrWuyVFO+SANpJGdSsP8rIwoJom+Nm42K2bcU1GT+TVAlyxvObDQ9Aa/9Y4/Qra3oz
14vQDuAVn3XoGlQGY4tK0eEXXy/KIu0aCXINXvGpjDSSBf1uTZCj7D5aE/Cz9FzUp+xGY6fI8fc2
V2WaFUu0dvVy6cSxKkaBQi8Mg5e1UgXg57Kvi9FPS8SHAedz/HB56Z9bg5qJawgPtGD6hA1TE02D
EYHWHPoGDr9eKH5KcUum3ptSr9ZvULG2vrooppwP9awb+plLJxPMI1Utt0fbPP4dTriFfmegRgpn
w2X7J/dkIzk03EDuBxsW3AcjkHnlD/jZEJ9TpcJJcV8muIPFcckKeWgf/YB855vRL2sPSObd1ZGx
1NBpb96eF72YPkLtd5IvD4JhUwsAIt/N+NwIVASFOdqeKtJolaP5h/YIcNDtVqQYOXbwOO7gnPzT
mEykvcpuUK9jJ0AUAii5nmuq0lOrn3lbTA4LIIoR+QgFvZ0GtYJuhFiJbq2LQD6jR2XxQ3k3h0ZP
nxQtA8dBfXpI8uuK4AbhENERRsNBqZzzdp6XhtOfzepYOkKTmZWgpnPKxJZ9uFNE/6/ACQTUQB1X
SNBHe/lDTb5xpGyB6sO5Qnj0aClWsqW7ipsnEYiu5w8+iln/dxAOxX/Cu4p2pj+WETpysevMAIdS
pU//d9Y5yHkFzGreh8ou2cf19S4wscusN4GNXtQQ/r8/igo3IE9iHQ0v2Ynf8PJfryOD+8bWP/gR
rz1fpzFM2Hqb4kaT/X3vtzeSy5YosBjudkkfuG/BmTTNbkNps4xwOPZGMzVI8RaYvdTvCqu97Q1a
P5p2MirclizdndIZEsLq8OObwNMs9zySZ7F9kzkipY0fz5LsEEZI143Jz6RUjzEtt1HfW8ZUoB4g
hFgDc568O2vnJa5zWs+psdMT8VCgwX7NEbIWAbicsRIhqHzWbRtO5XOR8PL1nGTcnmQ+DCF85vdx
oJhOyQLUZJkKx0q6/ffP05+JmU7XbzZHRl5uHOOvEGkvZbxsQ9BQSNuHG2dcJxw2SkNqYOMr1yp6
/04T10Brl8CFGDd9gkPANP8838Lfc04pCw0S444V8hgWZu/cXlWflAJzVsfVWxw5Z0qxu0vpwKnE
0rYeKK8USJccx+IZJWEYsfD4YMFhc9adQKMwsma4yKDpQnAxrRy8hFrCnEfIm7+eW1cOZ8Fkec61
I8D6fckUK2C+ZDDYfx+r5WoGjPcBQPHPVSmfXx3Ln0WtNbC/rGYTMcaBGdzs4xwgPU6JFizamBCd
I82p8u6X78yLeIKC9AcINQvwWz2m2KAClqJDw6RIUIO6nUjQcYjDafpoXBNlINxaISXqR59Go1dx
tnTmyWy1ImLz7b/Om7xMkvovupMDUct52n3MMCfukc+KC++SLQEu6ZnHLzuYZLO6sUdKQpuKz7+c
AvibQuEYpw55knqovr2+o0yNwcqmV7BeY13IqSQJ1ozUWxXdteJ09qD0wMFMUPRFwlD3YAc82Drx
903os4pt7cmDkuhmk7zGa3t/BIt8ErQdiiNWsYwt/xkmvBD91qo5v2mYnc0cukmnoWEo7xLMFEsN
wbe0z2B2wQa1Gd6tVzXtDKLUHqVs7GqTwNUUysLJqSRWOYD4ij0towN0WisD2JEiOIUwWjxA1NxN
kOH97rt2v8cHKVtyNcnh3ixl59aQ2rD7Fqa7w/NDZwRsOGDxHwuZkUGjC71LxrNni6PGwhLf8D1X
RcrVm8feud4BLye0RsHYbPZ/kRZ/VlJ2UnndlH8FeTornbKRvhnxPVi6F3xqhMRt8zxR3lE3O0tG
Nah2jOqV6HGekeSzSyTA0aL8wX90eViDP5efgZeh4PVjIx57oYOTf1iTgueCbemJY/NQLkw+Aet+
+GH9/X77X+aqJV8cP/qyoazAnlwzV4ZFwK3DmHAAhI8DSkAMeP3STWrS0KMu5cjjT9HEijsGAac4
bBSl5UT9wLYrORGi4n3NYY+bRdeuj0Yj8yFgUHChfcrgM9GMyq2muQy4on7EOTqXlL48/VmOlW5C
w8Um0o8fDIthqrW2n1YSTPaWODbOpNqVhtHFOKQlNSwTpJXhykrpbR5Yi4k/WpbtuzgSyn1gJli9
Xph+eFNeEpTvPc1EwsXuDm6uPU3n+p5QGo2r2IAfMCNKchi7c4fUjaCYbvMv1mY4F6SeB+4ByNWo
xFsDG+A8wTPMG56KZVSeOk8w3eKnnKHwCZUlv49AC7Ts10jD3UToUPbsdHGBxMBSKIFrxPwvYa5D
CMpzWoXVQtTO+7mtlX4R9F9mmJBtU1n9666upBfmrzG7cKY1lU3patMM2v36AWsf0S/FbZ44KPcD
v/nko8hq2nh4NM71lwgeWqCzAmYodnqRMMtnVJilc5SFJxRhJGX82SNMfo3BpDlB/Uw2bzVfN9Un
Aj9oEs40xtm5FL+bvrOGragMEphWDHKNiVfXHUdU8wKXGs5dtq57e96EHJcG71F5e326F+f45ZdN
39Ky0fxSEojEf+gG4rH1TfZknY6UyOGQjePOobGcoPHTBXEM1YE8J6USndinsxfEpwYFjGhFxuc3
TW46hGg68QVrFKq5mWKETaSn5nT1fWVdHH7i7opJR2AWRqG5kTo3xT+DBNiyXHr7TaR2AyrCc/Th
0lqNIsiHTGk0QQm7XIT7ubh8wisTMaePcSh3iq2g1JFHYNJ8YWyrT0Ofdq1ZscDsnUZ+9qsMwEcy
pqxPJmI3l34be9t8lhZidpA/Axo7cUjaOvB+JdQ71PCnWxGdKm6WiefD0b5vZQj0WkE4BxGLBxdv
CpL3E8nZ0UVCBzR9Gm0No/XAP1/kG2wP6WpuzmTrb/zLsd9MuoB4fqvi12sJS/FHi6A170G16NS1
pcB8QMnWHa9RA0uhc1ZqvheiUNSaHpYXdHUi+UJP3t0u57O7kWWg8YtEH2qlcn6Odbo33cHwJ+eH
QutwbaaYaPF2LzKTo8UmAnSUtU15e7op3Fg7kgPXIQ6GEzTEMngL+G0JpYbCDFRnNHyBQqdYdF/z
WbZiLawCFbTtNuZIkKx6HNBRluSg/uH+GLp9FlmCy1/JAM/OugQdXVUPsm6xhQjoxnLh+GMEY6c3
gDvtI7xw4fypqILZFGt0LA5UNhD/7oafloDU+S+pbPmBGe/vw3ZoPVJ+Q78Sgpmnm4AUOhbGbwzH
SvjNqPnvKMJhkY5eQnTOCTK3Op51yzQ9RXWcseEulTUpdeTXJKTBMa1Qg6LltRl7f6+CFa+14v6P
yLL33vUfiW0/P1NpuQNIKmiXtZ0xmQWMZPh9aW61R+1AYI0FV1wyhUA9OIr2mFLL3XJl9Ij1GOho
oBCMT2Mac2KL7IwRXItOGFPzH7jltaaePWWBG6ICjt7iMYrnRc+XhtTWR+FVO7HvHaKiUMiq5Kyc
u9+ehpapgRBtFasmF4jx/2+63H/p8jQgQHf0fh8l7x0tZrrMOYLz+HRNqyiPNAnGapmoW+ck/B/f
NO8yMtaF5Gp5x7D1yHc61Kxai0Rp/FjeQ40cnK2WIHFu8gTXvHZD523rCXzGGQtbAv193LPVa9iF
qJsyNGirXTvVwy53BV0xt6oxtJMexpzWGozvGpITXojuy3hNTdsKtHz5xbH61JhV1eHp4xyJN3zs
fi9eledkyvsCohUA30Ygw3zWnr951ZXDmQJDAp9Xw6yuFyNmC6+KlEhw9NANDzA8AFzd2/G3WKI2
4HADk/jIXLtL7Rqe0lq2Z+L8p7BNrMhSEvmnMtOe+0EFKSlVH0WspjyZADZ4m4IK6ovNeFm+ld4Y
ixNe7PV1RkCsRS6+k/RZYUCYxWFpG3cRol3PhFj7dfhFj7XaApXTiczGDzSxWAq904Dmea4ryzzZ
0So3YNcMcX5qzOQN4s3XAxm/sKB0sKgq8TcTNVX8peiIHR+LK5/LPR2P2suGvW2KDUSTYwhe6fQk
cDPkY46C9MKDwlyrGdFXz/rK40O6vtoBXnYNgtF4F2v46Xz6tyKVz9ahIhejMTyeCYxNR3DnWNRW
CZBOkMQ+fqsrtEdswrVozXEFam+UUG+xu+HV8HAmYJ8uHvX1oOsUGQC9XPVhbOx3JXTe41KKW6l3
Snmbo1AiMH5Og3OUuzav+qT5a1RpwMWoxKddAICE83SKFCna8a+Bl29ECOQ8x25TkL0xjecOapcP
TfH/rWHJCoFUCcm4T7ERh5zZg8Ucmei0j5hhiYcIzuYc4E5f1kBtafVKIeEcNC7AtSZ18xNEk5j8
FOKzDnMQp61Q7IgX8KZoHikkTX93h3xiQK4eWgVouIF/+d0kit9wt57LaeQ8gkjy0am5hPO7t9XN
1kJ4wLeMM4N1AZ5L0UCO/NRMt61xOckiZCncGAv4S5j7jjCcVx1JrntDkqgrYJ6v/sGoXFyBQ+py
icFZ9UhY905IOd+eFdAxJi9oTLzZveSy5a+ykSFydzAHsmxBzN9HPE6SIpcG3RJ4tMAEtjSGRdqq
sYu9vaR1mzECLi0q97wC7ZJ6lazBJ4y/hnZwF21CL5VDI2ffsr7bc9ZKPyrDI6MzGUBDkIKI7LrD
gVKdOKZbTFNCTYwA/zvyZywYPHGoP6wkrP5w4KSJSHMq0aC4bPwsUQbW4PpSvNcryYjvNjfYsxY+
rxDPyHDy9GJD5IIuyoRn/fheNEI+wKonKGdvARqpr0IfAkErr+Zh8fnbUCIx6zodedvhKxXKcUkh
DzPh33ukwaoEHt4RRYdBmQ0bnbAj8mmuhfDJwyWuQiZLTFcmeGB+9dBOXOZd7UNs1XwX2mh8BeGp
PTri5e/vAv0n4kquH3bR8sEe2WWIrUpVP8oeCTksBVv2XeUBrZXpzfmNHDB0iNFFYFmYfGFF0dqR
dq7Mrk7kUFFiR2FlFOzLn09nZLFekir034vXSRC1DN5y1rgzG8ggGQmk4QA08jc3o3e1kW37sAYJ
CgqdCzw5M0ZwO+et3/uQiO8bN6d7l56qomthRFas5APjonM39Kp7U/FeAF+7fsuuExTohK0/Kg0O
58W9fqBTPocp3UQGk6j66PzKsJ7mssphzt1echgvA9Ljqmw2rV29QNa5OtB7R/r8xjds9daYhR7l
Ot47gJ+FpCbBGNNVmuYk+8nOsSpC3+yI1C9adxhcxwzJUzNqQJ51OdrYuhR9bR4Wbm0znDZgCJWU
zRfObAY/pCZMrS/UuH5hPXCgR0cXO73aNKfkN4f6D4x8stnDJXOd3LBKS0wSa14eGFSIoSEYie/7
/zynA2iQggSGDIQZyhA9VyycDeQZV+1Yc5iuiZBKCysF7Af3YheG0KOS8NP86sieaFp5nkUiN4dn
erXneX73/zHBopmiAccjN7DZvfOz/kQ2qUdkDk46bzWONGNPsBf+XhOm4xDV/z8rW698j+ATIwQp
5KbaTzwDbc9+A/PpOAJs4W1Vns6kMj2d5ALTRhGGcGeNeKea5PC50olNK1R/ESFhyvC4F5T4QTrv
YthSO1hrjpeRSn580iEJ+oNL9+ca0DXa73pNBXy+Q0emmKg/INV0DSK/JZhFoFmlXGK4ClH6ch9T
+Ujh0MH1Jg1xqbRVy8whcMqBxDY8J7GrKVdyqrwY0l5Wjek1De8xqmV1cCN3V2FdivjX/E9JtGwn
ztQUm4gG7ObN/dx6q1TtSaIKG0Q7dxOLlFCmKc/ZL2Op8+7yLy9cpO+3WBiGB26p5B1cJqGEGpFI
fUZptNa4pegl4auX+u7aiXSW5zPwl1/mZJjDq4Z8NlR4dKUZAh19PC8mFIUwMQBd07ORMRTA1ayW
6pnkhvw6FlB4WwfQVYKc0WW/271FRRYzOkxuPTF2YwmfjgMTLu5DNPkzrR6KhI5YDenog89pHPKH
vp9ckWB68sbxR/4BGolfS8fZdVL1ao8tzcm4M2Df6FylfuY+93TSSP4YA7dLxpZ6eS/LmPPVfkdc
fjnYvaMZXiSH9hm2DdC3UN+UrHCnKubxwS+XPh3+/ESb/mILixAMkSbSfnIgU78wdF9JHMTE8EYr
LyS/CMPj10/Xzi8VZoEatPRc8SXM/q7GIOVVZbZgdrcEjhTcMcOv7hfn5mEfQbpWOury14OFgxEb
eQIw3Y0ZmftgzTGI5DTF4F9x4fKekyIHz+65fX/Yb5W7KhYc+uLQIAODFhaMorKoDBi7gwziQW8H
xJtt/zP+Y1b0TywU+Ed2RrvfB0TIE0IXucmeWRxIK7DaRx8XD4YuEYQa/nsl2gvoZXz4SXReLUpw
5uwFeZ7aNGi0aVLt3ROfCs75LmjUcWC/BSm8rkitTdIUECmudhSgbSy4pMy4UkWZFGwYBV0Ln+5G
1uYNefQ0BJYKMVl/byVgHWnbQzeR9W83UPIQt7ppeJ0McsmfJNz1ZpAaqdul0R1lYDL1PTUbK4VV
RVzGVisj5Yvz1/NHu4DNvCz8mpVdiS2mrOPye3r5BAyvdnfWyuiJWwdUC792td+wX7p/8McvdhxB
KVFnES0f7USargew/ZnPH0WHxRjlFKPs1Lkg6RssUZgjHY542Sw44/EHqFkv7IC2p8JEpJyMwmdb
/4pQUXRnCgj/DKhEiBvO1FXNzRdkD+rqzcGzMq06FY68D/IYbfaECNkIFFbzz7U8ecOrmGyaTD2F
5mMCW141TySxNFPFLUjk5N0itJjsi32E/otE8NgrsZFE/mgn5Axk6GsaZDyF0VwmmueGoTvNqOjS
Eb1fV5pBuAGeuu6zjW9obWQqtcuV00PaGZeIpcxnAKiQnsKwBlm4QCE4bZR+oHsS5gIGbQKC9Ht2
e1l/rZB0EzSuxvRduD9auPM+HVXgS68AnyxjUlbdwReWjoE3m9JuFsituNug5YEMXd0jeJ9GtSoO
qIOCAJ2GPbLsMRj2ikKv6SQYwdU/qd2Ixjp/fxK/c9875cDPS7FcOm1fWsrUZ9SgdKJMRsuBIoi8
4JaaqPP8bqOvlynnf8+iMKDkwhVVFWPg4tBrwhAaivCiX3oJ06bz0vVeLs7qRiIZdXtzsswFW8Hf
CoQ3ryKalWv59ud8Ty9EUu2GA80XF9LF0kuxhg0HEsNb9iXxt5yniwpzx/EvH+XK2D14z+4o4P1b
faMRlL8GHVpbzenV2PNzyjp+wICWgAn18W9JpcWNhZBCX1/BmXo57c5YpLJMhdc86EFZUOFf1MNn
Vsif0mGalc9zzQGKNOCmqryb
`protect end_protected
