`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RRgUO8Xpo/BcL44aw1KNtN1HasyQDjwj0r+vLOCYFstJod94vn0FzVoY/YQo0icMSJrLfXPdCmPA
1jilC/3ldw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kIpeUW4JEd0Oe+O4rD8VscjwGfVQdPKVElKIlPyIElqFDJ4CF7ieT297dcEZTPy6eAgCP23+VKVv
7+UpgrLZGVNHI+yV3dxZoh4VhcyIQk3YA3d9EuPDOEXc0yIpreG9Gbym/T63w7Vh3vlPRddTwDBm
Th46EHe+eDCEXrHpY+4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vUnugk7iLlYfM1gYiEFmZC7gukhkIJ8LSI6l4nAp5BnR4qshOljGiFdKry/dVBhcxe0o9oVrGz0q
RT7bLN8urviLIKefaIo/tslA9yXlo6gs356hPTWsy3X+brhRMYnVDX4rT+FEir4XivATJmH27Gj7
2wtka1zDLFSGkIfzG8Odby9Qgudx7AusWrhloEMmTDm6Yif1BXSQsY+4Fb2/8jk+pbGrihs3ERO5
OoVa8a7UE7RTkYORG5HXF3l1xxdDSdIt5ySpwwBemTQPpREFPk51MYbxRdr0gQX45TZLKTYthDPH
C/yCZz9s6t0aPgCHFG9QxOoVrf5JuPmm1KuiZg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mFF6ZJKG+24YD8ncnmch1baZjYuOfe316H55iPSlVuXjy73tm4sk2eiT3ovswtgKn76ocmOETbVb
Yh3Hm4LfVrpGo4idExoFOMba3MQX0CS8bQeYCUR22ez9KztU6Fb11WIl7Ppu+vLZJREpZD1s+zeF
3doBl0DnQfbHw0FWL24=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kNlcgKE6UUql3o9A33/4Wxv3msFV8soN1LIEw1j1tepSwYOq1to8sXf96AIpguu2C/pFF4+IvsAo
/uXEITCLTQi3jUACN2LWwG2iNfLLt+hmITpUNYxpVViazmibidwqtZr7/5H1+cBzxLv/puc1sJpy
3d6toJoJKorFLhp9XapIM5bzO8y/k8r02Vpy+IEqUVShP5eZBRwpElqZz0PWvI9ln0ik8bCb4vLg
TVRBdsjU+27JmS7uy/VjbPJ21m2Lufd9FPkKcCxuorMv24g+TAIWSX0MnbOWC9daQgOtjw+aqZP0
N8z0Q22RSMtU6Gn/3PxNgaXxYofPwER/FEF0YQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54880)
`protect data_block
/K2Y2uQ4KE5bVtsBzPfkzDqOe0kwfv90/6oQbPT78MK7X6X8gX0sLQ+4MGFqvcmHoVpXlbcm0xe4
qOBW7qt2zVg/sSdzMi1of745dExed+015GdfCrCHv8e8Jj8P1uWxZsw/XAVs8FRnvVGaMN0tpbeo
ChIZ1UuR/T3vrzVp3sE+Up5v727FTcsuIokhHpJjX9v6lVoio8hdmt5ZyveAdnKm1/pHogUtV5eR
m9DcGwCq7m9O/0jaIVgq/cC9HNdUokkEDz7ftS3RajE1rN5CrfKdSe0qO6UD/kXvRyJ298mWjJRx
WjdExkYBgArmO5YHZIASFc+86TgsCdkJjv8WkmTtXm2WmFDfh0HLaYp4N6LhcIqJy9B+BlCv6GmL
erBZcGrQQIJw8P9i848qEwxFS2ROTCgTDuQCUnD7xgnSHvZbj8RYe3L1lPcPA8am3/vt0isyx3hr
1PTvEeonU7fobZv9cqE3/nnMNwRwQZfILNTFOYpQXPmUUEt2jWKwyzPhvFfImadRtrS3G1U4RNbo
Y953iXWUlIYTIBPcYO5Hvmcb+rkmOHR9ttXiBCZvJc6TCOW72sDM+GVVtMA04leXbJ44duccRWy0
Ea2wJjbEbL3GPfd9R/hA1YqiapZ0/5BQL5OmtejRnsMXY+0c/aScXrcNTuDPqV4AorgtkIEk8pFh
RurvOeZaeCvAddDXdfZ/wEaA4qrIDk8bh5Hjn1uxUULimOo/WCSPjg5/kWWGOgEH09meitOK3/vc
JUD1sl6p2HjPYUhDolKlqakXinRAM7IHsx0kPSzY0GJzXsA6/QhuOuLnbcMS4VeoS2hvuEtLNfgq
nJKr+3SPm3/5cc/yGOoSj9fv4S92mY4YpMIx9acNiAHgnwkquIAJ56WvFX0nAxHM1XsBljRa2PmZ
GBZUy323T7f+4T9m/4WUsECUTB+S1BpNd7QTQANX53j0ufRSrsPXEm0PHvuVnWTAqYLX8hbZ7/8C
c2fOj9D1ovn885lpdLEbsk+fgUD3ublMwcKgAQUdo+/DK6ztNjMw0ln4NjCekhSDGcWHfAadab9g
y+QgzAHuR7ev6/1r+QV8a3BA6067AzthuPJ2/o2Anr6DMz9sz23iX9KxDsSa8uVULfc0zvRVIerj
Vhy/tTVNbbOzYrL2H8fG3Q33brXk7LzETRgv64+057tMygjM9oWxy/srYpFusnkmmBQu386iIzY/
DXN1F3JeDyyl9C95pvKKCb4LVQ7iX1MlbT/ZaZrdBeFbG7ttHpM/7OwmP99MtlLtqkGOKe2CF/2B
wGi7ucSQQbbs1NeR9RBuuNspnHUPj0WoRkJnYvEn2oo9pmLdlSfP/ILRNqpiaQL598LQFz7Tzr+9
xzef5fZdpxUjdN+YoWsn9f0Nzr3NV5ev1tMgnjPjTOUKjij3XNijTYZenE6PN4yOfQljZdZO47tV
BnYG2MLx+PZVOrqFis0Dys+XYcHHeoD85fAhhN8iQU+qcrICTytCsx/DPoYSvsucJ8BXsRLq9Ddo
NGdAmjBRWRynnNA8yeYZakqc0EPpDxqNXOECW9eEqi4g6fY+wFmjN+j1RIHbPqsW1rdPDlxNxA+4
eO9r6/oj39Ee4exKhFkZ50tTJi6b8DIPMcpj3H2DldM97EYDhBVQza5rAcPEJ2KQC/4ppb3jyyuw
VHTA2/6jyOBkDzgmtxBOp1CLIkqbsa+7iFydBFl6XiW0SEdmqxg5JNU9nNxQEI2YKsmT+/UA0X04
URNecgoSocHXUKFvpyskWvrBLxItbQG5jathNcPMvDb0Z2PuhI9vaYbyi96b+Z2mJtymw90HBCAk
sQTAkOG8fQX6fuuz9K073Q/ZDUFgkSIJi2e5ObR1S8fT7pTEPjTyMoYlghbWdReV2CMPN3wBOOX8
LtFYmrIv3QYcxnUWhhjMdM0wMYW7TraDLP6JlbJ0vYIweTNcz83pgui00kMzG7mSEm/okvtq7uyO
EA9eL7OFp/UxFYmo5skqDm0wk2qu5XzUARoDT/xGxpZNTjvjiZrWI+VAkEgJ/4iB1UkrzZRzOsEY
RGstc0dGZxV/yzjkkoMNuC4cu0nVPRYudGDtJgLtPwf5ZlU3IsgtwuoPHj8SopmTEfEYSxX3vzwL
Qq5DC7XvnEmo7/2rrgGtZjEksuwpmw6jeG0ez+bCqQbFc9zzbrmVisWPaiesekKJYri7oWeEI+Tz
A4cbPUIuDE/7TZ5T/2ZqpsLnHQxyRa/T7SwYh1AKyTqay2Y4Hoq31kq+5okpphYtHwjPVY67yHF3
kvMOJ+5dc0bfubCXOnMEqOHtVqoxslBG+nT5ESxO6GagmQeI8nnPxa2Msib9Xi+xdahj9k0Ih3QH
meTz6dnTLu6awDouaFRvAKTwnc7RHBAb0/Vf92PFqZ8WWh+K0AYaq+jQPPNVjF6g5REq92WCXJ7q
IrMRMza8zU029Y9+tt0lL8d1RksCHoVeWwoWWQer4c/w/95+GAdM/f5MkdMEKDA7bocK6+gym+M3
JcfCcS2jHua1SaiXHlghAIDChTR0v8hEG59EUUVcyUlKVySyqFc4Z7lgLfxp5Un59PAGhyetH6Xk
e0ybJRlTaV/nRcjOQU4/oWoUE+TuLQN6kEnnG0ztnOsFgaKXH1TqCtk3h5WUBozYV//CJOkIVU1f
/Ko4gLd2mS8nFd9JFEFEexgjAKDBNXiXM+Nncimx/FQpxlDNjcC4LMTzatXTiwmsynZvJr4jpYA1
4p51mqSU2QCQf+nxku/r3L12aZem6xYLN34O2BayEA6jdZb7+YHyyIMYKO2K7xHN8diqCcC+BEMl
Vdb5FoJUeM6YwlL523vqrkyCQWuZGZgvyStS/hbMid/1wG5sk+jKd8a62QCAk0utIQFq2XeaAvap
2y0rGRZHK6vlOta2zm4uFH6dCi5P0bNKMbopzOe1l76HtP7vQ1Jj3FeVk6UB4N9C/N7sJTEN685V
vSP+6CgLamRbpnbTMMg1r3TiWeyjnUkZfCPloZdWwhkQPQnn9tn2mwL6dhzYLuYNyLn29fy1PNuX
KUduBf1TfrpNz09/2jXB9ElWoGv6Dxh60cxZ5F+3//65VmlXqNdeP+zV4RpvFE8cxhC76+w2Wj5L
X0WkppBqFQY8l+TiNHevvi7ixSGG5S4//k+dRKqM3IC8Tc+b6N4hjPH+FopiMagkkOzGUeRsi7a6
0bLcZ1UhzCKJ+7ZRHUFXIZtfumJWxuUQEoOae3ebw9Kj1BNmYQLXV1h+p12ymbfOoRLenbmNMOeE
vj0Zi7OzUIl+D/QF9d4Z7kXuYVkdSDsRfg2kqIYhAX8COX/0KJ0LN6Ikwv2HftPZoL7Zd1CCSJ2c
jpebKPQ4Gm7NPW8sZ1olQktbOLc2P+L9WYr+xmEA3vc/ajNU+Vn65ZbMoKODn0WU0L1xHwev4ZFF
dvOMArrlSlhaWsNbSTHqtC/kAT/A8kgyMpKO3Trb3ErL5+gvM0ocbLktQ8iKA5y0Obd+XWnAo2T4
3NANtcWlWiTWuohgtzzXfa+66JpIMInvy4qUN2vLSwfdtAzFwPXy0HQW8bOALv4S8mQBWWTYLhCl
OyNk9UHWad8ujas2mX8CBz2e3DvzsVP2C4zhynEwAXVgaHVVKpAMcYTe301sOD9dq/iVY6dVAnU9
1nzX1b6rQd9b1wZ2FxkEcg46mgCzd33QiH0gRlNvq7QGY5YkazbZ/oAZsMgUifIN8AVdsWB40NH8
r4XMJ30VSvwPzPR/q0GvZ8FHXKXMHQDvPJgVSw8AUBUNjhSPssNnkAnGOotE4mUWSCEb5YIx4d5X
tFFmXKQqJw8gYPKwwSGGsUuDm4Kg0Cgic/xF82Im5Re2kvLaggz71C15v1JLbuh1OLujf2z4TrQL
n649Uj2UUZgi+2SqgyqXAhD+N+wSfuUojUOdOjouM+FjYI02SJNar34GFTwXB2iTxeBO7E8RXJkT
jenXt/ZYx60Ql+IrAcE6ibzN9sYycJBGz1NxVQwJVLg1vkRZjX5Q0ke24DxbSTj1xlMHcYZUQ4kh
DYsyK63ONjc4XXhVDwKS1zCU2ZLmKAlLRfmxehepKROTzbpZx6+hKdWcCHUB5Ag0ri1rMPfcRenn
xK+qJrLJCLlFBheXUfEZK8C70yxy5MHDCbtobl71oOs7jOycecAl1ETR/3r6mQWUvcWcPFI+Dm2S
iNfkUcCbLczhq++H7Vjaq3y17XzyatpzOAnJo316z7av5hMDRNbeCK6CFmvJ/VH3izSOoSeyoaks
LB0B4oLjPaHQ8LVzUGdyL4r/9v67u48bYH1zyy7oHwvU0DfVPoPIAt8W1MXmpTAwa+lcgHBSpIWd
Cn6+sZdtswSIJGWTTX59HUMArXnD0riVqiSE13V125H9w09XFdyYhd8wt8DHByNN8VL6cx0w4TO5
ufpWpzVNeEaMc6gTYjY5GnL79iYabtvLwHs1oGa7ljHAaoXK5le3hLsMQc7fhEuOBV5a6udutW/n
mCD/Hzd9V99mvBemaNDBSr5SatLQ9DyK3x2W4tmh+l2PzW7sh9lcuMOVoCVdnLfBlH/eoLqX4JLL
3OVGwhzKuUAfpt0FCu6pknr/qkvHJw7JizrSEeF7GSGcfecZjZhrHynqmcdyn18kxlfvU+vlJp/7
uJ4hjeCGCbt6XG1OAUf8lYsXtyN+ExJnnk8gXNaVBqW5J2N8Kkah3dPck8yvNUdVE30GiujVOwG4
rnfYHoq/wxsJ9l/teIJv9ZXoZUQl7JP+0NskyerAjWyFlFCbtWl7Qyl2gE9I7b2xnSdIAGyJGdLq
/6myMOgHqI1IT9vWliPfNLIpM5ZDkWiUsly6c5LAHoeIGza+9vVr4ao+kS30hu0wHih9faWVGLWJ
HXd+Tvm/A0KAZ2Tm18HP3Q02fGxYDPYg9rxY+QopAufmab+7sNo0UUfiOcmgJoqgLJvPe6mDbYyR
wLRtnPFTfpGnOYMSdWyrtkxx158hIN4dSoV+S1t4ybwF090A+uQ/CFnIPdB5jrWD8VaeKuk4HziS
8VHFDD47/MorCTI6mCQb74RHiY4lLSSuZ1BtuTYGfDH6ZKJhYSRbkmPW5vgv8ypg6L4C+g20Vemm
erIGxH75ij6PCw9tWSHSl0Uvt1fDb5eKm+lOiUGGjOIXkQsu/CdvnRN3NdHHWC+7eWvmNIv8zUnI
bqXMkHJSPbb0/2m7fgW7XW4G0BRSgBpmMFbLLFs4LuXMsTdUXX84Wmdhwfwc4wVbE970BKoAvZwh
8Ej88jDDk1UEWDL4To1gkel/uZ1QgrYjKrH4B00JqHIltAvQAUklI5J4epqLIytvICoQEEtrVmts
kS61EvkteoZOecn6iuy//LOAWjUvLXmP1HjMxH0bqFE8mrIuaZTjI3eSjB6U1KVTJfvsXR/1PDYF
ZLk32TxJZRZ0dEr93R7scO1yJjW5am2lt05Fe9kjvbWbRDya3gFNMkNGRYbZ0+7c9IfHIWFWpIib
mMckyRNUeGPy0DFsKjLgjwpICfi+bfpH87cjaTiShjzApQswJ9FLfqHfZrbFyOUQF8/aJq1BZVaQ
OniYmU5Jj8/w9vSvogmDLf/uYXrCRwAhQtV57AI7vecLCz9oLIj4QkBko1jHAhkCXhXkPUKzycz2
xkb5tWp6ilBZk9Ij/GXgngLnGztbnk9wMlLFgTAaK84Gy2OousQg2ZomA4VlHbDBaO82zEAPmAPn
cb+R+V29ESTfBSQ+9I4jd8G7AgoxM148RgcIaZNvyYWfn8jUk0rP9JaVCk6c9k6SqKUo21CwLvvY
iy9c6kX71KWShyWUOPZEhIo9Xid5cGuxg1/jLH6BrYkYyN4R2CV1CfsWTo9tTsBXX4f1fr5dyTzU
FXBTp59VpJ1bHWBIDKjTpQMMjitUY3dmfgKZPfbStn3/yWrsAaflv0DvrahxdSyvvtpIAvrYI0qw
XoafTMlDgs2eY0TFpN8b/Nlg4cSv7B5DnmBCSUldXCjHSeckTzxBhpjv1cw/7w3jWOj7EkxuUXPq
q/1IhAw+DO+OV64hr8aGSsEXfWEYbeSrtI9hSgpHicX0bOfSxkNfOhvJWTJPqaIZuJaPOnmzznX8
yspEo0ipGrR1w1D7IBSkTgbVODoa33SpASl5Fcu9oNWXX1tRsIYKNMI8pZzYadD22rkrdpfqCDZn
GjTzmN9B/gtKfzEOMpwKBTmrzBmEtrSDWPl3qVxfWh3KfcYqm7wbUiD5aXFspAC+gW8+f5wijGV2
fOvrI0YHxaEpNXq87TKW5/hBoNcBTbYBAEJatgyd2HtpNwc3LQX4H9Krplv2nWHeuZrSHi2UWnYx
TLgU2YnVU9QdOEWhQGbhgdv0gYF/fNDbB4FEGrUiaxykTEYbGdWpCG5xTj0M4N5s7Rv7ZHIWnk2k
okE8R4+YRDwXWY8SOZo/AHAumDle7K8ctfUDXrip8oPbBOPx1oKy5TPAy57yLi8lln9+Y/cLZIQt
+Bv+NZToV8dfrwvqD53cQ/icADsYxTsKJI6KEW0GRzlLTzHBEmPgrIO2njR2gZ4nqkiJ2EVAWmxg
35/OtLo4cx+woaXNUWxTPhorOg1shMHkNXGdFgeoUKBhwcXZiInfDVWmzxUZr3oEu/KXEMsDcXFt
ihybgWR4K9mRWEvyggKMiHimjEMX4TTCefZa2SX+lPi/RHZm5THbEhI/gE4OlMxGLwUha/ARJD9L
DQyFnl1qsgGFCbvDxEGNwZo7bS6BtouSJCBCMYW0lp9WQZdj34ViqfIZ2QkaezZij+33bMkzODHD
NYBjRXHquxdnYuwmrgY0ZsIOGv3I5j1JpnzC3h+zfT5X9K6kT5yC3DzhYixVpLXK2x9Doiw579QQ
BmFeO2N/P4LFatCAS0KLEXftZynXPw4CJwYdLoyptpz2hV6y7Y0UbDUjQV0HWjqGHESFBi4UOMf2
00yaNlAw+gANxz6g0+wcC29oQ9o6iz5WynvPioWZbY+SSmtzN3Og4rbbeFC6hswYLyZn3aggngCh
Q7/w9ILONA3/mF8cgD0Kh/i1D9laQVFgzwNdJtef0ItLRB7L10mBPp50ULqGVRgw2EEcqCiwCMOh
jp4eXGOQc/fy4CqLnE635kw5VOaLXWnEZdQedukpowV10Y+1lXK26q5OYxy/IN0l6hZ0FjYkUzhr
pP9Ke66DSZSy1eul7jnKAUs5RFxEkGPsKbRfK3RX/epZNS/IdzkM22CYr9G3HXXnUwGDS8P871iB
EbE0Zr5EDhpdvFTRMTK5emOu65aQLvC7gc3Z/GBZqcTbM7fbiSXyPwWY3O/u0zM89g27QB17myzg
GIHtjP8UghK4ClHLu3YJitrMLUWjRetvVnILAIKUnf5G65UuhmT9l0ozyNvIpAznhGK+bn4khcR+
bG/xDeDAhJIjQneGFoyuio3m3FiapNj+LgAZ05d3GA032HoK/WaqnAxi42C/DkDg6rMU0t/0/8wo
RV99+WcCNfnrINq9wpoKOMLh1Ru+rtPtai044axcokbbG6PgsoGYfOinCpDEyv1zt2ujGWgzKdov
zFsiLVOkJ2vi5x5zOxiXVWCS4ZayXjSD+T5jcZVKudkRjml8OzX/n5qv4a+Z/8w6uzyj/5jy4Klp
4hSv9wV2HGYv8zE/VrgDgUNH+4a9HU9DK+aAvDCAMuwHyWFlmbs0z46NyC/KaifMJ6VxCSPQdIyJ
bC4/KJNAP7x6E8VtVwAMoWdcCPg/tea36Ts9Tt2FkwQnMEPeEJeDiDZ6gNNkBKtnAwMW4MJL7ZHp
+dUbbF/xEpZls6x6Zo6+zaXlJIvDR9ohwE/fazKpW9msGPT2AzRW7KLiI7Yo4m2XwajlrqoS/nHn
yd0yCvpeY667aJSkET5KdAJ9YFJsQM4REYo6AN4fE9OfyQG7+2C/hXgVJcDNfjjhhiZpW12OV13L
Fh6ixMwAwcQkpX6U0z/cypPQtrS2lv6MeArHhAmZamb5SWs/+yBj9+gn9QOIUNxvBZlHST4tMVyc
x783+va8S3faKkmqaXBwP6cLmZEwPv4P03wwiTs4XK5SOaMOBssl1o9lqxy/WdfcBzgBiJsIEXKh
2Jok2tjbschODKq2vRnVxBnAgWjMkcNTVBjY1zQxes/Nqr8HXmtkuOBfVfw6LPGtVmRtmaIyjY3q
Rzhk3y++eqGmLCZYCFE/x79hA7nvJU4RDcu5DDijVdIXuwdqeOH7MGeC4hF/O54Se4EnzEBJGpBK
LBEhafDFZ43Ct7cWkoVaUWRRLxu+xCyQysAz2wnRVuKCL3SDQ/AWsiIeM7q2uQXPhsZ84xxhy6lY
dey+8DV+Li5QTHCkfXDzR8UJL5hDwGKXKF5sqGMyQCvX7Zhau8N4uTBZZOTDvN/AHAASxo1yTwMA
gVjMj68886JIfhg6jO7Sr5xLtaA7+cYIVpxY6x3G1Ojpzh1zUNhdjw2/AZhqnwGP02buwfxLPLso
f3tfUmoP7YwtkyVI4DtiIC9PCYU+qysasgTjm9u0RNd8pFehfvlb32tZ0WpFQElQPCIwmy1MZ4pw
szI+kCBPr6d+tKwf0De2Tw9oB/2lKDAQRBC8bzDejSMWUOcW7V7VtWWLj6V7tWIoBnWFp4/CHsic
dk9mTOcIFzFJQ0YgMGZ1edugL5AlP1iimHXLK17u2eYefI2y4D4u8ZiFQHDyjn3FdBOh7oVy53QW
2W+Rm3xD/KjX0vA3077QGIJh+eNKkX61/2sjZubklOk0+Z89dhkDVSqcZBnW3ZDkuxbuWj1wQQ8+
hmhssDcceZCzJ1HlxxkBC5A6rC/C0npYtywokS0Cei8WgpVxrzq6KYzQCZFcdFm3p4dZ0FxAm+GR
XmPWfQNdizYJ4v8E5PqFOyqXQ/MDaqHFKqn7O6ytwkm1Y7h5b7CIMeyvEO/45K+HarQU7QbXMxaP
W4MWsGvUfkgnxzLafIoLahAK/6BNQzX+X/5/R2xSa9h1XKHbc64myOlVk0wvtpEFltMSnWC8c0Ft
lGuWJEMubhdZGrEgTQBk4k5W1pklBIvpT1WHpighjsuM7JllvtTMZcNJ8QaJd4vMjcuLou9Js2KD
Z4bKVxsgyrbihwEy/svV5CnOWgkmjq71MUHH95c0I7G0KNHf8FWoteERc6BU0KceeAo9OCl16EeE
KSGyrjCh8wm1Wb1wPDh4FhXczCAgSz3rJ8LutNdqTeUnYmxLVRM4jRsO7ve6qfMcfmEwmT1QnK4O
/KnBXEhRrqy88TJpbas6424MmCSc/T4sWoUzAIHaz1EhWEAVrmVUobor1T+SYVD1TMjF+d91FrLu
aRbRGQk5Diad+cWM5SZUmTw3M04qk1nRKUE++TYDyYgNzPIz17qD0+EJMDmtPIYqdxbvwIrDUCST
OdIo07HsSZbi1eIGBtxiIgxS4+dJ0ic45SHbI/TdTqT9OZ3Tg0ihEb8SPxEI4RES7lDZ5Xvvg0nd
eSs8Okxr9T3m3yHwOzDP45LXzbIPkF5RxXbBqB3tpUosHGujqFbFpxz8baC/V7rtaPKXfGIx564U
yjzu0GgrN3x9zQ17H/9OaKnfM8JUa1OYM0CrcLaNp58RPzynetDS3cZKdpsnnwB1vvoLV9HUL7jp
cgClIvGZVwmRAQto6bC/XKmQZe+gj7oDtAUQrEe2aoIr3hRXGV+mSeR7Kjm8zrTa7HzGXedLsh6Q
3B1Z2o+PL+j6Gktdevf1DpnBSzCrTzX/l7q+4iapCBN2XarXlrOmXQtMdS9Qk+lj8RIfzWeGtBdR
XyIZsUUGD5sbB+eJxnq2Djquu+1IC1hm3UJibs4ylEXSV83hcjxF+S4UU7xM45mudLI5cZ8WgBfM
z1agQW9EB+AZDbyEpvGwkVC1MMXatmSlupn2NAXsAs0+C0E5NC2xN30JXWZdacBG1ebF1MP0zKLJ
0tFJg3ZAUylHWrC9Jl5C5/Mu/G1zgS14QEjS9sEuzZh0XAeIY1u15rW79Bvtrly4t/pwlpMtAqdA
JYZM65w+iDceJmrD4r8/ztMicj4ZlxJUkLNH88rhnRqZs+NTyBOXazcsZ80kvDuZKUA77M6wB3Xj
tll8+iUEWH6c+Dlb35bUQeoVNbVzbOjBznkOWgXV6k44XsgoLXq4eTwvnT5WI9G3zxM3MmjJx+WT
DDumiLYiHnJWb7hpJd+88KlZj7b81+sVeslMBYFEY5kg4kUcrGbQwhxCY1PITlUZZY13c2ht7109
JqyrZAD+L9VU1Koivxss52YlYCTI3SLWBk08PRRMmhUNsI9BJJlA+kk4FVvpLhOy8c+cNjzjVoKI
YHsCYbOvRTYjlR3w2mKyfSs+HvliV6Y8qMnPNjC68J/I0ZHCCG7BWUWhoVZCwRg4yo+b141AqWB1
6GUgYHY0oYVwO3Il+amressewROem5F0Q0dgyPXZ1NMBp1XaHErAGr9XMYEOyyZ4jQNAeAcf4g4b
BsKUE5vurDCdMCXvUHQCYf2Eq0/ZlFjKszuzhDVSoWpy9T/N8D58UHIx4+kwcqoXDTWS0Y6thSFl
UfXigkSUPPpVfWKwbzfOJqCM7r9h5Q9Bd++7fI3BgzBAVpgeFVkNBbmZaCfwfn5mdMONEhHvJWUw
/qz9hvlPAZOcwQMO9vrKNOjNyGMtWnSiJeudom5NQd/co700uiy/FZ64PEmuXbT5dv9Hzz3hatcr
UZNa0/XFwz+Ck1mz8iyaqUUcfvxfvRnKEJn2z7+4hlbzK9gYDLRUsU3HDrnRvVqXV4JTGj3kqBEd
Ga7bPZd7VQySWtzRJEtO4dUXjBIRR5ljT0OkBR7tEBNvbldOHe8g4DBMEqEbi6MV2EiBwAn02+Y1
+U55gOjVJjzv3aj8MqPXIVjNUsL7GprrT8evASl3kgy5J4u/M6YrqdfpWgnp95I82eT4urWNiRbd
we4v6lcVzsMPeqFin5IKztTx55Qu0OSTGj9l6BruY16vsoJ2pw4j9WN/PWzhISKcKjBK9mSQ1x5U
1V+gMhc3G+S+uZ1nPxjjJK4wT9viou608Y3cPtoMRlUfpDQJ39Hxrnsxvv+43HAc3GDZxoCimnf1
4pkCxNCI47mAOLVPrH+vi9j922A7j3v/+5aZaF9ytNSpNYoiXR1j2c1BqNfTAMKo3zHeLObqkL41
j4rW7sdJhtw5pLchWBpgEDcobE+mBhjBLYV1GydNbO0LkUJg2Egtyw41IOzIkCB4oDtearEDVBZd
RS6abGn/T19twFGrlbvn3OAE6rs41vQv7KRgvUX4vOkyBwKcLBWoOXrOxfbBxBOTyAZyPSeP5zXA
Mb+QuVpPutIt6twQGmgak8+7fMG4yDfJdE9JEDlMH44FhmX40sTUNV9N0d5+QWGThxIaYggs0yaK
dDryEkN4aCjp4xW0qooOXKagHu/GtMLstl5552LfxC3bTcvXNmps1xzNcJ4y/wUgK+qM4qhvYqCp
yvbgGQVsa1/ptwPn84KBAvEGj5j2sP2Wqrb4fntX7rox80VscTIgue9x/+zZM9i40k4IJKE5vvS7
0I6JpqSWJ3uN5w87U+WXa69R+/QwW6FvtR4XxupN+O3RJ0I8g41MesxbGqQ0N6OPMt9u07tHRXjE
7gLbRBEZr4hGpzK1DOxO/0eUq8HP6YexbUhDbtjjvyvd44aUbGT49VqA97UjusuU/GBSK+VoBVbO
MFkYGqmjIUAVBx/IBTgp9nUHGEA5niFkh8qHLRubWKoS4aBwM+tjyoG0Ylhmbxo1yY50/km4Nue7
b2ee5ko+iBGzVIfztSY2wWFzlboICv4pZT+mAQSOWApjtctqOcGnvNjnlVLndjWvfGO6JaC2A7QH
mVCastVE+zDVG90Y2vRrVOM/jn6LA5918AIW7JEb0zgb0OeOkSiO2HfFzcnAqJ9E3qs0akShbKUw
YlEje0NPjUQPU0wMSDNcsNck/+6rI5Ha6ugkKdniLxVIlJ3UYmFaVgrmKkY10docKmDO18XzKSaX
VciTMe7c7sF3dGbPdrML2lvVxZx33fke+tcKwwktSypG1Jra8z0HVkTYAycAmQUE+bswcG4ipU3a
Ols+iTZiqXXkdzwrou2H38vmivPcdw5BfuCHD8QlBAByoRm7CWyqLctWaAGF+6eQM64Oe8oA9lKJ
Suwl66E92QTncsPVkk5AMXR/ofdGhKvR1swUzDznGwBC/UKk9MBD1a7ZArHku1RZu/6nji60vV8N
scKoO7uWgs9FrXHvaE/E79kbwAS1R4RBcmivW0y3zu5aBwqFn8xuQndbh9SzrtifrpMUzSNSJiZe
RT3CsfTTsv+sOHAozta2tCm0AsRO7rB8emEvlDRnCy4x2ZJS7PYKipt80c7rAOCyCsrFr3lNit1V
UI/iZwMvznjOomLktPCu8uP1CFVb7GyzVcKiBFmd5E1bsk8cQDw0mTklyZlcnVUfZhoJ0fjsaoZ1
FBtt2h4OF6FqBtpmpQAcHmUH6aewn+nqCNFXLnNgGvRlcK45UibBXZ07kADBLOQcCcOijEpB0AqL
jykL/Ha0ybqnFnMrKi6RQXYnYCpMIKmGKVvlTXnUDfuOrhLRl8QBizhUMTSW6AoNGC6IG4rOUJu2
zCS3NV39pEf/WzWe3B+63b6y7WKM0F7qu8gdenktPcEa63BHpZjyH4pRIV7vyUqjw9UQvOImWq/P
WsPRfZcId4DFCc/AbvxXQz5gLXOI9ngdou6zmsp8zKJlS4BKLBzTGW1yjO0Hz876rWRI1wgHKwyk
BrYdXgz9QaFHjMTPf3UoIqlfXRR19U5DxpKzqaouP9nnyTYK+75QpzK1nQhK97IMr0fVBM1oXqYs
riQkwyzJ/6VpowAtPGnw/YCUEOQuzKi22RYXt4h4XxdhQ3bd9rmtusASuj9rkN0GBskMQE+gX6Hl
FbejZYHwAk+c7FCoqJhvWRmr5GymtZ0dIJfL0x7lj4HXbnLWGCOmsaVcHsUzMlvggh/9U/ZiBUt0
3rlq3xf6GGp/qwyKDwSnszzfudz7gX87FG2wwibK3Ulc08sNTbMEXmq6z/5EftGcu+hmWf/q/g3O
yUCBQfrxYp6KwR1M3hZrcbRfB56/BK+sksxXuHDNL2y1JGOVtHZZobTR3Kg+/CdbNM9NY8MjpDFD
O5JmoZlaIlwOuP9Mq5r6b7IDbeVq44o1kOetUOg7FRvnUNqMczbpWJTrp2AUNhaj0jpKvkxizoSp
8I87nw4eyqVPaWLwub6R/mUf/IeUGsYo3YkF2PKqPs8LPTQpj+rjpEz+LycYKO8blybHnTn7fMqP
pCdkc+pcKYTHIVVsprNYsqRoNWPORgxjJIi1vT8HadfjDdaEc23cDOQFgE1VJqiUXPd9p4MISfwq
O83LX3rxtz4SIHVxrydOXGs77ZZj2sJ+4h7wT2QZW2VZw2oZ42m4w9+++lfW/llYXllEOyTFtNRT
J9jTUgsevtzTva6V/PpxKSKSaHMJ1TIbVRAAo3RaKsOV1M3Lx+uVRYVOqZ3Buf1JZ75SeZBkk8H6
UE1oL8QIBf4ZOCGSIpfEZOd3PE3qPOXWMYue7ovA7I5t3PJMt9woe4lfRd1ypXSisLPJKdOOgfPI
9jIp2Y7uPCb3iiyKe/YLoJ48niA2qOG4BorMHkyf6Dy3DLzcNdJKGvavOAlQni/SD6x5MTeIJDW2
nLnXp/+BpoZcf+W8ljGML2xGt6WOEXOIcvrYSI7WfV7a0h/YMXLQl7g5XorBAUeG6DfvO6eApbCJ
ctQnEuOFSUclPAf6UkpKU6MZtV6LtsXYRbpTm0sOPcoQobVZcdaPMqdZqvxIEDdYias6MecexGV/
DOeaeFcsqIMW1yijRWkmVIy234ec5XeIpe/yWpfgEAfRS438m+PhNmpew+PQeqEmtI1syfGV7a5M
ro0Jb3yE6s/7zWRodgCJ9MxDYe9BVsmMsoGIXyHosjoOy3LD08DVEYYF1h8xWizMuCnWxHYkrCuH
CtNkxO1il4HpgKDUl0PGszr7K4zABZ/1Yy8dKMZtRmUECRu6uqpxZJK/TYUdbrI3TqMo1UBtayXn
0hBj20+cg5fZyaLD49+hhxSrCrDuXfrYAySfLpSLE+5jEEw7gsQ56yh7C5KKofOz4aDbaVC/1+Gj
oe32Gssfwu5Is1500p38qaMqWO7dRYqCllktZFXWiSeTxFZX3ZelT/B0cdacIUNxyThjM8pygWJ6
0lqP6ZfuDtFTZQVem0bB1FQ40ElZ1IJPI/01L1IQIKJPcctknEycZ40/Pa4W+Fh2FyJG4pOkj6pA
SeCnfP2iL0QBT4rmpjq87gNakdJ0jbKPmzIyg+Q7m+iwjjzHPHWO4Xl1njOk/DYZ9IbxS+lEL4wy
z2yYwa94u3Y6VAmdo/JAfQyfv13FmLK7xjFPcqRU1fsDysCSmhvc8fVZAN8uIXlnOBq0N4FF+6oj
4pzdp9VOpCWBfvEKfql5FdU01es4BlKhJbvtBuOhGe1bOZAUFdX8xNLxVy6vQXu0ze089vQeEY53
959qwhORuk0kov+rYTAdaaRO3eQJoPqs4ow9mKMH6a00zisExFZU4FhgvZk06LF7IFgfgMgO0oAC
OVkiA3PFHra5URbd5Rn/QdaykeRNNZ2wxsT3A4VJTthZUB1xHm+ofsxv78hf3OMMt1qRZ8wwCjr1
eSEETQ+oW3J7meyzEm84n1pGL0kWlCMkxn7S59ixfgzjmvwzVmQGYxrI4+DfslY1NtiAdQu+EGc0
m5kkFeYiAVnyf2zbJ3kBOEZaI7pH2lNcAcWsfFuyXZP4X4LV1qocCQxm9gxsQ+FdiUMKp/h7ikzv
XsJYtJSTvCTe41dL6NxL4ABIek3rd/WyZiZkgRI8+RQYH5Dk/a7bj+/+BejbDJ33Yx1BEul28x+h
RQO3OPdmK9AkeMRy7dMH3tD1AW9dmt5xLTvZtHefq1cEWSIBM4WzaolhXy24fQPpgiE5Q6sUqJsW
W/l7UM8ERe+LPd+aRJAxJ96jJIrvh8q0X/A1SNkLEEm7kcyrt+GxDa/p9//MdS2GoCt+Tl6nqgE+
JNtwiox62B2MDGNrw3JJh2ghefinMTO/eyTA4e8DMaFC81p/SQ7AFPj4pyl5CAQZTMS1qVSj3P6U
jMlEopW0ryro/aeXydlUwIjdy8pA9BnYGVxCibAjQhOnrPMJpHDB9Fmu57gDQimUiq8E5KJNjT45
Ghecn7S0/KLKRgFIjJ0KVLWYo0O62aW2aioR40nJRpUQN2QTtJvoAI2NrN4nre6PO9kEO2wzmtSp
NmNHSsCpS4tDm3pnS8zlql2JGdxxish1jZHWJfu/HKSv5s/ljTJBUHWhx3FFNUDGjozUoLui7jJj
mWfwRTNRzn7c3Tv1ixVLGJfVPac+/da+8P6uexnoFuedzuto0B7FlCbKzzvprBn9sYhibYXizxu6
e26uWqpz4kDyHmiFMrgr/JnASImud9Oz3KEdx3JtXmjLrplkhwQIM78LrD6S2EINTKrL64mt6nbM
+dy3pqdKkuZUA6s58hbO02Xp1JyAXHEBQNFGiKVLr+XVWjd7V7Qgtj85de8usOYTvs7JWpe/jGb+
QUxw3+9W13rjuB0PnHrNZXdDduPa5aNnF00KNw6aW7ednotpqAcMGKZlC2ygHS5M/OJEXMgbGU63
IiB08xrk9+l3dWcIJWHi43sDtGxP26XJjbyWe6e300O4nIm7LAWQhzO0FHYn72klFCzOwZM18BgH
t6yEvEuDmt/PIjxJA7UM+BORINEnXWlR8PMURYVR8VYWBVaTSaS6/WQ5zjbazUa6tX/z+trhRjh9
ELu6mQ8ZJsicHdgzynFolYanVC9TjeHSv2lQlJ31gjKBnVEXjQZz9yci9DesMKhdhiIiqkV5nogz
UxvvmayVAZRi2PIyVOkDSy9s3HoiChjgsiS+nOjI52QFyOvaduC/qDKhXYSFsu+ddSNXyyhmvvLK
RiA4khnrQ64FYSqgeIhB6SEMFn4BUUYvnUBlS2rnu8bHeXOKq4O8LZ2Crg8n62fbhYgRcOZ0vfaL
0bsrDoF1b87TmI0k35BuflOkmZoaZpzNsNPqF8mZsHiMT9hSz5as8BkSO+01JoOfE1n8Unqw/jm+
H5OmzzuAsJ4bn4IruJNAqTi87ZSz+glNA6RBPBkPkNCiwtwwdC8vM59ugTCuVCe6RzSdAPTpu6fZ
V/ETA27N4hIpEIE4p0xZhjx1+ig17fq5IXuS8N07UgSW0Kiad0q4s2u2fZe/eRwv1GlHJEJnFgcn
+UatRfdWV551Ew9myzG/FK+PN5CFvXN8YOyJFkmHoOWjGw+IRun3iOSRuvxJfWNo4oUIh5ACirKg
p3Z5OVaUj/r9Jd4HnCV1ObwS0T/bMsd8iX7efkzFUnoNQGomB6jFllPLWz3tlAKRHtvvI3+5ANZm
tVAy7HjCb38MqcV5i0c8/e3RosUghob6gtQums2Vh8jnJHcyFWMkAjakuFYfSfhwc3X7UVAywPQ6
GJpQ1WNDIFO/fsjebrKNa47TeJ1XT0a2mqqIPpMqQCEd77j3Ssu8rH8d9gsxiVydMySJ0M0ZVuWG
ijPH7nOKArb/hDzUoqajYEYHSap1qIrxBXut4n2dIYDXuhrznzS9IPdDjDfQnPlB7FIKaEhq/E2c
iqWHEilg5KynQxkKfnGqhA7Db5hFp4K17c1T6MO9+BvqjwIx6NjVWS9J5X9TtDubD4qrajABkTb/
P4m/B3qqnSZuY7jWKRvRDNYFZVWRDaLxW7rd4ywmYVrD9sO+CAtqcIYnLzdS2DzwPulKyGaql807
cxDtyFpLbKiDJx2pYRkGo+57a6p9YZn1v46gkKJobf27Wo173ZudRxAoK61w/EtwhkRgllpBGF43
QcR724VW9aWG8k7WqUD0d1HIVzN0XGRCZNdhkzwmM7/bRG7vzqp6fnbe+4+CmMNgLIyR8vyBDXIS
k+fj7NtJHYeC4UG+TOuZ46LnZeDd6RjX0ITsPgnj+noy6pVqo6B1d1W8F7i7dE5VHTp3K/gcyKoK
XcG0sH4oiGESSQvVYo5KO1slA8LwXtY64SAy7pHaag8SY7Vo3F5+fyxkl7tuVfVrE8WSlVMfVj5a
eYtXQqI9ibb0FnyDpl+YQbehUxc+IO+t44qmWDzPE8AOUqun4Ex/q586FLrQ48dIaNQ6GzcS6iBa
aVvMLTegCYHQsMuCIYTUahJMmJlNKHrByjnQZzBf5hMfxMvPAyyQMXV5wYEgFC0fQ6BVG6pDelpL
GtTozDYfBqdqALmxY2gHueY4gnk6SWsyW5sHY21t/x4fTiNwn65DxfqW5R5NkjK/BSXAc3MnXfdK
/BMYg0gjHMSTWcuweW8n44E6csr8iUTM6N/a5a0zbzhWvU3QAvKY+BfWGkoFBN6LTB/n2EYSP+1g
wd1/01sE6b5OYKBkF5xzLsmtNKv0K+q1nK9mC9wTRkH4zi5qh6CcI1/KasRS8MtWnuFr8Bky60gc
Sqb8Zk7UDVMNzOxPgtlHhP25BLIygrA4CC+KKnxywtRj6yddIG7cyxzlO5/44jM7aa7yfCnF5mif
/hnbWlm/Z5fXsrXxt6KDkIMIavhPWgZj7+n6m33fYYENl/DHxZY8JzaQhEDc3b+oFw/fbYZRlBCI
UwcFTwgEmSH8KSPUH1yGOPo53prHnyi+AX7K/PayenAb3sxWEnJ2rxR0aRJXBKah74Ucn1PwUcVI
M8vG9Or/v8qapDqhsZ86DkJuyv8ihbTYldJ8pG4BWThnmXlvU70piY98S5uuRLg1r9GvbqivULh6
G2WuQMa02FJzVx9mN/00DHEmruQ7GSmQkz01/V+S+EE4OCsW2tu0rYHyNF5zol3ohrlmXmvIAFa3
ojtSbRU6L7jmrTvc2nYKz9BHRHloI7L5jkRjazEtEHJLHAtSoNCYEzp/N9B+BHUxjykWplqCyS6/
1WYlsxn6/dy8hR3jz/O0jTOBXHvGMq33JEjpoLrhwkcH3HQZqUXKHOBHvK54r4+ptRJ1+bCch13e
Z3aX3LRHKF0ZdteqBM8d9NIOcU92WYK2MboVfhaNb1oLmb2hwyKtRsrngj4iKIupgihSTzaaPD7r
0qhldWb3tz+PdBVttB1LbffyDIQlWCNVFThafZPZb1Jz4iIWMSeh8dP79xq8IxyPPLOlKwqJxR4q
7PRSYcn29LJTnsKYZT+E/PKCRgut+i/kiPcbst+pzvf1P5l+rPu7t9IYzV3fYp6z2UzvOjgf6I4o
zWb4TC5dIngwt97lgZ6raN4NVbXogx5OXR7Xi+JNt5tcEu0iHxsLl6DsEeIy8FPOiE8dUVqfv6uq
T+iuBkyzJPQcgn9lRMCxaMzgU34o8L9hb05sG4qTiR9zjgRGESfkHO6gn/Dz/ofMGjWAzvR32JTV
nz+HabXIXAE6sCKhe5hWL6irLXBSka2vYMd6eUtiQUjIAn9RDq9Q0yWAdj0pg2EbgJovD8T93tx4
pGB3K+0sEDcg4pKjFMvOI/mQQypuaaRXg58qwlF/77nvR06fCCgRUQnGKqjdJmkLCTp1f2TuYzcM
TBygH6+3AxUzr1CXzNj95iq5ire7FBNwVb4NZsN7kso5fYs6RcRaa5FWppMvWGMrt+L/zVo/2cIA
Xp27y0u3NFt7KACQXIKcNYNy/q7KqSSyTyG8Qyp8JVg+yuYJFMQ73HJAunjXqp3IE0q3SBnFFWRm
rUXEttwm333VOPI5bcUwJsmzAbeIPsy7Y1iSSbUbzXSt7gCjg0BNoFNb6cs2KUsjCYzGgz285uly
nK+vuICp88mo0ssl9AN70ZfzS5VeqwQAhh29MXelXqKpZPlDYo28TGOj8d7z9SA3W22kpoCBRovF
hMkj57fF8XYKT8V3QCSwAMXjXX12UCHq2UGXWsi0quTfOXJkgj4NbOycjvEa+zzNMs1Ad8h88u7g
z/uClBOFjWeGPk5NtsltErRsoWPVZqvVBdb/eY4xvBfPwKgw/MByYrtWIZ42H8Z7hn4wXQUWP9Wv
2ZLXF/XTOoUtnGGYyPE/jdPGlEiw3+nmVXgV94vMkU+0vpJ3BEyz8EAfB+p7xr+KoknmznEs3wmR
dGfPb/KAGx5gwfrPlPW9uT4DYrNHDEDiq2HGC0IHzZYX5mAr4evcV3ZeqS8htLkNhSY7YPtO3O/j
8iWx35y1Av9p5sAQiIBZBbDk9GC7XO3AaxqEfHFhtA0UYs0zcwjOmuRcbVWJLLneLcHzvzgWXVEG
t92UeW33l48SsZDtzZ0mfobv7OoB/pQsePAzbrxHWYqMcWEmGYY7alo1ZvO3d79oLc7zy+dEDml1
jpArrEYIuhzshMgng9DsI/PbLZStakT2QdXGVQvCI0MzmQVLpH6XEcXra0R0PcCZqwclnToNmSJr
+L73TB9Quc87fbEbiD8BLojvJUMhoArU+xpFVC7pjQiF94CZ5bx3p8KnVifxqxpZVsSyIT4vkzyr
0PAFi/5JHAij31W6xUD/1H4F3fCK/0WnX+hj0LotNHM4MO6pE+0aKFryklOKJkAzzUlSAVIEc6U4
vcMZpzO6PpaTei+iLqmBtZ3spI6SZIauT5tf8PS5/FFAGwNLW3SDH0AFaRSdsboUAW19cJsWBb/P
qpd3g2cX0LH1uQL7z34daTEKnYiUYDVoQ6APrzSMMqo4njyaBW7IrnjWpY1jFmgVHe6Qma2H9WRQ
je03eBAZ89c2KqKe5mB2vKI/xO8MCXOYLWGbGlX14dJJBGprY9FIZAZpYYfjJcOIlcC3InCSBmqe
dq57JdBpQFmJk5VFKVHQEULNPyYiBdamUIvV+UVFnLd9k+kINvFtXCzl3PWqVkvTDsC2C/fbfzqh
ujrygw2SFi1QuJfUyoiecF0azLUVr0V3jFzMbrifTMEfFvm4QWW9ez84zL7hl20yFehk4Wkv02Wc
uYvmWanbpflLfvQ0QsOy8ewYG7wkFU4LupFvn6mIGpj/DDoyGp/LFuH0UDJGlhpR1uc6yQhfBLi8
Qttchpsue6FoZhXyYMK1y3xChN2ieUd/3oW+QigfOuf1QfDT/BEUI5OKfPsqRmdErL/iiuVDtsFY
g1tWYg/4qjWSHSuotL2yQZPJF9S9vJi//qeiZxg5x0WrZ6UV/RlLuqQ5vpfW4IxnaIm42HlFhww6
0CYlh2w4+lR1xgKpnk34eGKj7HesCBicmBgy6tT/oAwvRL0nSxmNb78WvCR1OPjAEdEUONZMyfnR
cFTIkBFb7kXKIDsPmn5SiWj1ycrB3/OgnFTs1Y8KvaYspT+1HCuhYzrUdQnOtVciTaSQz27KcJmV
4ZUCHRSQA/EyVxb0Uyav4SxYSpHkm4rm/oimfQFz+AjmMEeBH/hVH785zFL27pY7i0JFaPgM7jVi
LrLMc2u3+qmVV58RF6BV4dawot+I56YxBtIAsLzMoiqV2V2jl/IhQZ+pTYfiYZDhfyQzzPHeAsaX
6oI/uLy352Hj2PCxFt3CBuisAOfYnqi4cQ5i0Hq9jtzXhTaftXgRnq70/KOw6R9MF5KBQ4XwT9Rr
9zI8UJZFcyeh3o4+gdGuYbpW/ZzWax5KPJlL6KIr12MrzdqzcNWfZ5Qehryn5gw8ap4pRpu4AYjc
4wdRoR+rAry9PacULZuNiKwexwuYaXxYG2Og1dun3oiEnaOSPjvcbicDRItQM3WgQnhGU6ADL2W1
Wl38aZxvscXFIMeKz+3ZzHlmj0Xfld2/x2hMrdaviKH+Sfh1L5NABsRjVAxcMcwCT52Jo3r3SDCm
aVh71ymuJDuL7bJFeYQ/jpFn3ioY9ufZNv+ysjLtwMnC7lqkSEh1B+Mf9NZlGzgxcZknn1cDsped
u8ezK+BGznKnW37GpC15aksX0joEn4U4+JGRu6ESdkxg2QObd/urxmPO9+h37kgsywKbJqDpqGC8
fYUAJw8qdKGmJUN5zwCbKFuJEawIOrJDECF7dZ/NQYynN1o4+NhWqkz/G5SRSu/oQlaADqdHwTt2
lOz+3yeaL2zmz/4Yfox2GNr9o7W+YcSb2SFKHmviJxR+F0dsnO8eVtjNScHS7lkySJ4CHvHbS3Vc
S0vtjfZZoPq8vn5C2xp92OvivulBnFwgA+zRr6BVp2M5AElpwHAZH+b+2Kel9MQ9ifSlAR7f7YXT
LNiKruOLACG2fiwF9x8SL5yI5VtCWEZprxdVL4vkaabECBVhc7V/BjtwcX2cvHfC2QnB27KxBltm
pqACPNgImVefYLWwnn97u7fdsIeIf++ivl4/SHyV8CWN3trRtJSJQNo4Rmk58wPNIh0KwfoMZa2b
HVEoemR5X5FBLhrjo3E6SsRICLHvz6J68iyJzxnEbn+4EMjBkouYVdSOiNvylemxLCjD91D5CoKs
TFkV0BjdqMpQRi1EjbhtsX/iJVe86OqlhCX5ijEBx1roYF6BucxHerKpaAAKDwes782PVqp5a5UO
dngL5WDkbhSqmNwHsZ5DagpzIC7dumNMdXRBcCNbutjlVss+IN489nrKJIKQwVlMK4Bi4DHqafP1
aHcl2J3RWKvvItkYwuTq2sZ57QUJAWh2XnF7k2/n7MA0ZGPSIjUZDV+gPwfnXxVwMTphlbqmymgt
+7i7JZa75smybZNo+2tgjzpuyEe2bhRLaLDDkDhO0dXRXgTM1Rd+ecCMdHdWZhEJE3abdaxiQcqd
t5S4b5x/jQVdMpqB+mM0v8bgBb79WnVBQimMbOUneS95yPFve1Drc3UrqJm7vX6UvI7dw5i+ujE7
HYonSBW38cq0PhOdV9UHcJOZYJtmhkUSFbi4I+RnSO1RaOnccFkzb9PA+mG5LCGb+j0Iu0qaKNRf
Ztp6YW1Qg/VoCnFNIwCu/WGXI0TK9TRotBQpL7BSzT+sQ7ZoNWRYyK3lTwV6nfLmFSijPk8+C9Jo
anSuF2tmbdFvsbwcjqcp875e/4V8GDmBOFSrIbHlerULRqtDqZP9XIkf5oPzjLpB8MMppUJeq45q
2IfH7UngamZ5wveOeT5WHTUeLnOuCI1kp/UL0+QKN1mguP9eCoNYtDjMMwQhCO+WuKf70jBPtTO1
oI95eOumCGldk/3NgN8IUgT46UjnFLP582RTY+GEUz2zxb3nYg2g4GNbytatcW8DdYn0hUMnrEWW
PDepAUYCOh8mGQY/bFHNlnfu2nGtzU+9zEc4veiKSe6l69w+dHd9Hygx/ZzgXrS74QqAkcWDHkVc
yTkGU0h0bEp+f3Cc40ITj+etEv7a44bSmw64oaG4yXZoVKHCRvyR1kkwwWIU1UOB/EDPHVzZWJbD
aSVFDhPYVkzU4CQZEu/IE26HjW538EQupYpebf557/QN4nslhM4w1hGAFlYpBizdgNB9jX4h//zS
ORsScHXh1Ml2zxP+yHYY2S8sFNK0lHuiQSh3YvOjnUuTIZWE4SP5A/T/+OB/TscicySop7PGD0jp
Uvv7MnfCd0dsy+dijNpc1qOnKLzh7w/kwu9INrVpKsbigbZVNb4SK9bQ2+Ze0qTzjGVKsHqmETge
8bMLenI5eq2CmGLiPaCDZ4N4+cwRLf3NyjKAxQyQd7BV2vRniu2TDvPAY25FVz7B3ZB3S7TkWO82
na5osYBu4P6mX24Xk9cxSFyGhiBZVegRcJ9nIeQeuaJUkIf9ppb2uftquZp2SBYXOxN033jcBkA+
OiY3/7+mdUtTmY3iCZy5BWi8//gK5pwmFVe3n8U/H4CvIqj64PMbXJxj5Qota7HEuxbhfbhjeGFB
A0o98OEUa8mnsMmRh9/EftNvyY+PVlgxb3R7s4WV4ABzmrF2OgboN2s+aEV39fuzeWC/NIbRGQ3s
EHHz+GAxvVOEwjs7CYlLk09wlNYvNP8H3q8FiWkn2EOSQahRkfUS5WJY9HH4HK5TWQmuBvFJsJB6
8DRRkKpmqSM+ywsCADxeOrShDJNkm16KWot/yD01Ds0LuroXG0kKhS96w1QdCEaG1QtkG3/BbDm7
YZJAK8yFq50JUefch08JpjdzOqxS6Oh/iQpHGebR5upkSJZ6sMveN0+xLX0zZDlKPBWKRzJNCdgM
S45UXscR60DwQ1hPbGGZ7G9VZWZIrWtmJshob5YefC0Vn6EMMfSwr0G3x2FZ3oz/Y3q9VN7Pv/WX
rURKCx96sgMv0Pd05pOKDjFFH+F6orK4rGIS28jBnosyonG3Wpta+VpS/PLvF2otMfmk/XoVPoS4
x9oegwgk3h3itRamhrVWbLpi2Cs8HSd7+5YGQEPeEDMQ25P17Ygsh2cKsEf6hIH9PMnUIxvcJOep
8iuBnDayw+Voa77UshzT+xjpz8GPxJvouXyJgCXgiDPFQsknUNNtmuLCp7hmZWH82NuWBkHrVqL+
NKWwIxUvSEfdiJHPZyMvZzZcHHnDziLPGnzzvpTl4+tPaN+OAA+2cRYCHud3yPBBU6swqXD+5qVf
kP9XhupaPHr/9bzxKRCsJfW+mWrzNQj7D2OkOkE8Cmrzs4Es1cyTQCeecmZwaNR+ySJVLSmWlA5v
pMK+ZOhY+L4MMdFNtmIJ4MPfMFACFz+3YQvfLuwTqbie9nXwfLJ1mJnUOLtVUBzmvtiWxrrvb6WS
lAk7By7Hb39PikZhjH9yRUrRvJtDxOyi6JJVkWigddHzH9o2uyYVeZnXbloxEOWjoTCdq25o4jJU
/PvoUgCsslXYaf3tYDYe9UoqpBPiPHO1s4+l3hS0t+sxhdhzvEYOGMI3rcSnORBfDS54d5fMAU81
pPVzdJ8/2CEJSD+XlKIfCGnPj9ZjFpcRKzln9JU+9ffmR6Y6LbP7JAXt37MSiwjz6eJd4n9aF+nF
LgMaX0f02v0nEcwyJ+BAIemWErecwR1R62ZdcY5fUX+5vu8VEoiGQImQ2JK4mk4/E6wc2HVpFDey
yxTXwls2QZDM6yornqCUu/Ba48o4auFrKhdCcF1ZLIcdYr+psI/6vvCG/nrQUskCI5U8XxKZS+0O
uM4hQpoxJpVxb79Y5hhaT/VO0XhM+V8mamTZ8c7pblEKRIFJDC/e+1NRP4/kHpX+fmaM5uBtgEth
9eLqNF/auq/+u+rerbLUHkSrlxr3UCR9o/waV62/NELJFlU8pbk/VR4zlnKTEAW7mPpFuEXJccR2
kyxS74Gen45bp5W8oXXdUG7Yia6FXrcWq25cxVd3kYAU8VRj4pnN4emWvVeoYmznBB+ZQUKkeqNG
QKGYJ1amiLfKEHXizC+6nZMv3e2vmFbvRuBWH6gThYivKgijjciH7bM1GgzVocQ/jXjaqiNWhFc7
a8FJW9EHF5G/GGZhip4/zqgXVP4ASDj9ODGSBn0Ws/8BoL/4PShquEhgR4/RgafYH5D+Eqs07m6t
PfJeWfwsrtLz8tNQ1ciZVquaE9i4b+LQ6fBvuaFgjHOcsOwh0j45NsJoiuY5waiZ0Md4+/XYpv/9
2RGq47opRy2rhv3z8+uo7UfJkwDNNmQ+huOM/43lb6sWhhICKpeBpTgLsd75NsmhAwvRenHxIeJO
Bd8SZTkR9Qt8gYevsl4fFjRBqMUDQOCBiGpZNx93xh+Rjrtane46vuElVHu8mLLfvaNcWImMRfXX
rSKr0IgHXRvv2xioL8fULtcJwrjPPJFJDfltM3qwe1OyYSrMxcZB+TQFoykO+5tiqwp0926YW99K
/ycfBqgqEFOb7cBAkRcID7O7hUmyzhjHcH8KfXQq+YGiM2HOHAw5E11jVSGhSFo9Z4OS4gWWvqqH
qUxHPlMi3vAVOL9ku0DAejY42iufEnw9t/Mp7XKENCQ7/Omj63Qx7aI7PWd4ZZPNq+eJ8ExosXtG
5d9rIoDu60XMP5hDlGfKhA4w/nqb/14LLV1/gnF8KqPkj2YCBUDq7KS4/YbjIH6OaUNmDbAAU/3/
0OdXfREKhMftXtSrM36KY7iwXGD3VQ2ovCJuRepbpXYITQyJate1RoEJxlVzMsMCz2Ovkd1Wq0Bp
fzd2zTaV8ZzCK5KGtKMcp2Fuw7LbSNIS/qZg1tumf3gTmNOVt90e9/PrxZix9AK1Bv/k2RAK49DK
381aHKui0lTirYqv+pjOWeleIJN/O134uGOEXOfNi69/k2dTMU9Bs2iARzD6MEurWqAawuqgPU6k
Lyp0gVtrtE/cmJ1EG59VP9bG7jLUiok60mBJ0BqzyAt8wWZcPUYHrHZdamkAYhT1x4CIJk8X6Tmi
x0Pu3+KJFaxsA4YcPUu8pD8gmlyJ2ubpXCMbdt3vHk1pOzHmcDzFidjywobBlwdHpF7hnojHUIXF
gKDaCAsdmWP3J9YPZG53DOqptVju9BtkR9jQ0zSYRQiyOQ3EdpXyAoG958JTiinTTgU95XpaMHN3
lpavORciNkuzsPPRJ+4KHtig/tGu7PXarc691UkcjQLt1V0Wi1aqO24EBYgC+PDOetAoeUwo4Gv/
JC3r/cq5Y64Ntm+sWkDMSoUxEAtWnm0EGy/m0/WfA3JoP1Ob+W9Ixt+4bkh1dqmDzCPxhSElDCaZ
5XKGwXL5dExKj5TOqIdFeWdugUjFDCwo1kDchq6NhdnO7voj5pHeuCKJt2IzM9c0qg2R1CzEOGMp
pBXUb5aPy7BYaZhX46XOGKIrVkopeNUxLufnGZZ48cLo6uPF28dO0iwWIDsTchM57PtZfkExY4VN
DL46M71bbqF9jhV8AyytbTCE7qZEj2/k7ODKLmp8KgACoTmRUOVAt6m0oCSi7GelLN2gILQnge2o
ZmDrA3uAsazbN8FzTAmOc0p70Q/qoFeaLfgqDEilZu/LoajLZnx00eFJBElD6LRdYGAkCQqNY9WZ
wSPw6yuD8sSLP86z7RT3cxml/b+nFDKscTIYGYQgR2L3JYhgXwlxu516qfWSmV3spLZ8KFxsUZPz
BruyvqpW4J6DwK4qganZj4mOIdRm/tfEIutWE4+5WHfSyysfGD6vJV8Ixbjm1GMf1UL+Mhv5nTKY
onO8i0OY0Iue5ZN++E5EjFdLDMbdLht4osBdSikj53do99eKKoBc2NNPex7ap2VYRsiWKNyi1yFf
NZlkca+eiHuDTKD0R/g3JKq2FIAVz9HxE32xL4Ic3tU1ciljwZ/gpiNkYMFnODaziGf0RuCtDgW/
Cbv5WTmsHSHkPOqiHPseIcbod/aaHudD6eddiCzi4nCCH2SaNHMtRRTrpFQ4J8gI9U3X6PZEik8q
t2Rbn/vR2sUdRnuthBhSBNfC2AFUtuo71ZN6lTFUVqqmFvvmP/e8FE6S++r//Q8uywZkeQ3H/b9i
UjcRVvuNHXGbZpXsh5bH08P2FvPyt2WcaES/7EdgvlYEoqvLjZjGDpkh7LqvGuemyH+1f0AjUxtn
UYxl9DGiQSS6/rus/+vCFAHIfiUxTdPE1C7yotG1AUuusWYBIjUXl992JGmkqrY0aUvRxO1sV9vB
GEzDEFBm1odVDjPhs6r+MVKLSBCgioV83NpkqEwNS4Bo2P6q5wKCUI/1Y2bl9vbnUsf0m+F25C+2
S1oIN3tCHM5SnFZg6g5rVE71uDDVo0HJ1fVFAVhwXFoKric+XrR8WXPesJ3nkX063Bxwyb0E8a9i
A6I0D+kPKvDIbJddWGsh7ku29xPh/LUbu0BsObdM7yRCWxHRPWX+fsmLmHuvhtsC+Zwx+EYX+Zie
peJ1cnOgwG1+dCMsxTVDVzE4ChvOP2tdpqKXREiQeprApn22WqddnnD8q0GAdzApP5/Ofjbfbo6x
Hu1WoJXnoSD8R4itAteD8KKxGMTZQf6I/H9OTRoMJiBP2RHZM/UMC1LFcKL8Yo+MQjPVFu43vhI0
28WVbij2J0S5tw7dnr6X1beEO52I41QwT64KQ13iL61oGWBWyNO5LDi+wMgDVLzdpwwUiGHQZplt
OH1Wt/uhlpFJoURBrT94uqaTGQQl/LQYfWY4UIPij+VFwVGYTGHPfbEntcW1GgH2qDNJeQ/A8RiG
6T29zj0ahes8x5oyV83oNyA2tE2tCfycAHD3HNFCreV6HIDKTH916PBtBQGr2zX5Su4cPrlIyWjN
qsv5ULlBkmfxIKdMVzbjVM+lpagNBs23KVtfG7qgqehdrCACnlplRDA0LgMGDnSsF8PJOKUiMLZV
YOEIB7TYx7EQU6edeYWHI2fa+yEOJGT21RpGohyU0Ockyk5nR69aCVCfjLT19xvEyAqyLpZH+SpZ
YIfkGXoDN/veOY4zBhht1/hXTAvDAukK/AxnWP/kmF/wDVmiNE6ZxoHk/MWpXdkCc6TIXCs5VKO6
/R9WHKgG1hfOka4amXA5OvpoWXKpyOsfHKmsHRiSLGF1SSz5npVgGAX+UoJEQ18N+JWV5bV/I83b
pC3YTp2Qrcvbm7rSLF1e+ASzcUSPM6p3zzTGxrMuj8FH4uVr6G/zE4ZpcHlnOd+CzLgaffmZ6r0H
kKGVa5wOXn2KCkFKpAmvKLgSvP0fhSeSbYR+LX/19E3s1X4XyP7LP9sO7cXlpO+jkrF98MhbZu3c
C6NPjonPMwMogoBKWHTsW0RQw5zPjAICfb2hER6aHQyLYJtQlwd+qVnLjk3tzDVc4TcTANFJq8gT
we6fyIFM9j01bfKfujnYxu0YWcV4wTptaMrvy+cn1MqbQl6x8iswF6DwFLeSmZEYDN+vKaNB6UYx
8B/L2ZfU81JehzamxcdWyC9NyrNxOEYp4SOQNMYkAVkTZd+0CiXEw2pUZP2Xar1n5Ozf+w5TLMOI
NZZxvn+IbRHtKMgO5ggymWMH70YVZFMFBNpLUn5d3Fzj8MXzvvLSHJowkYhi7+8HvjxWXkUeBf1o
91mjk/vbwbqJeIU25EICWWIR0/HuQm2bpXdWugEv0H6CxO9p0lsoGyyLSbORk8+qCICiHgdNuXUV
IuQQD4fSKORqLfJ0Gy715ykgzCmuSEsEW+6vd8BlVM8jHfMzz86IRxF4xX/8+FHl8Cg8JKTUtemK
Hzeq+3I6add7nXwSiwlB2VExDY7IfM2r+aLI7eA8MVsKmoP8Ay1ME1aUmNlkW7zzR6SQmCm/UEXD
xd6hiQdeB6pdxVdlPqQewt8mE1oqCRMHzLaoqDCW7OR15aD2ycrFoOzgG9viwSgu8vMJQ6Fl412k
VumJW3/UeO+XcpbsXcnDpT7Jq9aQAe0Vsln5AtAWOXuqx3U3O7aEKZ+dkDL0rXqPRgSqmYqaX1NT
ltk/h3j3JnAvXTlqlj/duLqWd6MZ49pepiL5k0shpR5fK3AFANr9RxJD0V8nhX6JS46IoxUp6iUl
J43+ZonoCvWU+uC/BlUIz0GLgM2H0JpnaAcpItEGcmiOu7ZFan6svj3WXI0z2aaMdFTq2j/R8206
VoCbtTvjB3xUgOp+180jM6JCvZ8IZniFb/UWEHbcyLrqNFCsT5P/EOA51DcnWtbLQ3PMsoTTEsut
LoIhVyK3ccsE8W6Wjw25x33c00t9G/dASFIu4tLmIydJTL65/1wKJVg25jwHC5VxwsmzdKmwQCfD
dxyddqVVn9LV1ei1YyENNlblyX8KTNhEhNz1y4nZ06V0XmLifPYdb40I1YEzzJd4Ntsa4tUBCjJv
aA0BuO4Hbu6jJVyyE2j6uKWbcIhm8Fvo10X5EpWikfX406Vr2e1jbLv4+hHBk7NzK9rys5w/4hfD
yxE5MzWfWnlh7LvY04z07HtajuUESJaFfTeOsGjyBgXcbWs9G8s8l1vo/k/IPVnJ3GBz5NxzqRtH
Qcd9OewXT8krNCAYl50L0xssOX82lMxmr/WzbiAoumqk9HCLzx87D4V2NUupZUSTlejkSBCevsbj
R1aApa3/GrypYxgmhIwSYph8sEH78VshlNuxJcb6a4N1zeSRPG/qBUSnYfyTsxuqEdkVBKMyn5Ll
qD7GxvYzq3UusE7A2ZRfF0fpTLdWg7fjMPjrSDuSRZAGbVPpqJfY7kETf8R9WQeo5cln9G4k+SCu
dJT6k1DyY0AAMz1yC8va1zdLM9zSrpzGuz730Pq21cuwI0fv4c2Apd3S3f02+wDFZKDYClR9pCbZ
p2XIyV2drWVdFCQyQsvmZgBSuM3IZI518Va4bJHcURxPUqkcpqHPqPv3NFQbGrFi5xFHAudiEluU
M+lavp6PlW/+nK4D2IvhGn8Jg9+y6zJqSuIu9NnJykLN5i7I/t8u01fwZb/HSIHM485YKw7mfz3K
qcSjhLMjcV0WnGcpQxRlAGH5qwugSubjRPMicMxe08w3gKzU1aM/6yllxfy/enxdpAubkouysXHr
Dkr3Kg9P43IhYFQ6Sj22DbLkfAT9DAZP62Wq4vMRpI8RvtYzhZeEf5n+hUOet2L/clHYb2b0xL0c
s8BWwCHXj0CaPT8Fp4n+x9yr67iyXBwVCHxJRmwZLJOQJTacc7Qd8gEvMBJh5FNeUY2U7100BJ+0
9Stf/2Ff2Ww9brMCyDKndoJ9ITztj5LDxLSwZQLDxdJsX9wTDZExnRu2gK8jxKSBC32VcShjpP2J
XR86sUEYY6aOCVRj2417VXQj3NPi3mXxJYQc8PheggCKfU1OzqNBM/BG+U5fEy4AAilPMFVPStrV
nB0CYTN37/Ruxrki7RZ/jeiTFgQCZ/SE3IXSq0wMAaO722nXSp3Rs9e3+dMSrV/Gr8lakmdS0j9L
qxPdWZT7QxIaYlLYWVaFbJ3d2fVyscVq0yNMn8ZliNKkcAdVqz6VoCfoxlL3ovqRxJifbma5sB0e
hD+zppZ0Z7ELGkJVCpahEBPqUUxaV2Qz0LA5WTLWi/krGJCU89PMTwQ86Q/nRLT73t+8DLJirPF4
yMTvDR+ERA+9MK0D/CD7QWxvnnPl638RusaT/KHViKdaln6gaaQcDk3fqTbS4uWPhnopMkZlzBYR
lLcG9RybaYVbKV1mrY7++4AN92i35uGlab/HKrSiUDptlPhLamcUnBiWsjpQX4CVB45ngRM/YCSW
AYRI52n34TN1liKkzJJJxsyjORPRoBAGJZYD8iN27MUv36V+GZQZD/PdlEtJlClfZUuCRYg7zPZ6
r3joW5yDGGEAJqkEHKsxye51Vtiam0iBQA6aeuJ3vuG01LY4o2PpfHi9pWsONN3XCSnWwv0LFWVl
Ea9hjs9dDvPJadd9WarZ6nMYGFHw7MJlhot9bOFoiLqJjMFSAxIkuINFpUkIxVgv9fKM7xDy2EPz
inppIZYecZMPfxz2NhPDJLlgJOocK3z1LZvAv5E3AKJCWhcQVf62TlarnrxWJsJ8QoR9+AbrkljY
vvY0UahvCJzPJA6lXDlHllSimBRvnP2t3S8YWtuMq1PxZvALFxsZViureiGoHSDjBpgEv61taMgy
l8dGUA17clnWUGhMnZfwBOHbXpc6iPAisRBf8MURenC1U8Dv0BLqQkkp1eCJgkX+o6NRoQUiIc8w
xxONREcMpOlaUjCY2Ih9sta5vzq7aDsr9yuXKKC1Viu93Vps+I2Cd/GMbdYbvP0PceZq2MtqyNFm
8O3BFMpi2J38R3k+udqPhdyb0fhCqzluvRMoYFM4qRR8FLFweriI6rxpdo3Ah1YTO9qZr8OYJf3j
qyHqYzZg4DN1ZXhNaAqJpKqc1lTv8aEPJHa4aWWVjwfgle6WkxpueDGRY1nDQGVYl5GWhC+3q5gn
snpFp9oqyS+Otul9XUWtN2iAjlzR0XRgwVdltFikMybBg+GkQ8+gIOnp2qDQmQq7qoBeLQqKCXBa
9fanAhQoHVqGE0k6TJyQoahxiRJKUyfAw4ca1k8iqQE12OKv8L/96DR16V4XZTonXH5yU+pAUdb3
M2SsaPEQ0FoAlZWE1sIWtI2mBwi6QxzE87Ml3EbsNheu/3zbb/KADy94+j0by9KcZEnGGJ3E72h+
2C9w31KJIZQLRPFUPBAgy5orODOMy5HAy2vymz7Ykyazm65+ZdPEgkWj22jFKttR2xNt8vfjdGgh
Kt6viMpJuCOC39zii5NPeBFcbflNENviR3+ZfMy3SJASah0SJ2qWEwEf0O5LMQAda15xqTFM9bow
QPueXM0Q20hx35xwP9SXCALB/IYTCFHSUazrQ3Mml/lx89xFv5kY4SZ35+9/VxBM5Zmw0yP6N2bn
U5FTLRNxBF9viulunZ7jbTO58njcpYJag0nsQqXGNKpV8pz8hpz6pkzO3cyx08lFATOLlDFo+5BV
03pi3S3tn9wed8f20vfCTGjUcMGWWu4VXwYFNcuLGmGPc+I6ZHaqTNb+/9Yk/KTJMGDE2hoKZJdb
QVj5r667b4VplQE06IgPeU1A7giY3p5jBgRc+oL5GVt1bmIO7oaWGwIPOJsaMiPy7Rjo/TddEeTF
jnyjw7P4KTHx6I8YEDCkjcojb0ffsPmvt9vmnUW73bVn770HXCscRYLtBOBFGMwcBCQ5EL9N+iVF
3IcknfKBEyecIbklTKpG+peV4RbYgg5WlJhlxjNNFmSEcvZ9F3/O2TGbXiJUWOoiTwdIVUwntc1O
GXfoKGzdPuiHYVPmUnvHtDb/lusvBYRmEu5PiJP5uh6DA8B54wd33FgziddGkHYavTM5uWRQ9FBk
a6m51iQMjUispkTrw7Zjtx2CpShENcmXtjcKfmT3wNkJRTHeSzgrsIJuhUGvxJUeqhxvmrEQbC+v
/vzlfbAc7qw/1AhFN3CGZ7D9VOVm4KQb6AkAsWmuj2oywGTju3smeGLXoencMSupaGpyyIwHjzff
QY82VbPCaw80ljiWh5CAvqZrg50Jn5aceVjacwiMuI+SnSOrG1Ru6dBLdVLTjvXJCbpNXlJRdMpC
KYAubBeg3k7MqJyWZ3dgMGnG5YYzajW98FPgwWQDKxrJApsE1bXkI+JoRQp8uh1Nj1xbEUOMiqh6
lTJfNgm0HvHksG5jwXyQX2mJ71GoBuNYM7mBfgpO6TZaVI7AHYb3oJZBbWSFWoaa8stuP67+tzcu
lgNAbfN+aZ96oSnPRZoNfs7DuNR3TVaVeRCQIJxkVNCEPZvKRcWSUh8QUPhpmtTbuZVyfJebCzb1
OwbICNt9avUyirf2qfYHFM9cso+BrE2f5YPTxLcSZvT/mibWwYjRfJBKX2G9CF+TarYjqdp3W1xt
Hoj92citzV/1WTHIMBUWzUn+dXbOKqaDN+bGA/xD1wRZP0L4eg18rAVekSxWyC/ZknqAu2knhQL5
yjnDz0XJzB4sFFEttRJKnhxt8Wx5OUFiyzjRg1aRoyOrDgN8JJoFH7YM2pMtrvwylgQo2zfdlUhM
P1sH+tjAcOMeT8HFk/TaJbO+zKWGR7NUsRkPrh4M3nnzwv2Kv6UJDW1ET0zrDrCVxnV1DdITi0ER
HZbzfVf/W4H7XALwCOfRcIbxX8rM0wVa2zTx0Ackr7mvJ6RDmVAqJROSlsf7mJ9C4QK9DRt6p4BE
eq7rCTYoEs+J1uMItaM1lt43CIGrI5IHoxstZ/8Ks1XTkD+GWZcroSmFd2HUbRGMSVQb0785JHYy
f5ZGrduXDSWsfPui/CiQPEE5c3hBgJfy7Ud9yDyiY4wAsty4nsodPOfxijyFU8G5f4V3IH157zon
8DsxHFvjQpyQhAFOTIwHt1IKqKNM6a/UFRp3Une0qD3zS0kK+DyVRkhol4I0YE3DeygPXZpfIPWg
yZD3HbDI9HJ3Ve+YeOvWtk+FwgT6TBru9XbSM/YyG8ywhhVEhDntDe75X0z4jFckQKqW67n6vLr3
zTPzYaatFYapbU0+ld/Y2uLXVSrXtenlwP02qiTdbGga9JIAXSK/hBK/gWuvXn8NfZiBocZmHXfH
aFgZYWLKoC9ThHY5CnRwCp+zdG22q2KlDasfuN2cETD5cwTLSZIQkhdR/CZUubeIxNm6nw0+ETHQ
O+k5XYkzQW7r8SoKhf/CIiYeQ8Br/kzuggovn8tPW8+o5C8aZhm5DgD7OpvxnN43+6EJx5507Q/d
5h0IXNyOZBDYbv+IJCy4hRrytU3k3ylNaMhNBoqZZIWeDu9gu5xGKgedbqEAYYcF5CsuTK1rAEO5
2TmQiIHeEWjSpE9p2+o67T0gDp2H1GDZUjagn0D2L9Pxhp6iSI6Q25rWv8UwAt4rU8utMteBmuyp
Pc+rPr0cUkRanxZEfn93KOqESKIUKAkghNPxxw9NruUOzdaDA2Lxj8CBx+UnkiuH57E0dlQsuNpY
4ZyX26S1dhBPRlLDV04yiV//lWCnKwh7k/d6yBPQH2KFl4oz2oG8g6unaoy5WtW+kat4uE4uv/0b
64jaBNdEA9iHSYRhQ8xYV+iXII747/u//LSPLQmRGmOs4ZGKzmTAbezFoKWV7y3Avch8yxIngYXT
ZgLIcSuGuEToBEBvz6n8dJXgI/rn5k03w3ElB8dzhu6QOnYmevdmDf1aT3O7Tzf5Hnut1LlKaObJ
aso3NUItykcqy4iKOm/xrlvn2l8UlyF8uYjE8HcIxpLRAGhUaceGrXpQEnFwOjQN+YYusgKLnv3Q
Awuc+xt5NmQZACD+bgr9clUSmIUZdOw/ip/K8Uvzs31M9f4jJDmyNWHyCIh81sWokrHXmndcd3X6
PMflTRg58YBdqvCtO6UtkVkVGDhV+a2JX7cs71+hLVTbfu87QhPdjzZcpFbI2R/XX3bZMWMAnEai
lClGb/euuNHNtHT9/6phyOuzZ2YelROmDjwtGCJoM5npQewKRC798lVQdyrKaZzjwU+IKMrFvzy0
9IyD+O5ktH5AZBdWV5BnH17PtoxRc56Xp5/OB5xObybeP+RE/6Mm3ofI3NFjRiGUitqJjmMruC8O
SvxZgEyHK+ZUgMQ60IbfiibBqn/mFgrlsqml0w3gMUwxZu/F5Lev2ZK5hCHS+ugv1enSY6Tgev12
nMZfGyBcjRuulU3qHMdbC2sJ6/4vAjmOwLa/S9ki0wemdmdso+BKrxU7ZJabviqwotNUMW7Y3v1i
JMl1IrpCbqCmBhv4JIDJaGi/ONXobm9ReRYD5O0J85tbQremSCUaYFjp0p+iHd90bKbk7lMs7dDp
Wu1OsPyoXhDRN1axTS3i2yNDZr1IBNlg2UnJ/WFq08YIT3kSsVvm5qDu/z+efGbc2uktdbQwjQGE
hYBb+tHmLVkAvrrrYlREsvNJYWMJ5tScAvTUfNBcQDTEo0rzK1TcJcqGBwpldU3bn2oo3b7uVq7U
7ibhg6dk9FGWvM37P/v8unxZi9kMfX/Ph57C3bon79oGbcj6YZzicCb0sdm/cPbOIlqVeAZyuIZv
t43VtQcmXta/dKSKlDUKGqxt5XJDUO1VrzfOArJpC/0oduW43gmiffbPRsL0PKTxsjr+6GOPKTRH
374unYmLIx6j/o+jLab85/Wzia4f/aoUhLQt6Y4mpZ5P3eUXS3uDiqjezPx8GN6uIj0+FEumUgS1
f7uAOw7pBV0fahJkvdvUyUE8YR3KxQ95TGnj+KSyQAQYoagwW4vTpa/WHDHIvcpPgcnw9LPk2rgf
LpS43amSJNLUUlfDondsJCZnJYQ8XiLvwlvEwD9TJmIv46utq0AY2+0Id+NcBON1+dCeGFgrtm0O
bpEgfBLsbZiMnFW70v+hRzlFaXsnJ0Wngp3E5ZRbo6R5W3DUaRfFqZz6Ge4MgEQBcyvao0LktqGP
2BqBa/3nUXL9GTEnTorEaHziyIx4OVOh5AHsVUxpHmCeeuD58GVwWFgp1pxtUjhuHLsEbY+yn+j6
JYFL8UIvs9ZJEa00Wj7T0xineOxVliPH8Pg1ciVjHL7lXOyIyasPBMLT0DYzZJUPLiteJAg7Br5C
fXddifsstK/L+D3OkqJlOBoUSeAUAZn4V4MXHkGmt4YHsu3cXsJHLs2xmCIeuLnYNe5EBlvh2cd5
ukE3boWH/icgrwM/wftDY9FbG/lS5fw4VCnD5ve7Un4Tn5pC0hgStTc71lUcvMy/VHrQPv7eyz1E
5eHHVcZLXsmdD0OYL7hp+NM8ErOcv7GOOBRCCfgWaezeRxyyBb3e+ZrssBcnKzaxAUCt7dVU4xS8
8MzDNtYU5gM7GfcWxJ3viWxpOi+3kymfAj+lxNP8U5/HkfdS4E48ZlhMncaEXNB5GgxhvZ/Ad0SC
00vNmJbyn7qoPnWdkRzPiNFetxDC3WrXLyMVPWFfSnBuADZGc5joXHRStpIH8Vsz3q5FuTSo+TI3
t8Fj8oplne+xvGRMyQ3rA9EBvOKJD79h9XVyPTrKb7ExzoX/d0uQVj3pCVrZ1KWZ6L8FeUGGCk/K
PdpL1AhC7SEF3Jqsa0oMK0IsNmRmdzTz3gpY9VbKxQjkCmYE5vaMFoQGpZlYvpQX1Cdav0iDDZXw
71aql0AXjQQVN1ck9J9j5SBgQ4idlrkCClWV8vZvd4d6ZCt/SDZAY8qekQfINrR8bv1o+oC87fBF
qxMy6mqw3pX8a38s6/zeOsLVFpG+k/BvAZ2KK3TezeB4CEKOCN34bTPvJtOPZSr2TAPBu6SpvrAY
kx4Rg7l9dR5N9drJDF90duIx8FXTZpm7QAs16E7TREtSu+6W4GUHagWBuFpFTbA8ZYaEzfE6fNrq
9ZfvpQFRm7Av5eh1w4n+6CncAQe0MPPP+nMPZTBwxmA1p86OCzW+bJgLLaPjbhIptZRFUjzp39qp
82hMk6PDrGe7giyBto+x+CNdIjmqCpyt0rHyztIDrOpLI9pIkIF0OYD74BeIkECXr2FLZCGYg5rl
Mgob2KqdJuUyiTmdcWr1b+7sbgVboYgZRWh0scCcxgsXV3GOotPur42DPYJPe/huU6E9M3kABz7F
Es5zGUVnkdbobN1duxs8ZswANRxAZOya+zFRo+XNaw7GWORU9h4GAlaDJRFX36+kJm0+gP9Heya+
42cJ8PTYfh6XTorM+adqMRdZzcfaY1pDJX6mwNy4ECtRH+Yi1ocPWmbXS3MrO0lhJtHH7s/NoYIT
+aoBnry1W2A3ebTvLEI3P92xjtijRxaCmaIfY3aQRLjIwH+fFrpmft/Mzp1u3vExHCIp/GJ/sTmx
/YoyvW9y3geiRStZ2Y1o08FVgeA5pxXjpByVo/ksI2bCBkDSva7++ttLxLGiZ5R3ACBzrRE3L2kw
JZpaJcGqPC2N6kE1avQ4KBfQG3uhPh9EqRZS/0fiudXgSEy+Jg5f1ZWCbR9aLW6KrynH9DZqiyTa
6/WkzOxDpBGKJE+2xwYqcOcbV07JUVbSC65+MZn3KCw9kWk+3l26fGVbbUnP2K4fD1VJIQXP99Tx
EGZxDTZSDeAL2QWywYcM3ekA3xd9pYRF2lqzvhzDp1N7k1OUrGz3ThT7fYdXSJI6is+6w+kycamA
N4vJ7AJbNu0kp3uO0MbaEpHhnr4ll5azsIT4QvdWlpWmnBmljrgWmh6vzrFRBzdcyznAeh4WmQLx
2J+Ek1WrLRCfI3h9gsrfmqmFhb6xjb62DRNrsZcHMDGNUG3/RNd98AuHcE2kxN/XODGoI1gM3SSs
7ut/C4HW5dxT+2XE0jmmXHm0LcOswx44QK8GZp3+CHHWTxIjj2mnKbs8KtsrqchpW2Qw0pWLcYb+
iRowPu/j3PPjGT7sXEg2v8mm2zjy56v1e2sp+tuN6gdqmIQhiFwRnf5I00hj5SoZFWJGDFA+qu1b
bl81mRusU75rPYZMlnggNFR3K5piFCRly5RyBl4r7lTpNPtDJ2O4lF1YlLlMv42iOe6EPUUn4G+w
ssaV8rbiMTV6Kk4GUgEdwAS7UFy65LtTn9YtTDIwYB3ox7JTlM8XY3QEOevc3TcPJcId/J/LmGZC
x1/sYHSSMKenfEaDJa8cLYaNu+fuRxmeNJNZf3CuDMHADdXUGhgIk/VlTKTNhiI/3R/PYy3sda9V
BXfyvaXzC7KA/G6SglR8FuZgvPHEWxPqmSuVBd6gxGgeldXLhWEWfC5joWl2zT5BvKoRY4dXWVOe
LyBNHZQOvZbzx5oYHaBTU7QyXV4qRc5h/E6lzd5IaoXopclwQV+fPdEumVUwhIP+o12y2XECA1Ln
+l2O5j4XlihJPlJeBJchUPbsqY4GnKoa8J8AtxFXIpMGsfKlhBwC855HQkxUpBTJIM4gyb8vKrFA
zUbFFGZn2GIWYTP55V23qJp8Nxx22DU5QUxRFkFukd8OAjpI6p5QYWDy5NjcW7eWmCUKicCFPku+
w/pogtjxsT2cjvC4MPLkenQNvGVD6ULsVphMp33nq1VDguITfjSruFVc8KV2WvAqnWzeBM7oaT9l
kBGYTgkH4l4l7zdKf6mBMG50WP+H1ieGLSrHQE3JhZ4cuEH2tMmCpDokUs0aIsJdpmQij8OuPY43
0U8GRGkN3snU1Eb9qKnPR9bRgvhHzAFkflelKpYY2iNRoJTx+2LrRuod533g8uuJWZ/TucFfvj3I
Gsh52pPHIsNTVB/XbjUU2GEQf2/QCyqRjkNVlyX/69awoBhQRK2qbKvBPTvu9UX0vtLA7m5cp2+M
9KftRG8fhiROw3RokCEu9AKmMgYwh2gAQkIicIcSWtYJr0WbOJopAXzb8WMleswirQ2VP9yv1kS6
ktTPB0IwkqZNNd8nVkVlhX4+M2iHqr4xyyBuDNd7ln9xPbzLO080k5hhhpd50ltaHdC99Mg/roAF
VhfrYc+isCwUmdBW2NaWCCmRnOFHMfh1w6wkGuVJmESsTAOjDznHFr3ahFmlT7sMO7Er8qtcdeZ7
Mch3C92g5xYvQ2TJMJLf+gjLlMl4carNMnfLY8duiXGf0ePFKnhYqpDJrzOB9eST1cNwNzNSKHzL
vmndOHJ+NBCAD1G049omgGy24lIu1/pFoSmD8tmVIxdcfzuPObV6rC3HL57RfD4xCpB0UYLj0tnh
B7bNSGcLveviJtrljsuzd0nRkNyH/9Q/IeIBx3LLHhKJiaZWeGn6z36dPdbqOhcif3jt9V4DDbTY
EKTnBZhDiOHKpDRCddOltiFBzHh/CPCwTBiuPR24hxZqVwlNIiR+wlfvXP94vLbULsyMh6H8Maew
7XZXzO6Tcp60v/GNrd5+gQ1TPtQ2MRWeTlFIdsAUepLeVuoTY3KkTE5/ustrDDxuX5+EcOyniks0
ubLYV8WMmd2az2k4671O0DAdpSgOat6hgJYQvzmqeB9ibRD/eJYjwmfEmFP59jobzgtipR7OHoUK
rig7l5636uPZB05XnIAQY7XNfGbej2+FbzBRTBUuICDbCAFSUpOB1NT2vs1d8vTJxW2J/64c0ls/
MW/8q2NAC97Y9MSMr6oEZ/XbCsQee62GyZK35islZ8jJU8la1qH8c0iWGSuDNTmrHb9IxG5Dy+pG
0VtYU6vUDIyb/8TaeNze/cb/VdxBoOONC4cHzLQqVFlBmoP7yM4o0lew1tiBjcYPQbvItQjJbbHb
UlJpuIzULt+EQGCME4/IOFi9M0EZi1m0E2nMHLt92CXfcRKPIlZE0FJ7KCTQmTIVi94V2s+PKEt3
pM1DfcQDwzRYwsJzYs8PN0c48837gH0wbNBDrU+SSerif567D6Qgi/Bu60mDJp2IoOqQB23gUCaW
e6bef6avX6MRxo+8kT/bJVFnmoO6+HyPWuZdrcf+Mc7q1PtSV1CItBg3YSg+aC7CYN+gARab+NHo
LBCk4dzyOxwonvpL670hubtAumFdImyIi0pfLqwNr7RoxIiTnCzDj9sHGo2g+DUg8FiId2dc9Lmd
xa7zcXQyj2RS3tIZhFWVuekjuRFUXBzu++9YB2YhgC+Ec75rrQokD0r5HO+zEyo/hluMhXLdomUn
hvxOHDEq94nfbWFrLTujNddaPuac1ymU6ZQmDMU+4JzzqTXezkqVp0huI+o631ESUjFyIgqhuzJa
GuPe5yKt9aaJdz4e9p4v5aNFvm5a5AHPfu2Ri/W8d4nRTA7OVHF30+dQnRTpodcfK828a85qznKo
rrS4oRSp2+7ETbP7pGknlGIa+CFswMQMST5N6h47X8TOqfU1VmklKMcV+3UDCsEHtMmoIhGuONLO
MHGd3xx4ZAtymQSkXtslxHiBuimRZDbkcYi7Lz7Fr58QWZoiHcrkX0wO4JLLxUvJ6sS7IcM11YcN
61saTeNcdrEvTFkhq8RGenxLjMBleU9hJRA/XvoaLx1kaMdl+NkAXXLd79n54LG1cWYALdp8cytp
4QD7ELX8L+h97wmv+kBzwiLB6BiyHl16th4O3mjijWA3CUHb2EhVRHxsvsyPFTTdHDufebr+j5+m
XWCXE/K+KAJVJm93ZV0NC97vnXszRdnseQG/JVErDzpaC0G1LZEm66zzlTUw0wyCzGtLqoHBOiwI
iX+hcf8HYNAWV2XBN+8N2SyxcBmtlXy7dj9+5K2ESmF2l5crIelPU8BPYMyYPRLv9xWQpDEXkmlQ
CgggVl68W2hmSpLy84RUxPvfqlM2xBRI9jUv+NOtu+xnrtbp7fhzu62434Oxq4pV/WArI1kXVJ9T
oA3rKkbQMTKLDTnRWr41tL34dUYkJv0xA9k2UJr2Dm4eikFKbFd5Pd6JYdABe5jageyW8/n4CmN1
64p5ZZQdIF4+pcFxeTwfFCUme0oqqLL4t1KRDWA2u4fvZ0F7NxFnSuVQwdL/a/ERoxUqV0pYBluy
b3v+0gldOPQXPYFFPfPQccMg5rEg3uvvX5GgcCpIO48D81Fn5DK7EUKdQ9hyk2dzpCWezy2NyWnD
QJ/UZfmoFeoxB8v4ytMcv8sxkkCgWxj9ECexFHhLIeB6akw77UnHoQtOXOi8gq6H9KoLhMj77JX3
HfeQulkyFOfKvc3xyVr7vBSvPaMxfiGlmGgQdgntJi0GovRSE2RoqITBo+BxWMYIfnlGQ/ZECyN/
xI4lp8XtJSYAhnq2/ym6WcRWYHzP7NitMDs1eZ9C1bPRazROB3qBgUMPsMkH5phYacTquNv/JVG4
41mX8imc0bHw6z/HeRR42bRwFiuaOsNq1TXh8E5UUBNaiVCKrx0jmJ0ub8iQbcdSrcS/EEmXcAnY
y6S4YIlWLNwAMwmvnrn9krc5QieHnVQRNvycOZxOD5pxxiisUKMI7ZvdE8tQGUqgGsv8JGOXsFWJ
MmRNk69yWI6V+ld7Y/nJXrNMpPehAvsphhl2aA0SEhUdzL2S6wW5GRgss2oYgcU9dQ/aW6XUe5Jc
+YqVwab/kuzPHh2qtbNstFrgpe94GLPn6P4lhZRJMrcPaTVgnGKEdJFEMc2eVdloUMiNC9leI6tL
mUKQmsUjmk9GpRQ7tk5lSzSKJIImSWHMRhk8gr+SJY5/f2oYWFHoXJT5hXfWWzAnyFuHAzv9+m/p
O9rZQcyGL9pTGeCT3Elj2Zg8IcPCYLT3tgtgQhj0jQ4NNUqfDycqbx5lST3rLYGSJe8AYTHSBVcr
cIWbM5xmJgKAgqdzKMTux+CSoRn9zejhXYb8lwrfR3A2jEwbYYvvhk6cYMUmc2jTPG2MtaNlvPEQ
DwTec5MzOB2uJH2qtQbXfFb/nbY2X/Q9OlG1xtZPInFsKlcXR1aRsBFrmOc6tjVWuF6El4QIFpXC
r0C6SdBa8rBX8fDU7CdoAVPk81aHWC0cdp2vfQZ9iafNMF7Tbx33jVIx6nbQG1PUFKT4cTjLCeny
MVinTwSQlrAvPjDbB8yTEv1mUh7QqvEA7ermu/dvQw/MrQTXMhYz2tGzsulcecHNFgZkdyh+U7YR
uN7RIqZOSrjtlX7JAJeMWa09yZM1BOAfIRWkVUFlfQBty6eHmvKm3WSMDNoaYdLOby9idOJau90H
CUauC6mqLwcgUt11kQqDySmyuEIbtwQ6mNkvTPHlnLVkIHLHJkv5MXeZptfo9mcADa9D7Ikq1J45
25JMqCtKl7cManjtWDTKotD6GN7sm0vfObC0Mta4HhUcfrDye6u0SoqAzQQIG1SALqIs7fVHFxox
F4J2FA3qLgfn21rsTL6zvN9TGQfkglIoTrEyFAijeDjRALDdBUqlyKr54dApvwcTtYjmeCkYq3Tp
7780nuDGhI/L/ZiTWPq7TXlHsUydiwbqoJN1hHlxOvFQHROSEPYzCBhUULYgS1XrShHY0oPWOKWU
egdeQ3Sf3/RGYn6bD5P6PsJ5cOw7cmmhzMOBFXFwaiIS0h4gWTPtdR89RdnFCFy5copOxIANe9zb
i1bD/XakDcLw+1StVK1ddbm5oqg+PoeFxreyzv+v/XxpxnGmqEC/Wadx5KH33CAZz8mAHtsgQWji
2Ob5DFhI6r1sc8pL6v2wIccDzwMvO+v2+y5OQEoRPCQ5ap/CoNv593KSwPdPHpS+LJDtwqyZfc3I
u+85L9Loi9drk/76efKj62pGylgY9cqIzEDHEEaNb3iTytPL3XW2GTzQ2wshoNIaMEWgjg2nMyYh
UV+rNDzDjy8KW7jOM+NGuEorgK05ECSsYjYXrTtrf8HOGLjND3vKrJt36S4t+xeVjm1OR6XGnOYp
wdRq/Mu4iWYGZkUSrXsjOe9nZcrVo0eoBRcsvl8KtPwWiR5sJ6qVqiIVPa+NWVBZJ44a65FAUm4L
UcgCl1oc6sLmoXl+lk4+W4mlG9AZAh/15pgAu7iM13aWB2F/gqxQRheLGvDLy5iUVO+vorlW8XQ8
B4RUf3TZiMvXuBs8I2ahfcJMVG0v/LkoLzq3n7PYtFg2wolyE9FOGylmVnWztF6tQE2EFfqDCzm8
uyH5nfRukm8H4kdTtTy+Ah+tTUR1LOzhDi7FfZwKVThSG41xnL4ymWeEjxQXpADiJFpXPtJNcD8Y
n4uJOgnI2SHcgGmzGWcxV7uy2KCz0mAXcyq+ACOFGcb+vRgNCIzYDQ4fzwuPoPbHyv3hv6TK8I3Y
DWCfliusdggJA6NUJVto84EAIchAGwwl2ipuEi92JJXXmxPIiGaHKoj78uDX4GXbImFH9z0nNRnQ
ucvxHH/0dvBCEk1D3XmAfUkUYROEIXwaouHPHBHY1zLuukkFBqwE8sWlg0DRFzJbJJRj6KI30oOA
GHeakoRiaftfx2bhMpNNNB2L7yQIfo4J6EVo4xmgZyRl/TQJOJESFUK2tdq7k+qIS/cHioZoaZnK
7ODvAeF8T6BPSDidE136+T5rrYO0iVaQn+UMLFIKrURmfvdVtq7GQMkW1yVad0hDHtp6RSs1M9uM
erBRPpmTRhebLNkNrJQQgnur3/RFwQjTMeN8+ki5WRaVOCviSUWYVNGyNXlpk7OzoxM6bQAtD23n
PUlSsPiSGbVSNz2/LFdYXssRuGDVTIrZC4s2rjJihstv6BZawlecQRwjPkSbhtq3GKbAhNwPZGzR
QVCPOgBRmYUGN9Gi5wVb9LIDgxKVT9WvWeJDfzuZ1sjZfi64qyEOwaEKL2Nba4oo9p5t0PYhf+22
2NRYFYhaB7nfP7W1JRa4QMWGcF4FaU5PL0FuSp3qKiRePI5tsnaTYMqFWz9lPrdGWEzbkzGfE/wE
GCbsPofrrVarLwur3T1P4hEqmxp/fe68TPnB0RT426ezgwX7sUi4jrdOYzIzttRjQupCMoidm85P
qercZXV44TEv2vo6uraWXecgRPVaZbA97t/UbZykHRXBnEwt6ShvUBHKx/u45L4OKJpTetNnpD4O
/+c7G7UcD43j4Nzrd5sHLcyJEEKgFf3ny7PprckZWZiY0JeZ2MEXyxD57Snd4U5fIDpWDau6dv57
J4KE/L9TUrySzWbcJUmbmRanZ+sZ6Qd4pR6oE42HLi7LFd0ufabbku4xQVCDhxwVOQPoBbhRlVXQ
Roc4x2sEYXm2rdVPsWcfbyghDqE6rp/pzFkfW68GAZwuNPQ2pCdha/k41RjozMeJpbCtXyxy0mjJ
zcdGMcbMeR83hzkwDdKjwbpJPWDJVeLkNC5sducRDL4XI2Rytqripe9TOTujS9Jwb4bA00aVUtZ7
WzwDeX9q3MVsuwyUrfpxAlNUGLJfc4qcUbmVubnsPvO/4+JQ4IT7uEtiCO4T2Je9epmzk+sPCTLD
B5GcIs33ZU087mTADSyW5Js9AD3YWucpY6qhTc3BekSgNL+Jd0Libkl/tVvU37vZo5G746JneCXa
CvgsRjG5huQveTYRcKkkn4CtGVBM8xrmkoKyX4s0I4pO0i/3z3DIMFtrCwZwAX75p6pQoDRlf69l
13dS8rp1FrKWUoex5Q4T6btiRp097RqKbdI+tNXeUcsCXohHGAugP/tfQB95JtXpI7lJU7EUMGDL
JvFdUyxCPcaYLpjapEU19+eoVyk1v900hOusYlKt+bvxPHONpGW9bW58nc/cAmgMtaRYtXwVx4Kw
eu3DdbuikNhNBBb37aV/4MN+GNGTH037VaNeyQw0pvuUqLZxA6AnTFLDfRzTopXE1pUmwq/KHnkq
04+jL60IP9t3mEUcKRrEFxEvJMZTj8k8inN8BdFnio5jWvEUHG5LHJ6M0plZgcrUldKzZA6gq1wJ
w1vOOcHugHxfgQzkKusaRHriyGRMycHCk9yGAwRjDvxaNfEKu+wavpmgquFC9+LtrApD63nkLLHT
qHGhvNx28qbdkjFlWcMEDBXGPzbHi6BJrhyQ25dTdcYo8RXgrKqg0EWXtei6o0xxW7Rtbw+DIMlj
ZxDnBmZVQDClOxqGh5Q8vueM1vkxtUrkNwhmogc7oItqFiBv1YYgIL8qRbYonKSZlnh6/Q2jnB7L
X9LIxTUAvlU+Sy2jv9JrwZCXp2HmI+/qW4dpNUkuVAcJFYNZMnYII4SsJWj7Yu3CDQYK2DGAbDWk
/FEtN+f3NR/XYP93vYDdyjASxmjGuuBz1M57T1LurWskPuPEIpoGcrpN+QMmWxgBD1QEMq5mJERW
eFrtokVGXI/gwBKAlZ/xMvfKQUdrpZxSNatbQ17COyjCX/N3DJ4aX2jeMOzmiIEGBZIFEd+1wZUN
RFMtyo0rPuQKIsJ9uOxw5H92WXk2krbi/hTqRdN31j62cHaJ4sfgqZqS411bkyv5IJvgOtyNMNh+
gz89JQ0qA1On+YDqH/+M48hm38+8Xoq/41ZAeDMbInWPhtrEPIHd+q1wGB+5lDYNNRGM52jFEjlR
ay2emrCoxd3N1tqWXKD9sSazbwHPDxOGHx4UqRpgKqU9V7kdE3qHgwX/D4dVgvfC9sz8F1SAL1Yl
S0X9/jrU40nDhCIM3PqBqcJw6qb30gr1cq+JZy72gHnQd5cDRzmGnWZUVckXznzMr0+6ukU8ZwLy
Z/DNmJjQYmu9TdpuynzayEMsmjmqUY2Ge81FV0wTMMHuE/Q5ZiTOv8gwUdbI8UplAmZnR+xfnDYc
GLs/oYqjv7EKeavdNyVFgNSWkSVTCq+bpF6mSwi05tI4JGbIywB7xh4LQ005kHL2RRtdu3xrhgnj
1uEUx+8TSbpSkEZNlYOtKs6vpAarut8VANf5uRvtay9w3fUpaULMZ3XuM8rJeuzzb3tAWEsGUaBR
6OGwas6m+9x3Tmn3xmLwGc3s0E0fPaB+0TSJlPUMpOkf65s1SCwm0IkOfpKaQsU6Oy2tsWLdD5aY
uIW9R4jtzj6zg4B9d6D7P+yTjJr2qbhcROiKJN7tLg6yPDXYUDLNMXddJS8H0MtUOapzQddmu1rl
+4ViMVW/KHARpzyGH0BHIZ5H+sNKnyHs2A2dnTQALHl147vDTd0PeqFjR3j40cSpCZquVGhIj0Sn
q4IMotPqhjaQHp4fguqIEX505uiCVu16BDQnQpbV2ZHdtbAFMCqOGJPvZ7Y9/J8iF2ijBeuIbbA1
N2DhHCzNX2QIoHc3r6y57/mklDS7jS9Us4CbKkT7yvhe5UxVC3Z05+40OmHuvnR16zZZV+EkJ9WV
eP1JslZWQM/xGgmrdgoqQMimDtVzejJa/Kwqq9nUM8RNYX8fSM0F78mt7HHnzvV0QWN1xBJ7faNT
AJ7ZlHT5zAX3ZJhzRWrxpdghctPgXDNFIAz++7xuV0BcGOfOGPlR0VCRuUcisz4Ws40sqCTJ9ACj
PuO+ZghXE06eXUHVC2QI5RUn5BBkQ+XLLDGwpVBY3zRPZi1CPWdhm/UKMJpCrBisN7PZ6ii/mMYJ
8WX7miYNi5Mf/PkJl3y6JAqB5CgyXzgjpM00+DLXqZPZHhKztMvqZfwiEqdmChtSKaR8PiIrMfMs
qLhq4jiR9TNdoiDjhZn80pxEtHZ0WDzjxPSmqsiHKtmsbUJNDdKRr76/HBt37401W7C9Yit+BMkR
fyUVOH3I5q+/Yh/5tgqxjyNUyUS2ci2lc6geTa+boXYhYu+jKQSZAsQIca99v2JC1/yyilmMAwCH
dteS9RyTtEjP4mlaPMbYMezhBttOmR1kxUO+d+PRIcwW9JSfRtCte9j5VRs450NJh69MFBHsoeb7
+gwpVvneNeoEPo9+62o/SaKOGUyT74YteOD6tf8qcOQJPKdZ3WXuSW8Kn4uJHjOJpX/BolxzgboW
FP0LbCLg1AiUuteWkGLSWP92Q7ShjmJCe9nfim0gLdW9kkKcPMeo19fF96ViHH6kTzvI52lqLNxL
6ZA5tMsTwTPnjgbPdjWQpKX2He+dRq0/h1sXtajD/jyBLPem0eFIH632pnWn2gkUg7s+jzeNFuYY
P3yGZK4sB1tDt/ftBA36P4Dz+cwThx9ZsKJ30S+wk6cy9aaZU1MjvQ8kXOhiL7sabRusUP1JiRxq
mYh3RKZ7k+zmMHFTq3GysMk7LE0wwLsj7jBD7iUBMlOYY8umWWDId0MPB69SdSxgp8UF5x//dDCM
aNR1SRl2kFeyKaZWOc3vmP8O3c9ELE5LhUmt5XxTFUFqBiw2VSyn2EFPEPMFVV8KNeYk6TEFioW1
DOuIAeNZrHrwwjx+gdKsxJ1OwXDdpy7bGYxIX94+xxTjV0aaRXWqtDP7SO775/hB5XazKSQMSTip
IN+U5ecRo8440TpBV6il9Kv3PXLJNBz3DY+aexUlybjK2QKGag8mfJH7WYLP63MZvxIynrF9XQj7
kzyhM/0f4ugbpiQ4KiOjwMfIp3b4tnTvc6IsGE/G+dA4yD5KzpcP1KGgJRBSyHbXYYf14liBR9z4
icbxxTfbasblNZMAcmlidzhfQ/suXfpmT4oObGw+LR4NVfNolTZAHfRGmyPWLzzUOLKs173v1rva
fVk061euRnj1SNNpgi3CE89HS112YXS22v6Vfz0zTjKbSEv534/KNCcJ7FgTakc5lx8vSLzHGcsw
MWPoVxwqw24GKhYQJlLvJQTV7EWObMQ5KXCpKAMu6GIsBHvtKvpSBnmlHYLXuKyrgWXQ5TrA6TaV
PKoorxYYDnnBV/10Wx6vyN6RCcb3nLYj7TP2VQsENZT72c8CTGU2KvqyTkVpIdSznlyd4AM8jXh5
pBaGayFw2TlMMzH8eGgPRoPV14GqXBuRqDnMiJOO7AEw/M3sVMgM5XTVzayfQlcmgvn98SB1XKsA
H4lIbE3BUMuaaCzl7fCpIs2hzP6K5f3ZZY9lXMIitl0HqNpA0f58Jv0/JN0kT1ktsR54hsLMdBc/
mF7fR5TeuA0HkH38OEl1hVwxRM6Ij7lL60Jwhh5+RqzY9+jgEoTFVYWf9Gz/shsbZ+VipPnFtB73
vCpyab9plQJ+6IDNna/MCziG6Q7Gxh9JP43Gq2nFywnlnhUj8kLT1VJJs8h8aIw/sofxKF7R/b80
zZfNRKlTS0eHzViDUN0FR2F6og76Gqe9Kg00mb7XPZx+61pr3Pbi/zQo5BXp2OIvRcWqT9W3MvXc
DPK10qCuFhzBQ7Im9xTq9vrBAGDZ5F8qaD+kpazNBpVOY8M/PmC+O1nNiTZ9BYM8f6X6ng/5lALt
pqgXmftjHGdAe3ZEofUPkaVtBb93a+dHDHNarMgTldl8cC+dfhen1Sf5I/jKMxir7Qkhfp3ROMYS
aBEQ1EQ1zX3D8GGERtViuJWq3QJ5CwmQp3NS+Elsy5NeddCrcDgSS3NiAocZEAeAp+RySr7u6PtG
qoZ7nHQyQbbcKzwKUFzOzOmu/Btwrl3eMpXlmdxzdLsE0pVBILyDU0n5RGFLpZJLfbNKn85JThPE
1w+MEUgo71fBdAZMXEoNLkkPT/p2ndeFfxGGg3z/xcA7fGFTyWFxNnfQkvbtH9lIju+C55gOlXHZ
QCpdrC6kVyjhPQuOpiZ18hcVUuo2/tD7a95SStUwE+iS8mvHF4011D/3gDQoIbWLhd4qtEYyG5Nm
6882jw15fjTvHkq7dKZj/XjcFpQpTk9lz9tpG7jlpdbpiPEGEUO6V6ETiyon9xexuh6OFPLopmFz
4n4IksGNfBXqZerrmXg1ZES8o4EvCA77Uet5CI1E9zs5z7noESWChjiJYBbpTCf4ETHCrOqrY9jv
Q4R/UyUxKKB1XPIY1AztQ2qei25XqK2WiFb8elJRTNEXwxXuuW4fhg4Dsab0iDyPjCeBgkVkE0tf
IooxsrN2EDYu9ZevGsES3k1uQZ0RCcoyMW/yEZ0ox7A0oBKsYz/ZI80FNTchslFQ4ww81HYmpmhj
lOd3Pvs8WDIIS+8ti3WDJh/loNgEATXEShe2WCgr5LmhEACW6jmF0IrxzGGNI/Od7PU0ixJ8+sFD
Q29g4cxTj5pYchW1fLvOgsbji75KXkvQj2rkd0Y+9MsqnvGvYotwPAkUzZ7z/XBxMkyvnpkgs9jA
f7m6Fe71UXOL0ybDb6RlfsnN1Ow4/ETEhK5nfZ+hOByWZluLgcTGkfEp+VT6nlcXdGTZxG/hSlgi
3zM13FV09dL3T4jEalQxUknuO5ZBzOOx6iYCidfG8iuzu4R97zbcAQe6/OBM6x/witkSRsAjaiii
6R/2MrWHnON3XmIehwhf/qFKcbTlP50CwuZlIl4LkNrc9CCe+YSOiyIlOmj1Vtie8XINQGBXm00U
0vxeCFPaRdA4vtC0lwFXpfmYc6s3MyDm3C3KkSzOWIHB2dfi5XOvi1JaXubefCQmUqeGSJUo/vkj
wPITGfOeWMVXXmy6aGfO2fedKvVZClEnpQ07D18W7x29CmMDbK4mtnY3mOJMSQMdsS+NnTojFUWL
979+4EMiWF90AVKuoV/bzmcZlXCtEiU8CIqbyKp9AsrGe0R850zsZBa35O/ZLo6hFvtRm0NrLj41
U9aRfjM/sVICQhF5Zps80OoJs0jqITM1775paY0ofh05mAIIGbaHd0F/ZZG2/Rh/uNGT1/KoPPS1
sKKdtMZGG1dR9wRsE4TnjOJnWUNEdkpJ1YmPlUBdru02IrrLAb1M9p/AySzvkn83B7dkZMfIj7aS
UNAwUl/k/YUbG2GymvApU+Pb8oL726uEUcoA9fIs/vLCYcui8a/9ewlgV+/DEYwMXoRkmhyjj7JV
Q0/Xv9U8TpgBLAlA6N1MGY3o4GT1h0gPO/N2dseTSx5hOQUyQVVoUejP1wCsjWKRK+VKS/fbaPuG
ItSu+VS/m69njPPP4/gEzgXeoF1S/183HnyX5Xzu5s7TN/9g3nxrpH48uOjaUejQ5XyLH72yEt5x
J1fbwjme8Jyvb5LB4XRSYsPsV/qNAbPl40uI+chK3/A3KvbxTnsTtKH1PWoU7KjGDkcmVZ9XQS1x
tX75GUxMQOMK54uuEWG2Fc3THyQ1SkQDvMqL2dxYgAc/e1DyKQ0271kaqGlWrgP56bBe4hLE58VK
JiWvfncoyn37j5PAK9IlaeRn9ISc2qGXNPQ66+Bqa4d1JH+rONW5Qkf9Gw46o81MeO9T6CTPVqMD
BrgA5vhbqQZcI1XNpwDCPcHDN+eCiCImTgnTkYSbTowjAZGTHDvBmYT7D5UiF4RPGc/7ovE5Htm7
dYOwEFwh6GtVXwlFH8S3n5WhjX43Rs6UX65k9H/wbNbivLOqlduWc33Og7LWLTCNGQIDu7k1hQgd
Z7ThlPYVBSr/aaUl37N0vZJk4ZnMAVF7idhbFaZnKNFuPjErCxpRMb9/p2Nzf/7i+5AceBHl1qLH
J5EqmsleNUwXaLQsayjkMhXiBgX6u/BV0Jkdh1c3JvniQAdjfJ65Il+1Raiqf/8hwtyPRH+Pei1i
YhhPABGMiqxcicD/nHZs7zZS7ILd/XUWCcT077APdai5Tq8kPpwm9/Va+OTuA6lRthQ/ccBzxwE3
hzPmtuXLuPiBi2IiPW+WIDgXUgVIbEqUlwPcluIF4+5mjIxPkCCLq5igJPR0LZendNmq2BXEJZCM
+8Pl485Hy0RjgIiWfo689KC6fkQG3yjm2aQmBSx0IiO8otsjCkgV2X5ywyeHsUAO0kqQa91A3ovA
UL5WgvF48HDlqkvJtKheNREi9ZxpGGnak7lFjhO6ecqSFpuZf/xEqpeojlrKabV8+TCjU3bBeLdf
HnS9q8alYwBfUosHDlGvhjIHLXUYh7W49fVivNGb4rGoVLA71Ts5loZ4MgxiXEz3vNsuQNMcVS14
2ffxiGPfsYNVRjJvYlxhjhWrI+IFLlVRxJ8royc/bIBdxz6kZCZ1fQf4dT+XdJ39cyvj4Bp0jduH
t1W6/wKjFxxBbhqGdoUk5fvwBYykCBJJG3bnuTR/k/jMnxkVLCG6kVtj7BQZIk7OLDUOY7mJe07C
EzugsyZCmu9y4tjCPw2oNMmCBRol2rzTJ72doAsNzzUG2TaUM4B8h+X8+QKn9MIugmKwyw4Qu0o4
IFtAJfxsx7GPWzmdXws8MhWAy5ZGzrLsh0zbYDgeI8JHY4l2iVutF6AqLNfpuS05L4eF3uq9uEK4
6wOTHIZoSMElYnmFpB5aL6kEHT8WQ7Duk7AdekJTO4EYzbTh2c8zF1POS7j57qoKpVJ1+YNptbpY
vj5stxs8AujSdgXHf3u/ZMXYr6L2CqMXyYY2NupWAb2lR4ndjZBTX6hZWPGVx9CgtoAyJxWO/V9L
3LyUiUJbMhUXlBCXiaRJsoOKcEJJ6JQWB8x/H9/GlG3nUw8A15YxjoM9wdjogQzt3r4W6vSMUSTZ
vLckHNnxsfbWRtumTY87vtfbASTgFjwkAPOKZ0jOTKrue47b9keRmyc4Tivs98wEyuzD3OTXLcST
IrkadsYwC1Bwix7J/241381Znz4nTibtVTNuVnadf3DsUk5t0xou2Shpbba6izPcR8ss6r1QHtSj
T10EzyO+33NA2qNg1Jd1ZD3vltITgiiSeMkeis+6XFFaCqUJM8g2JGAwU1p1dLNfM1fXZtcNbfnx
UYg+dBoahGRCgV/8Hm9+cbCfbS5oAj2C7YrF4nY92OzCtEDhPkHXTPhkAQeEVSEaIYCgwLxKbZpL
e5e57BX55ftXSOd0h3FQe1U/ieevSokPeXltVurdQsX9lk5NptQEl8GhvQRxin2rzg7fgGm1XD9M
XfJZ47sP2WZR0ffQvWcHJQORW8oCZWFUWa07BFtiZ8cNGdtMMe9Iz1TsFcE+woDslkwDbA7wRY9J
yk0yuK+h3mEThaxxllmuLn+C3o/4hvtWCZ9dIv38WS83emlFGzRMHOpOHm30RQmWR0Er9S0pwpOr
YAiwI7hp7obVB4RFc5eP2ol9YkQ5FJVBtshq7OLus03BJ7U5+wDfDsLx9Yrb74fZBUq8ZIzEH0CI
45uOuXQKVPT8EiV/oVDOp2i8BHwS3JO+0VC9GOD0pzfT1G9wnsbxNiH6bRodmaYM8KyXlm1Fzalp
Qs0mYTscGKoh9XOL7L2RFLO0enH2KdtG/NvkjpmzLY9ua6O7KuMV6szpGU9MwiTojXVlpQ38xB8U
ZZQdoFPB9RkXWOWh+SuyBxvMfeT1bM2EhOsXXTjzfg5zEJ7IGH8lH1t+XYOpYJeAowoqUcFK6T3D
YlGE6LI1Km1yHvNHirBZuqtp3HhfyibmJIZwq6V5LaeXLXJNReF8D4I54rvXXwFME0/Y9zhYO2IV
f2bQwd9o/Dt5m2ZE7/au9qqVeks9S8KeCUwEXAoDPKDk5wXvSN0ilhPuAUEzIAJW0ku9LHTCUvsy
/XyEfw8QAFcw/9l3KHZLacVgDCF97EhHeP/yZs+GwAeSrz8KuphsRNBXIN9BttreTE88qE0lTg11
32cfsfXxoEun6lgWSUBwRkgaW9wzop8EdJI2Yw8OQWqO/7PztQEGgOcLtUMDOJ1a63EZqRmtCalG
1Yej0Fri1jz9XL2LZ3NoXksLJrtTrrLD1O8uFSO5iXKlXM6lJv9OO2Aavi2LA8kTWZKSb1r/lC12
J0yH0Jw/BC1BTXMYrP6YmIjpznHK2tVq8FPTFe3ylMs70+umqms6cCsPDT62bws2RJhwxIaRhKGq
5BnG9YXRnveujLWCBdIpb2LaXt0Bvj2zNiYqmMmvrKJnsuNNUeyd/uZnEBNbmWfozI1WDTWYDPcf
37h5lUu3vAHY6sJs4ao92uL1rCtcD8sK1wn7johwzovCJQHaPKAjJWpxaVthARrVBlBO/YPBSfzy
GNdWghNzd8RGXCPouWLdUhUpoKxxqRuM+BDsmBfAAS9s1rfMhgHdH9DL8eF35Nq2skzAZTtXcCFC
qKfMXnpamBCt5DO08lvQ2RgeBh9KBOklE7ThjQmHE623B0THov24diq9M/j9zx0mSEMqhXCXkSEa
qO1z2iII0H2l7n1y0bJcWW+KZTHBhGSNZ1NfVZUs/rSi10zzpUhWOQOvVfktPHI3yvS7X5GYDTJD
2MN5RPeQkfstRPmzJtepsETB5Y7V7JeisFN8u6KuXKweodDPujdKr0TS3TVdW1hege2FOm7XnTaS
3RI+L70/GMFg7y3Z4aW0MGMY2/3jWprpbB6vu1w1NguOFEy8gxsOvxLqP8wUA8UfXul/TyQuJyYJ
WiYomup2lkVFteZnwKpL3ZnzePeH5F9crk4/D9lUMnOMlEkt3sFyqvzs5LZ6Q5h5Rv60mH9RF2Ke
n0VZ10B8CPEKtcdR2SPS7ydzK0yfpq85W8BGNp02T9bX749U8GAfqmn74+/bw4BeG3JwgfnBsI3u
2keQCE5MxzYFeA8lFunfYq0BA0YiTol34SVaCtkenouBbULrZXMvhicm06aLcP1oeWxo45BHmuzb
5A0juL2Ctfml6ERsPKbr6gFhaoVQ3lLrbjq8tkFnTviToZQ+Cv30Osuy2VnzEyEyrz5co/hK0Ivh
UAL+d8YzxaXzwUYm5vAUK88Zo7i49neeP5ML8ihNCWVtoF5MCkL3CpJILJDKUstUcqV7T1+Fuxvi
dErUUEPT/XRcg7CocqEsjNdG73pkfmFwmLKMHK3yMSsiHUgaLEfAnE7RfK8fSVd+nPkBpx39xisi
793mnIbkKZUfGDaMbaPhhWDmDvohoCd14FgYINoQOmBdr81ogEjV5zq0oX5o0pRkTNixCwZ9pD4r
zFDf0/0wSFyeexqvN5wu5NmHgVHcgs9e5a60m0NZrDYBKhGXWwm+24Jm/z5GPU9jKcJeU8YTWsvK
QRJNy75ZdYEAO0c9IeRa023WRMRdGUdpGZGQTT0/yLq1/Ekfrx4RSxBtrirZcJIz0MvHMLeK/tjK
JN4gzDckJ+Sg4eQwQygG9W75EI/yXU8l7aivb8K0K80ideYalJxhc+hRLMyJ8H7XUnUjLOX34j9C
yLdAUM/7J99KGwU3fGPX8x05oLcsMKYJ4XXUyVzP5VjscBWIW/dSK1GPRDwhsU4bOmiMbEfxrKIg
aE2h5WTrbP6/AKHZPb24pn1w7+hAgF/kKOi7FLwXquUMA3kSwhuTj3ftq0UX1w0KE8+hd2jJoDTR
aa/fJKhXhDI5ZUYSIX0JxQNyI279ukJFxBTAbZgLD50kavPaDimSb/0qQbwVFt4IxNjPVfDISUP+
S4EC3yBzNCzyDV6SMkcMuRO2gVijMgvVWTvSuEU3+YjYZF53tCki7TO4caIMO7eD+dVCuaulPXvC
SeE9f3cw3nzRZ5sbBBZ6+aSYDlf+E3WFVZDKw4hygUm/f5xDelMGy7u++JkEyTvuiC5Uun5lnHU3
g624XdQL0RYx6ZX+QlNMO2+A12XEri+shUlml7NPmd3FXQwWc/d5GaOWwz8ecyjqPlHL7Ie7zoOA
T+KgEB1CG2BuxHvewsSXtspY/fk5y9LRLOz0e9nBZEnN0Dg+hC5hXt6SEEDZG0JqCwacGPJUg64u
fVSaPEFxCuTsQtem09oBBLEnZ5/p2XKFrkEiexM8i5jKG+1IGk2dnKss4ftcTuv1wbtV2kdNSiEc
QUI+KBG9qJVGUtsuQ0LhdzXP/+5gFFEvuLudNa0QnpMEXZOh8SnR7ijTHIVyLAv4/Jvq52o7xqtD
kWn5nm8rSN3SnZL4n42ZPgKSpNDUyu240FbYjC+yPNhAU5kSy55al4FpeKN7BBcEjo9FhP8f64n2
1FW0mtGmgyP26adczaIslTJmqGNoX0eypI3DeZdviFEfkGHVnc90M+S9pzCqAlnqIWIdR9mt/iFh
olkqCLFanC6yHGM/04j9mQhwhPZZXoKtavl+IKqRgxtBt0xCzHwmZLnTsQue9JC5pTtP5a5Sltxy
t2ALlzjHpjoX6GR6MyOzlzwYm/iRUpZVCCwB47mRxlCjDl4hE2oEQi1wBqeUquuOKVQK1YUWH+uc
13lQiVd6eeSZ+Ai7f+pLHgBMmS2EZNrqTS5W6F0O9x7SX7qQLsodGN7MahRTMxxjHZTAFNK2DyzN
eiVG7VqAbdtGMz5Kuic84g1hVS0416a/RjeqPDCmzHAbY0t3yf2h+zq3mG4VjIjJZmBrURL2Hlm5
tUn2D4B7ETTdrcyAhz07G8WdvtQ84QrnzF5Zchk0Z8h37hqMETf5jTshnGBAg7Pv1lGnOj9PLq9E
aTySCFfla8c6v/nXZ8yD6+F1er8DthsyDKFdv6EEDCQPzm8K/GM7KnHGZ9RS4J+opBLpcus6BfyP
FSmdqWH6rgq3/y3BfNLzpDiec3h331qT6ZvQ/GeXe63XcrnEDqBCp4sl29D9h9k79r7mhPcyLPmO
7XSMfZCnVEihiiohO3N8iGUF28r5ZkVWx87RRVVYLo3gMNDQkl1wApvEsveG+gNA8qesDAk+02I3
M2lExRRl1wCLkarwD2csQQeksvwJM9XrWBG3zNo3cFC/K9QIi0lRJ15y8EDzkHA8DiclECt4Dj5r
SDonPLCcWWI3EcbAXlLE4ltE1+fnDf/X8k2wffzn1jo+5NTZSAWarEVG2h2pm1p1OagW+1JgXXJf
O7IO1WBXj8M5QlKX5Pg5USNsRPWTdGCcfhgl/q17QCs5MZhNES3d0COC8Hm1pftZmQQrbmtQ+CS7
wdZ4yo1ca/IT8PkBqTZjHYHPASPiH5xE4Y5s1wZA2F/y7LC0Ybwv5Dv7lvwrPa5RyipARcRIRWHI
tOdIGTmYC5/v7iipVBexkVQXtWSmGLFQq0fcMlL+Wv721Ocz8b8Ip3JCD5sqdFOBIn8peMY/+ro4
cJbGHilFt6/6i4p2KcWB59tfTjEOBUnkyqs212OBoR3OnVySTV1ih20/p4B5giJlzUgRlBBrlIpA
1vN+CTsWC/WWvc5kpZDk8yK1aSCnJkP+AWMkwUbd1bhtE3ci9pfX3chuX+J8FELGpZKLJZQWjP11
mFCWcnM4WRUun50iUUNICaUYP6WKk2xWj8jxubUWYPnYyvFSWV3Eg4ds3QbKtNfbYiUGFH792djH
saAKKI1Yln5w30hFs2JWTRixGuklYgQTVPUIOcoINFEWFRTqZhDBbbMYc+rpaiFYbWxC/0zYbCyd
ydbwkNeLpkkMKnZnfQa2HghqpDGTJyNHsh+Rrb1GzSQ831ip8QZy0ko+m8jsnllnrDkP2lJX8Ifk
4U4BSuYZI6PQkYhvGfbqfiABnXBqANuSqbTd4h2zRnMauZ4c9nZXjCYbSUy0Emc6cPbNnz4fee7h
AyKFVzlsZ0RyLYqYbcw9WnSCHgkMwMV0Ti9eaoYLwOrCq7pUwQEUtEbMAhGhrWIh5s8X07juS4wJ
Apa400EBURY5Yb8pbN2ViyDxJ82LABZlkWy4BmihvYmwCAOxRX5YBWoEBP0HWeY6b5nUnVFPglaE
QXXBgn9CnSoWC46Kvj/+5bpJ94AbbWN4ODs71LM7pCjnB2Sca3lw1SE2+piw6pRSUmtBoUQxd/By
2Ffz6V9WP+FlW4XMG59WuJCUVp1CetOSITW1eshsN5sBJy+1Az5OJcvpvJHB2SqQe3uHa0I+xMPk
+Q5FrPdcY6+RXkvPTEltuYo3mbNfbDhlw37wVqAfJf7zTcx2fxzqC3jrrAA30u5fEvblPPKTQ9qV
ap+feBaCp9a94i+Sm1cLS9nLlkP0Gh8GrTTpC6IxyKxuye0zO9rlUACOU4DccKXLA7f4cmIFOC6x
AOAb5Bu+tQ1uSzeQBuRYeJ+D31m1XhBfrsPPJd+c+DfRbNYwI7hr27QL3zXWWpb/ZVhDgybLxSPF
bsWOHwhgozM+o8Ql5c5LZ7lLo8NvpZqh0/HkL9o8Fa+S0DUJPrBME28qKxgoT4NKN//ncGoosbqf
+SLq4Oxkv9O1zTPKeagVE8K9jJHNG79/+Fwh5NfohJvtagMFUGwdIFQTE/rtW+GUEy+9Hc7R/aar
Pl2oOfx5pH17u77OhU+BGbVgPP8lSmjI9Z0GNgWiAag0uWLdJYRDNcmLt97PbLnJ8OaQUxA7YMcR
MHo2iGyaEO/FYHIH73BkLWf/UjUHqjVrEItgpC/EmDQu/eLX7CckXl8SMDhsan4KfAfw2BBC133/
YhkV2EUxwEl0VxPv8eDMz5xMH2sZfUoBchqk6AIzsy6S75YmGKa4GJPHzxr9Dz0JspQor5onQHTJ
nThcqjh8N5RF7RjYHoMC245Ug0/Q+z2H+SUgCR91BnGoenRo6sRkbrTyiOC2dbJzcDv2Zf5iFszy
3wzuQ9YSDpy5cEyYCV5hmEbWXc1QiM0zSgMm5P+nrPrLuoFEJY4wbYmHuvlioOg/mQQ9A7PYgao0
KGXRFCcMAN0V8a2f7zdjB/SAe/SKtggvdbzM852VhMAAL48Ky0PHRW8T8yUylmO+feH1pL1r4vIB
smra751ClX0rHbaermdvAbo67o59Q88RfTWRZkIvFYMTD5vfCdR2PbWhjpz1Jv20zBdu7uDjFidj
f9trC0j8w9c2dYlIL/B2oEXUeRXl7R8+NGjTQl/EoKmSO77TCgD+sq6/qveCvNgakxaZTV9SqBZ8
1OCe6MAY1J2qbg3Fuve9KUmo0WVlUgePevOaJc99cfscG8GX1ZH726b3IFXTYwAzh9HG1JcE39Yr
GEPgMnrTA03Pg+2ko/Cs743MFUdEYeiSRDBDojALfNv2DFl6yIiZfITio98aYIvd91XJwhp8feRS
jZEiFiU3KvOBfNXN35ubnItx1FHdRpzc03rBREeu4RgU42PSWsm4D+EcQ6o/PEp0slMJpuVQ0f+w
F4ezNqGghq5FtFy2bV+e5RB4OBAzsPTH4Jq+65gTwHlT3TuiDeIQdGykMO2TV/Lc6pCkntIEEUvw
M9Jt8C3oJpCqh8sjyx9zfOk40UBX4M19ILE8RD9P/GEr2zovkVA41NEMTdYibS/1J0nrdNx5kd/A
+N4EimCOWzfMghUAMcArGXyjCMM6+NsM5jDEZVyxED2xgfyRo+qdaNZaXj2eb/7DWixDG5hIdmV1
+FKLbdDqPAJEau6Nbl/iwXOTu9BSbEwJ37AvNPYxx25d28L5e5/Ff6al+0V7RhThKWsYjQOil1PN
owovVo8lyhKjTnMB4TfrJJEkpv2L2KObH7Go0dkMEguOMT566Y3p5CBSGlJdydD11yHfT2TEbGaU
b6gvy4RS5jJnKEwIQD5leDriidS90JbI8qraeRAU/le66f8Uw8x3oUr2Sza//nFCTSVoUs5/jD2a
fhfADQzxb9UUfu5mqH8Mx7xvnu/l5368Dm419xaJj8rrpbdDR5zRGlwcR2mRE85NJZrQAGA0XfJO
d1paA+DjMfID+sbi5OHTzRrFNuPWOGu3QXhwKr5ph4S/rNdFDrzxDVBYy+OcTpHzmm9WkEbHPwJK
NGUy4ChnwecNEbD2WH3ZPK6vRAum7Ni+2/yReZqk7yC2Iwdbgc3z5/2aIKbguazhN2LbCsk871SS
ibmrb5dSKq1FRhA4t+ABhm/NfG1SYinaH1Qdh9PA7WjxNbgx4T31d9XnxQ08DlkIGzaGsIRtzWKT
AB0dZCh2yH2CjORAKtBxiUrCnh20pgqvNK67ttfygNMEN2vsKyAvp6pAtI+EhDyf0UYt69uC9Mv5
iJULAp0aOjtAiZ8aqJTRRuRNY+GLm4pps1g+c5ffNtpCAdhG9rHQAob7nB/NzN3/+zPhuf0S8KrF
GGSe0WQ0pIVNWYDrU6mbh5RlHnYbAlRCyZhp0tPYeMMxCM1mRfANwr1rytbwpZXGWlhKkWZ6gd0T
0PEqILZAFbRDtJkmyW3I8e0BdE/4Sn+y6ULWVil7is7fXGe2vKBitfiVq9xhjqt4GRlZ+I2IfVH2
/lJXgCNJHxgtShX/JAmXaxmOs4Nnz3P/oZ9K8Piez7tRkHkbjIR8/VAksiF4q4amSfqp6XU13ZlW
AnRZv+nR4oHcIrjlq6x4i6bJU6VrRqw1DwVrNK6sho7QAbb0FIvhdWAH9M3tDuHt+83NvpRGoyAi
sKE4uWpXmDjcTWoqK0mFHoIrOOjSueOUPy9bOm9aUSP4pxebtWslX1Gyw7OXPG2DDaS8u2BrZtCY
OKscIvdpJ1t07SALWKYZ0rZwx+tPkn30Rd3KtudFYHiRYXMGV1QswvIqD21Yw4QxqEVCwwHKmcYp
qIa+c0JBmZ+xBS6Qw0de1vfkPUcGZ7cqFi5TzgWAhqEUrWtKdjoFVConBBZlg1k6/7CViNys9/uQ
1A7zMu3ckHxItQ697jy1YKtcIu2j5vd9gsPa9yOCTH5SufWucDFoK7uTGZwRm4w9T+NDwwEHpxMA
0emlIQQPyGIaSUx8/8hyLnMQ1flkIr4vHXt1jymlzZ+uRBke7OiY0IUS38jVSkNUmY526I2VprOK
ILLxsVJfRiO1hz49Eg0i1xtQBN3AJTOJL6haRtMMRsmtPeyWDod8ewOGV5zoCW/Si+j1bgadjItv
E7zZVYjIr+U9Hoa4o5NMqLL408XPFgsnb6L0erm0aIzjNgB/mJExrMxaII/vAmJphY0LeSkNT44z
FBnEMJ2SdHeTtxsWgOzwz1+vNYFcK/u5rHnypgKUl3r+BATMgD8Vd4GDSj4/uzvpFBvTR4/E8Jiw
ieqdowFI2DbNhO8ZJaoOPWVO4cFhjisZmRz669ok2ak1hH2bakTwAuoIj7cxcyzxkmEhaBC22qRs
86s4eVpei51LkL+gfpN5TJ+bSKeTFFWC6Bpr/ywDy/dn7F5tyMP0VDzQaFusW6OUT6LHi64w7c1A
7efBZCZt2y224+mxYTLlP+27Msi8jH+Jkzm38SVWAjsjQqTLfqJ9pIN3TMjenEwRdpI04Pdh24RX
42cuoEvjX1SCOMgPt1o8gmAy9cvROO33gTV/8shmiMDHVOsDx1to76rLBA+K+zpPiWytsVJT49Ri
CH2EW7gyRuLoekefHvJY+2lEwhc2Ba/Wz1Mg1RxQvpE3p8bYW9MOTH2q1I44NOPFetBwI4JtaSTx
0BdHSK0EY8ODhO6QgXG2BHP0BvqzqUEycTg9dDWTayK4G+naxP/7M9vbcbEiSifmO6wLE7nGfZJr
5WF+DZyUcH+0t1ZkYHQUhgWKGd7Jo7MUE2ApyVZi0XDLQScugCxNH4MehsMf1P3v7dj9lncyyvD9
RAckid/0KXGYqVeBe1QsF3pEQ9IyKw3jXewfFGpd6HxAPs3DqPWGUUSM/528BfaoHsYrWSlozIW3
INtnFHGyg4emaZhF5zWQx+eWsx+4VavtZB/Pm1fl/aCA0QqmE48QXDkrJkLyTYvYPxUey3JhQbOc
kkupVt4uXrrnUteVRiWo+Mlk3AWU1jrsHkl2HiG2hS1RMKp78reNpbTspPp3OatYEtnCO5eC0M/U
kSPgPex9JQx5J9nzgWSlGleMkaeIr3x1ECA2NTp4pJwWR9q5gzM4exrJfNTCarGIwryoZr9RMD4U
EWyq+st3ouvccB4Vx3pwVffmXnHKTi9I5gLPoqXKppdD5MIgyfRrQtESVA436n4op/SWP1Z+8XUe
PfE9zcd23yKe8vZCE+GwhMOrk+ACcciUd96LYCHut+yJ6A3i0JDTbbnQycbYG5w9CmN1aC832v1b
Q7fXFyLfxg3B+Ibn3lHKts2JEc84jMV3AKhSWoGoXUsPn4wjCsQojCqZ6mkblxOaF3idw/my6W7b
yKFZrXrKtZagdN+rirr1nXveaudkz9n35pSDJH0SOPNzuO0FPFol4VCrV36GjLbAF8VwvUslp1Px
4XmmyVOqUYjfAyRC4jk3QIn3WSxMXEgjQ+4EKh3GFappJb9I196T57gIGONRsbaYeOpL8V9ETWQ3
GTbwPlKIivNQeaQdi5iT60OlB26bpCB/JJYSgjCGlVNvbXMqdYMwQ6pPkqqAOTND3ZEJfnNSuKJQ
6VLXTphEtu8rbHnJRXpUyX+zzodPckQA/Rd2PpZwXt/CfNcQai46m/pMaEwaXLxu0dXbOIxJPMiw
UcFdAYV3cIQ0uidR0yBsg1ZPl/Ggs2IpYFjdUh7Q1nBgO7t0C/70DcWp2nUNcBLc37AUf2VpI+0E
HWNEnYgS3vQZFfYjoSenwamKt17nURUZQ7g90XdT3Ix/EtDfhQ+gp9ymGU6zO+Qmj9jb2qmXeHvT
4Na47B8wW+gmz68Zs3sO9w018pQiBX3yAh2/SGXQ5KZ7JOvvhfJKGp5om6Oa4ehoPv+4Tu2UDX48
MovrhaSct0rwws5GMiWgt9u7Wh91P+hijSyj6+PFa8+TFvn4u89eFQiuaHPEi0eiRSb2cJmrOh6L
6Ehctfe5WOZjTV9GKIuKonp/HSfMepsqa4qyzwoRoKiGaf360KqXlnEsk0LUZ2XSD21INL3560VC
fVemJZv+mBxSWNpy2uI28uzrO1JF4fBzoF6IC2R4QP8iLcYaIbp/WaKBL8/cd/Xg4StvXIhapgDa
u20SO1GSrdroOaR4dIzlVoapQw0Xn9L3sXqJUXjo3yrH9hAGYODYprQST5Tz/PDmdwmD6fX2yowP
+SAqAUwR9Y9NZqLUqYmwvNOaRzOGa+7092KMQ3iJ1cW4K7rRDyECBvMuYqvpNyldjO92BeKbzy4c
DOIiF9yq7qWm7kr4Ggef6/5watqxB3lvS1qLoGx8SaAjJXuUV81K/+GZg06D/EZbwfPWIWTlTE6s
GJvbUWs7bMacNgKqJakFQy2DEHVqLViOCRF9qFsZHik7veCgT/ncKPRujGnZBHdZ/KtdGWj5EM1A
8ujr6guwoL2nqSEVinGSYjhnXazZIzX+mwPjEkpWIuUbHpn/b1EnsBgSowzTzO5YElyU8K3++8fe
G//M6C6XUQUAYX8fg66mvx1Q12PntDNfX3dpILMeY5KuTWV0UrWYRXEGilat5aEB2H6PhyeUobK5
E6xSvI0QN1DpRRzPzntR4ft7fot9ZIqu0aQNfSjY83Jv5EU2Zqzz4sMBPSXyyjtZkr0dU40nqVgP
vbQ+2g+RlmqjYhc6aoTyAs2VzgBy1pCnfAWClDR2KVVHG9qPg81nocl9xHxYIYxcnS9UEy7fokWp
eoWQSbSa9fAB2gtGBzrY0HXwDBHTOmznCXXSw9iff6gpRgNOSY6rXype+oQ1Tk3yWigNy5Ity0ZL
M46wEKZLFCdvFbtGtB3jBqnQdO39AKOFFho40xVSmASGPS9mf24F6LI/gslso7kO05ZbokJOFAKu
4e0Y1G7YDupelNutVCj1UYHWA+YuerwutE4SPI2BvRHFCbkiQ1AAvL2RhNTgG3oVbWzv/6fbAiaZ
6ArVF3YA00dMFbq2ioBOCPwugvtmUyk3Q0l5ItlitOvNlvSq/rdpDf686Us3FhpsCS7t+yqENcKS
+bMYGU/9oEYvPMJQif/QVgGqDS5efrjWICyT8yGa3Lg4TMcWZ9OEVDgJcO7i8XdMbCCY66AzggL6
nAeu3/dUlJPeF50/ORU9j464LFf51qrcYIYyBrCchcZAB15+itUKvrsTd61ihDLthVAfrjOX6gUF
6ST8MX1Lda0k6uVynyrq8qDXrxhDIxnFXJwq1WDWColtf/4GtAFvwlnCWKDmw8rGUgQG0YZWQUDb
shY0GWNGcBl0w+g6XHNXFtDKKSXfbEfPVLPRELtLRVwSTZJ69kxIJW18uksh0x2M7qSupU1paHwT
cVorB1GDHqJuwaYpcCbBMVy6wp8XdpWWb8PCVh7FEw+2dbiAFswAQBYn9nAbezUAORYyZuMlWd+g
OMZrgz+8iU3GRcXMJnFMpFRsUbV7FrCrXQ+axoT7MQY081bvYmjmlG7I0odMAzRyVe+8g+MuHGPU
NwuoWv5ggperR6qa+OOiJYXoVYBuPq1UHCQcOXMIYJCimZCDQocT0td7S4c6YvlKVEcJfbz8PXPP
tHROiu2lTJvkbHptcObO1B95Q9I2kr2IrykNJUuk+4Om4zJSMuAlovPrF3Dj4cuqEIJwrRhGHDBx
vsYrdP8dzgOUfvprJoqomi+r/vSVuTMBkLaGxdyXZIgPK5WQL9u06cTRcvomLL0U7O6wL61XYc+0
ARc+rd+37AS684/jrEQetrMMUgjx+THM5Ti0uX/EiEw5nM4sR644eidowuiJedGEhXJJVbT4U3C5
8VtiVe0f6oKpbK8s5k+KpHRS81GAER9bK8CLGWoS4zNeDiYte2NKtG4tmmgXPrMgis6J6EYvunsp
7XFEHeXPhmjfsUcThm9AwLrm7VK8jFNfOFakizBvkZho0N2dAaj+AAU6lpMt6N1DnOAfSaxw2lly
q8L49papUcnb3HJ2fNBjIIZKqsLTBGjIAfsor2u/n+WuB8crL3ontwV59oAZlc2j2PeIxDhTc031
z8sbHDBPm1WsCIFF/3l0QvlvboGl0spoIYH3MeleORblF4719QNgAG+fUB+5MUuZwoZOjbnh0M6Q
YsU120+5SJfj3bMylFbmDRuHxBEfmz5iGCKIPOlTEdu1bCeVo8Sl7471LJeju4OCIwhOHPfM6i3E
LKEdW+el+glwQAVgQOcVblyqXu+/0V4vK17LjsW91nNumROJg6t8szYDcXhgei+kD5dyKZY/GDtp
YYA8vVo69nrzuWLSOQOVmGUSKQxAh4wuJDw673FuwLk1ZOJw8xdvc6BF5w0o5HNGzMFjoPluKC4g
xv2iBRhpD4HWAIHO16TOqhGnG21f/KusMgPDnotM9iVbmZt4NcTqRSx2BxMIawO7gvXUBfzrUcWf
OwcyhYxA5OnvfcGTD8AX3fcAG2IJledyBvzMYQtsPpqoR4E7yV0LPjoEQnjFETwsaNcape+Ux1au
OhVS93Jz8u6vpHbPYn5Tpz+XS6fx0VgSpcbMoBdoMIgwbQWekNp9PxO0iCXI9IDOzy96BPa0GhQ2
7RaELVpIxOZ4/bYUnDuWgksv7SsWBb0z+gkhWXsUb+b2nFVCEH3QHD1WRgQA/Z7WxJsOPYawt4cG
230kaVBGf618WYF5RoX3Ls1Q0VfW4i9lUUqSq8eR+wPCwQXp0lYV1yJdKG87HVrmfX5H89LcBDyX
y8fdJ1IJ0vH20Af9EWNFZEI4jlyEpRB7WuMRD/4EPkYMli9zGHFzl0sfxbnabqLcC7nqdStMyE8q
ytlAqJ/YK3KiPXFLjIkq1AjAVVggBxo7GAAQAvs9RCiSlxahmfKhOZz9Z+IvpW3VauyD1wtPe/SO
rc0E1oyDytJkxgI2Sb/hGoaUMTFXmgfkCKEbhliRdlNTW8PPDKtqYFRFxC2YbQxoPm58oXVQPuK9
dgvJgdacble+UZWkGnHk7A/ZNUqM4H+Q0Bn9p6VwpfaRvesuq807uj8L7gw4lec/gjiJQ5/xqcmt
Fs9gHbDZpf4NNUzuf53DgVUBlqvLqMGxYZ8vYrpLnFE0dI1hu2xRQhjV8Tm6nASjhCpRaiJqBRPy
pob8cGLL/U37xYTOfdlyZ8SGixXKEYF3YWxZGwJA2KCot3F7bnpx3NU5meSsqiHgMWxayenYdVD8
M1UehUyxkXyqhjJEpdlwCIFLthOU3TtXRD1PesiE8LxwuATBzKcHkMXFsDBafn832JS9CalbxMgs
rtK1tdY271uP57U54aKruSZF7RXM/tW75xdetKOn/vLrOBtM56vwBAj3xfLEGWAa3d2O+zxdjbAA
SIl+Hp4G05KyLxLbtLw+AOp5C5woIVVJwaD3EpdqzfQQa8Qk36PK0l5y6uikox2xR4WJ2uNT8IL4
X0Fqkobf3MgPAqp3LOJPC44If8n+uHZhfJ3vJ2Rc4Cl52RUvwYf0cjJQQJ5aB4pGqyHquiPPYR+C
CBk+tKxuV4xnGZwfTV0vF1XIqsZAz5jJdodDESwZ+kymesv0vQS6xvjYzzV5L+0uHIlbJZrAWl9D
44chsxbYetnmQFIigeoP4TPlpIULQ8sh/JnbbULpGrBx/RDbzxequdyAPXWoXvb/Q1E29na+JKqR
4ZjX0MRBhBi8E/UHcapETUHuCylzYphyFvygU4yoLwqFp+XSIPv+OgAXLbFh1HgaFClrjbCmq6z1
ZEVZePpgitulUzjlzssbotRPdAAXVvPwY8NqvazcgDYWcu2pV3TqwYOHqdVEB0GRCr8emmU8Yf3b
YBukjs2mu59JkljdwcR6RuiuCFqbK577i9U8rq1Aq5AhKILUV/xJYtWEndojshxpGXfCCfLkoZ5p
LGP6BlzKzUTf/6gq6yvbaBeElky30Cx/+J0RbDXKRyeCOzSzOwTwRoMUHStcRO6PBnSlszMhLzPr
nCYqA4lO6zlzIsC//pa+CQi1RHS45I6X65M0u92HDKx8kdjsZws92NWPQ2kEbjzoH0JNRf+pi9D6
4q3jhGbXQU5a/NGhtVsXBCPDeJMdyEIuiPsjKO7Tr9MpvDpa+pT4BolMCYujrSlP7+Ia9ESSLY0d
7sda6WcaQaWKK5ktyefPm5zuF2a/xBH5sksU/Ufbq1Ztn7/0MfNE4Ptxr2O5mxcCZWN+OmbrbvqV
nwmFfb6ouNd+qxdKzO8+4/k+kPqgsLNPKGtY/UKWrGoVI1C/EjCN0Tdo8ldyK1EkZbg4ML7FV8sY
tskxu1ramvTWTaEBJFS++cLlmUcPMeUDYoqSmyU8WdZ+t/rJBE950xqMmX+oavQ8H+Eh/doA2i/z
nPCEM54i7mxzY+ZoPVo6qw1R5jmgaBs3LELyqcskYbGnv2CECQgg7C6dxeeF0J3SGbRSCoNZ4KUc
O2lPnFVBJuvZyoc22u+MUTw3EhsvVqL0VO8erYzTvpEUZFqoRpvS2xU7a4yENgdkU6mNu6M4VdLe
yEvGaMhG4TWNhrfEYivxPDfyygvsTlUn39U96ekYg0ekgJo/Nbh+HikY+Zm0xn7CRKzjxwXGcRmA
yX0XPreyXccHeyR6ZgpN9RnAkUZxV5AAfHglNUyXRxOa/+z+RZvDfDY011hmDHgM+a8B4CjIl4sv
c9tPSOLHLhhDuMVSxHfuKRtOBbdtocuWyrqp4u7rnqGiYqh+f7ItEEbuFm5C3W6e2EFWo+4SQhyZ
WKpsv9WBVTASTIqhyM9i1I58aAxlURzBBUzK+UmA9JrnLKoTv9DTPvVF0Q/ZklzYO1wieF6dNp5/
A7DYZ4hv9UudOIyK+2IU/MgDjrCk513GiEhwL64Fdeh+TwsmHsGJvGOsEnglhj19PYZNY9beD4fE
OA0xwNBF58ozNXDeufJP2sTQKgwyg3dPx0SDwr6Mfmi0Wuf4HVtgwHvKE4HqlURtiK3CSsjaZjHA
74ZjGNIM6fX/yGnRfp6OxbnuFxQk/cJSTy8kijd/XmQG7LOFUPWdnhoUySeQLpzOLz+kb7bXVCP7
bti74SGwqVuj0hFQYyxdZ85nrKXgAuuxqGe9OrzJW4t5XFFBsxDZhokkhwq6gxUJHa5MSGAs3vn5
beccUPo8UF/w9gkn0U2FUMgGFlq6p+fYTPvvmFygmb0R7O3jDpE6fIJBgG0Zfkox6rCF1pBJaC0w
TzD9yV8VqlgsNn2+f4EwiQSpoFvlkTTKII9oQtlvhyJufszVVFED/teCQI4dmk0z++7VEEqkFps0
Ri4uEc1/g6uHVY9n81+myZQli8GDCjn/Dd5dc3rZ/YB6C4PxAtAZ+Q2hHyXXoJxCvCoPTHcs9+vJ
dDJIw+xftfusbSrqVqmNRv0r2hkM30WnYxd1YDf0cm3FIdvUcq13SuRqAgKJDa/Z970k7r/w/B8y
Uo++bl8C5zJjsQurwlcYLhpKmw0QCDQot13qhvD4BZKWD0naCtJQyNQvjPcimftB3C8ycMNlnnpo
vbMAPDJ/77dWZHnxHItAJsACK5MWjjedSLNP2GJZtje8I7ZOl2ko3mu7KTX9TeetXnVF51RaVKTl
rrH76fUyuZ0RLyOcNPY5bkP3CfO5N3T8qkaWe8op/dfdVWF2yO4e2s+DhAz199tKxWPVaC2ap+6l
1PNxC+U8cB555qJGcwpkdEGGd7Dbm9wi4WjXdk6L+WjFJ3T0Fcv+2igpGsSCXwU2ab0Sd+J5FdiN
YWmFUALy12Q4x+ewzKQFDycdTkYyQiMaCMARuBRyzEdAmI0qS6HSGQ3IUp0uTmcG2k5NgqEsqHNs
R2L/tiId8ebYdz7M2+4Km/cGyX+v71jV+u4F5XkAfH70ctKU+PE9Z5eDuG0dEEDiIvC6iYqiCUIU
QN8V8xSx9MCQh/qYeM8Qg3UCHG5kBhUksCfAj1/4Dqfg++//be3DfcR5sgQdTeH9fBeUzNN3Jc2O
rDtznuLvZVc0N1KWVBS7CCRsjISF7ablWk0HP/Hd4UXBI2poHn8YYLJMa91AoGj95/2bZier03h1
vKUTg3Jy0roBvm+FHFdu8twghKJhBAwHg63rL/zq9FDKFghSHzVcAbpYXurEwuIa0U1d/NWZAqAk
K/C/VhHz0EK07bT9InyDoF9ZgZ6DuCfHfQM6tsXYU7TjiluWObPsFVTJyDSBWlA5rgyNUWhlGfjw
UoWMOcWuknND6OkwttoZBHJUC5Xxryks2oXBsY7Cbcf0D5lPmFpWOpkXsLmOyYbMMN8kE2GKcXR8
QF2u97hOhtn3wJNGykELNqmM/eKjhYuxp4U96pEB6OsHJeWVdS80jNxptBMzSVY97xKSbS6Nn5av
9c697iN21I+NY5MHNi4QX6v1lsH6OTwugxUJ7nNIsPKUYYI+1Lq8mhWaZjivjA9WqXXLSdQI4vHm
KxAZaBqjpexa4LH3aEcEYetAAfSztkUo5weVCDvITQ7lPScS6ophC5v9CMM2gynZ9TqUl92RBaaq
GSitbjSUc0n/qjm1OEt3FQo+8cnHT7arUKzJwTV41pohfA0ha8phKf5ztZNpnkvtSW0noWdT47Du
zasm/z/ZU9SVzafRhDVS/Ai/YC6D77X9/IBAxUd/hzi++EIuHRjlDbp9GL0v4zdYekp0BdVVpbr1
XuLZvbPBvBdS9LrX5cdvYKwPVla97noz3sAqkeVYfi4PasXvLbhwi9NXTJPwv7wgU0fzpbAkkWv7
uaiN2QMAqelouRvjNoc5Q2gDIqCKwEgOMIXOTF4nyEJD19voQ5ujaKkzDhRkK5fg01r1vz78ivMe
XD/fnASQqBA94XdANiwGEFAhxSQBsZcZAAb3QXr32FFn/IBzfNnG5W01PfpSrcmYdsqgo0KY3Bb8
vI5uatgzjHJcyLy7dXS7CpZ9U3B8oRz0IMzkwhBnpZhLPCJOvsO+MA49OZ+P+XvX5EhD5K4hxnGV
4JxduRWHPp2dh5KA8eo9jrWUUkEUaEANzod8R37uYXy/D2mkOIfCFgiCNlqW41ADeSQK3yQyGbVf
PhuzluLVK4alaMDfKuKq6TfvljEbYgOFetsiXy2v0t50JlFNBac4rLz1geRd1TKH2NcYRWDT6c9R
Z0sHQtYG+bOTVGQj/1wOtkU2REBkG1Pu8KWC8dyEjeHoDn8fmVzEsPNjAI8Hnp0Vp40l+p4oxZT7
BECs7CHykdnfKjcs0f0y8zxc9yHy2K88iWAe0nol7uSQDctUhlleQeXy+fwlBSu4mLQLxRwQzm70
/WsmWk0fWNnWNRTqiPBrpJmAmRQaCPnuntqFBy1SC4aD3DE+QjB2KwiNfB1IUTG8Gc/WMse0r9D1
N0Z4ComT9qWl7vPSTND+L6IufH1IeI/C+wifOZgj+6LbNr1oyk1R6sn4fVetMw/rovanLQbDFsre
YQAWcpT/G6UnzfVAhyypy4LXtiePSPZR/kchCO5UeVOmA0IO9i+4QlD5LAAqZM/d88i2d4lE5LdB
1irq6lJWfviM6pvWen4Mz6dSF7eZdof+7YD/OCs7MZ+mNtHvOGpxw6TDu1vEsNoeW9gMy9cFfgC2
3CeFubabsp+EcZPfiaiouctSZq6AqSXlauah2t2ytOYd5lwbeDLga6pMKtJhrjYwv3sbtUJDXZnd
UrEKzSAUiVzNaW63Mw3HXlwZqnNEi4+j3lpx2YTcXddcY69wLOWVZs88YfbCeIURObm9UQ+JV5eh
nUenG+mmbgpz+9tCyqYH5sfu4brN1jBNb3j2QkKEqlsAwIG86uF7rEinUCA/yIfbRv2yw+jpcLey
7P9smleCKqurG9L7JGxrRIiQqVltRHwOLfdQuJEpJeIxmDs/VwTXE8+lNxUduv61F5NtuEPoTc5t
bhF2okb1wg604LNtCdWla6+Nqik4ISAs1gEoxGxfNfpIvww/jHpL+xCsSKM9FaxomBmnrVxHCQwM
qJfwLTKk+DXMgdlE4hxdSknzvtmhzLj2tB7ccDYx4TTfc4LOGgGHd0/2avAI0T/nWtfQy8H5qJ0b
3TDIMK3EdODVOcdO66AjndeXxGoul11sTjzuGVL66YDPPeGXBQw1ohy8stVqj/U2f14fsMaB+GCx
AWZ36rvHnkVhWOd5TPuZOJP0XsxroGRl33N1A6nDkRVYshSI5XjfHlixhs0zCm7feChpcnh8RnS6
bYl7ZHlxliz2zTW1bawsdPFcN72wV/1G8r/IVYqlDD9+Pr2uu+NEaAGWeKMgYob/Cjcg2cQTGtOC
NQpLYTXk68VOOrwnpHFQ9fqq6flBeg8q326K2XQNTFDoCRPpGau7/5UI08vgf9Uba5Pwouwjy5Ou
FrNPvTlnh5xU4+e9C2dldMk5PJ62+niv95JrUMrXdSs1u35T2zQbbSYJHHMQLQlu10o25Oi+3ZPB
1ksp0N9NLB4q7G4JEJNXdyjH9M+ovbemC5Y/hpif072h9pit6CvYUQEhGZZ1Gd6YGXOCnHFrNuxU
KStA+8NY6C4FbmA6dbtuyyJjwv3dP1qycZ8LnW4WNbpptHX/qcgIFhK/pl+lvo24GZJMRbWte6EC
Yanx84zz0y2tU0/jA3eMK7HsFBsRg/G1tkcH34yeB5OU/rZVq3JMjaZZNGPJVVW8IR+3OOOcE9XH
ZjOur0mS/67KP6HzQ93JnzWPVl0lputVHV3ap/RR43a0OVXo8/FRsxkNETbDpOB+FPEEGOiuAPMQ
IK3q7hhPk3LLarM4R3k8Kgr2Laqs6qCmsflcLhlOzcZ32LYhhspiHwOGM96kpcw0mS6f4Clja6JC
D4nvpJjcp7ZbYjqKxsEIZvctHg5uhflgET0PwLSoSkwaGRezSMt+OVMzxSDnxLlUJFX++OMp3Spn
jdcDHmDuK29QymBSafXlEeE/BrheM5ewTyhDpJHlmX48Xt6/hMFSsm/BkOcHrkoN5XZu4CJ37ACX
nV4gJNcp97kxFG6Q18XTJoh8KKq5SR2cZy1ghZhQ3HPsRYEP/I/DlrrbHzsaf6ARDkbTb23w8bUT
gTP7jPzOM3JiAcM2BgNr3lBCClMAtcMtBDQUYVxTuW2XHiRkiTYXko2eliM4lOM2zoB1coX2jUxI
V/K7bQoy28p9VKvMhPZd3enwQV27muRD12wP8NLIr3M5OCrZbOxGHVRly4mJAZOw08fSc//zJSxE
UKsAz40rgNXRLHD93zLb5Nbmtn0wwB6UZ8WPNVcxoQ9JxMRBbRuLelZahzK36tpv/OtaIHzN+5t2
OF0UtK8wHvGA/xyMwKOx5jubah5dThhjPRZesF8hSgisPxu2gjHeNxuuQ48tVi7iUp15BA3voWek
kvN2BMaUjVTeLjg6NZL/dL1mKgkBj9qtAamppJv3bLdPLUrlgRJfc4hJN3NQwbJiLhSVetYYLNWI
lV0ELdwYRvsSlBf4QxsLMJ/Iy/3uJoLRq7AU6t41fefaojEMm8D2tgydGezIUD+PPVFZiZT/9pvi
d3yh5U+9GHgj7kxoTpUVGS0ZT0I/RFvI/mMCBj8ATO5NMp9RThrKLKAxzs7+vek0vKHdNgJFdZLh
Drpx/xRY5K1Ffvmj9Kbv2Yetm6X5gkISOwFqzTaXcwBsCUzXcuT+S0dajsGmX+zBHXaR02ijRpEE
gT9nzgbPPRCR3by0F5hnngapzNmxpjW0GeBBMI8m9H7ro+p8o1zeYHd/p/f0LR/Muk7K1HiJYbnH
J3p4Jq4RaWCNm0OJcFAtO6A4/jTzUyCPpV1Bb9jgwzpF9T14dPf/8jEkqeRxByfRkQOkQ8FnplN/
YusmFEJx/fWueN/fSFX/jpYDKn5m/gL0e5nZ3IoviXuZwW4MKSy+7beDMMb77o0lPvTT3TqcLUPB
uNzvb4ID+cEgSICp+hFKZWQGKR/19FEf51lyW0NcdpO6canH67jDzLqLwbYrpyKlM7T9jMYrHF71
Q8b4L4MFTqIFGR/eUZV5hzQIF46v7OGXJtQDRrD6z3nXNEVJTghkCVBWDxpvEdEBqblD40P9Oxx9
nJ519RVmIHOPVwhOdeodDLqGfmud5IosIrcMPs30L/O2mvgiKS2nYuf0rVbH8YWmkXess8oUCfnT
SDu5lfCurX1kVp9H68UBeJ34GgA9P9rQ00ZeuYxCfuHtnii939juh5oUp5mZdqbqQWU34GZ0cUAl
9WR0oME7nv7G4jQvZLTUJhR1F6B8po7sGE6zLsKKKh1eqPV1mW9YNf381ACWBmSQBfQhqLeXcUJ/
fWlTNA5nNx6AaFycQzkM5dnF+P5hIy+Ad1/dvc3vsMNEB5iUUO+gXuuMH7dWbTMHroWHR2rASHm0
kNTi5HPbgfg0fiYRwiqL0HDQ4NIRMh6INiTRyNwQ0wy38gKduFeYmA0On+1SQV3cfLsCeSl25Ee5
0d6MN6h0uuUhUMzN90saxsGs4ACVADaYCx/f6aVda9jgDRAun+RLeKw+DTtLL/Akn8UWE5RXlahD
+my/OC66vJR0Qstaf+huPHQVOCN+iaEecYg+Xq+qdBqfzywxQBdz4NBhOVxz8tO9rAXRpL/UNX1c
nFHieB78OasainWYpN2ZMvT2hbaQtcXJr+5yi21NGEzZiiU0ENEm9xH5PxjUa+YQUrXLnhxQ/HiK
EQUq5CjHUMZoIqUSDgsX3EUNVlNDaJw+tq+tsVk4+mQYINzxsZ6iVM/Lw6OgHRuQhZPxFuMQCpkI
wBP6OJD4UxPIcqZY08waO2xCcMPO42QvJj9ZCdml4EbnCC5j394L3+PNR+WrsZtqbumIbiYjVmmt
ePEQaSVZSZ77GhLMC3mz8JHhmK4O+uNZHdT3s9ETsewLE8JD6uPv6yqMqB6juV2qHJhAV+XqnodB
dVgcCJ7DF+3XijH9KiAOYBaKZHLyPMMRl27djIPSvtaoFDedOeHQE+pDZVnNB8Di9hL+ErQtolWI
J10R8/Sg74dd6AwffGDeeauyZwx+bedTbMSIa0DG8YK6xo3CrQwn5fMnkixXhPEFOAhHCqBwZ8Wk
BMRrHRMH7toljsLpjV74ZEEK/JSUApaK94WOrV5NmUuCBxjd81d1R+Ute4A/8pex4Z+n7n3Uhen1
qtdOLf7r2V+e9ToDuY1OrT/Zi0eAfSKkFFOWd3r6jA6T9ftFCx/D0YMEw8e2IwpU2HnvYRcOxv3P
DRsOab3KpNvMzpNv14knHLLaiEd2I+KCtG/2pjseWfob5DCr27Q60IYkLEHtcVxLUCQHu4b51QTd
U25pYYtIouqChhbaxa1tJj4H89HWcJYKkOyzM3WCtKVMq5ba+U2eIkOOIGt1sEF74bvJa64Kpro6
W+zAo56lcCXdBZPupNYeBzrcGsysWXuzfbRaTmRvS2z9RjWuqX4pE5HlczuqH3gYJiWKdeHA2F+x
bXSMg1FUGHSjstDK3yPpP3gWVsWL0C7gep37zBb0rUO9s1tlZk//tD+MeIL/sHb0A+OJ+WJQGMGp
A/m07ETYnVZSZ1eQFr7nJpeeuE+3fAFFZA9JwliSotx2dLtqz44EUjg27msXcDjoRq9RxfACJmLj
mPsijweTptt9rZTi6ouAoIW1ebENBkWDRmxUXLv4IHAG+Dcamc6SwKHvQtF4pnPw8y3ydKsfiCEN
IAS0LcrHy6QplcnIZEELBXKZgCVAHzXeq5aQXH+OY3k1LCr88VSpaX7T3+RIVf4gpOJ5DvWxWIbt
J7muYtfTt+uya/sovw5s0l0haxzm5g2mXDNULwxabKGf5JURwbzQUGFK64uHvWs/UQJShVgrzb9U
d5s8iYJLwIIa/vbiN5luNQMK3G0rvnavm4nqZKl7YbbCgWTJ1GRxrXyOusNkmIlDnTkGiAZOLRQM
8AWY+THHg2m4SEQI9WjEdYRz6Sssi7DbSN47O9XKjRhroNrIVXhBtikJos9BRbbjrs/B6dErDug6
9EPzU2NxDGK1e1KxbdgnNYMAFAkG347hCYm0pkaHNNel6lDZ+mzrhXRDarqym0opBSjbxlz2Sfsp
tzIKyIAkR9WPdDJGqhnfIc3Qyy3v16ctaVeZUwRyJErSccAaeYmA0SLErCopBu8yu+PQpvMgsad8
1tkIENrP5V1wW6s8z/68SqgepxxBhvB1QjzVnVr6gGDWx/52sFvm9+7FwI1RjeRZ3UZHEGlSpe4t
oc2NkvtI4K/0VqXiqeEzJMiE/HOHZhjGWDjZuameTNmFundzXZrDyBWa8I8BBryetZ50nX0HhF1+
GeRWwcfGEUoNNHoluvDWkkI5MBHehoCi74RxWWc531ys+6ow/AccT1ArtcP+R+PW8DhTb/003tFs
6eckTZQICqbILqEBYnkV/eAbt4b51Vl9xy96EOJnayHdTwJjw7VLrXr5vbT2NZ+Y+2F7vDoJD7El
DgoZbmicuFg4viBTFs73pFiLzx/7X9bgfX2lyYSOGxgg6FAlBBTU1wa43RAmQ0bzLhFOdVq+3i8T
+mPcDBFcdbqBJjUzhNwWpAxUPVtwYOZQUhCZ0L+MTALLEt0YnCwWJtDIjn2tJQksXMcQNmw/G/hQ
4zyRhj69YmSstLBgqb05/TuyJGmw+sv1xMYLbplUGjiFjacO4PkdOBwzYvkJI7dbh9YKJypPYXa7
i+LWKtSLFXf5ZiUqggZd3YodBRQNu8aKGWSYCUmswM2HZrw+3DsBIS9CZHK5cI2jBerzgTiSbsfB
xyL0si9mJHY5/3Lg/BtLGtrB4H7RR6pNzRvvGFqrXuYFIFB1i/Zh0swljG0eM9075FSwRxj9dcCY
VQXjWOqvIAszgxDJgLIhVw3857cgu92AINpuycG6nis0QRbootHthsryRo81NOdODgykPubE2wmQ
h3on0gQoKFg9aU0DYTh7Cuw+8OGtXp5oSKDFJEsBGTyn/Bh7hfva1qFN5lc6OXYm+TKnj1xMRFJL
2kw0bovwNKZoAOZtCPt6b9y1Dnw/C9766sKEi0ln7sc8M/pLI2W4CKAcUljVWWM6b6zLv0C6p3F6
VvDncwFrCzo1p+2TPpHSTEu/SYrXrC1guNrVqp8DPjVezWMR29oj8DPHlIHTNaPua4ELf514VBQi
9gfH27EutY7vwGUeGhj9vNkIvMralFbnpwLuhW9puPoIxLnitUIHdgB6x5pds0Du+LD6C2dw2111
UTYb4sWm8LZkqP3ccAS7cG5mtaHWqYt/yST0UAClMlZtaMY8+0FcCpGFo2Q6TVZGvrchaMDIi683
yXyrmo2yS4mm6CTz7OKR6aqYdwzg4Jn1tOPjzxEloUj1ZeMlHEY3S032wTqx+Wzr8pQ+EiW3vm8T
67oP9cGyakKhV6dZSqdki2mlb5D300mi1EUSSmhMR71don0HlpGOtB8jbHd024gw+g1LueRq2+FL
8FXgPlj0lCRy3ejDWDmxqein9sOuYLhnitGsRL2l5TguuJUudk9E75kPWVpe/nhqASs73FCrnkuK
1mIebS2FO+BL8wN+X8SVH1pLUKqU7qqKRiOaMyAHOwyqqNOv7YRQLakQEhm8qy966NdInKniZoDM
xGXTfOopOdS6Lz7FQD9wv6RGio/nEdlbrhfYGnQ0RGYuxDzVUDnxjbReCkD1xwsuz+ukd2o3YWg7
YgPXRp2Eao2PgodZAevkMMfohV0x/zpb63WSl5M6Sz+EexVORQsMWHJplELkUcYScmSjyrmkOEIP
E5FdU09KDoH9oIcQYclKCNPDZdxzEcSVa3Q8aqohzXURfmgNOpJg240Un9tRxw==
`protect end_protected
