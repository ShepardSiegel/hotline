`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hPl+naUBZsqPksP+JeUkb2CpfRXWNFVNzN/o6ZssnWdhaPz/2ejA2/w+SxlpupK9Ywuf+5snfCAO
f5phLb8SYg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pDoORLwTR3Xr8IlQrU+pWQ+vd2A/FYOw7BLmq5PpWVcwaGmLlsttHyYQZJKp33POKZwgNlTQM4Uf
lX+ak08ig41M1gbcKTZ0bjHS8GvrO2sUAKJMbLkF1f+lNTcu3IxOFeClQCMzO8l8XP5Qp7bu5vcL
t1Dp7YQebq/IMHn5iwg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lS1SrtdQOBnrj2oV4YEL9FO1cICe6HblyvzCUIh22WSLvaT5M1NNUFtZqDDcp+7dsjrL+XQcUc9y
Pn+fHMqj1zx3ZW6yudoCIuQY55ywR2CGz3Rihmxwwj7DDt0WxCfBIlMfHbrWMhFopt4zXkdXc6AN
IeQqcJ+uV3Eaqn3NEsG7fO2hN0JaZ0H3IMpRUSxc35OE6CHyYpJAH4NUNVMWrPA9Gy9NtAabN7U4
TJlq36PI7fEaRcrbCOevLwxXyAirjO4v1lO7pzZjI7Opyqgf9FdvGthojoKP4kE+ZxoLSNMHqedE
eqkyWmPqLeJiaSr771wxfwzb88JfwtAr+RQv2w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HsBjDSUld7CHGKAa7SfcfBMQbBpEZ4MQ3bW6xCenI41PC/k8brS/zJF/9IxHG4wORmEpE4qIdrIq
ANcfVDkdYaCJsgQQIJNjKjIJgHBYLzTiPfYvU32dkNYdwcz6BcVflP29E1CWb8U5INsZpHpe2rKs
NIrGyj56SWCr50MfWuY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OCSNH0NOnvZXvDBZjxtFrpxHSDsv7eNmlWasP7+j3rb2z4lY9GplCYQimgfm62h6ll87U3HXSoeg
2l254edbrKSc0GKWEyHVY7TSbN6mgslbMY51gT4224RMcMVbqpQVnCzee49vcGsfDVw8GUGWkSV0
RylXvkFv2de1BzmFTTJhaeaYeRwfmIJfG8oWN0zCUuaWqhQZ8qCBvG7iVAEwjYZsXYZZFIZhGCOr
2pCSq8EQJWUL4BqqNvVl4AOloxbo01shUuv35nIilFnUsVMT1G8fv3sE5uGNxosaK563CzVYQXOM
6YbYuGE421SXgJ/f0cigSCMVvqrqLv4d+vD6Xw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23344)
`protect data_block
mawIyqR/4mr/B772jTIwWzkL68Lb6XthQK+qzdyjWZ4zU0npXj1B2IiKheEjMT2H/QSczoDtFfGo
2JmdpBqgEfe7cjnNV70Zj4Naaz/vx1FvCJLpRKqLEJHeiqkqgMSp2RCE3D9QaYn5lnapGvuJlr58
oSkrVi3lDO/d97eXpi+xh+HuBxdtJXB1Qa8grhGT6XSQ4QmAcRtoomg5WbLXH8shx4UsIH5764fK
fhbHOatwc2op+BPGrIgrem8VsZv3Drjms3VQ6iy1FR5FRh9pKTWa5FjsioupTioKWlFcf0JX36IA
p8M91CyWlXr39yPrgaR+r2PBLzZcDQesfzg8kOt+XLz691287Ki89P2YMl41tcOHjc2fL1LQ7GUM
UR9ujlpPqiabD3JLjIma3uw8sX9XDmaPdHNDjdt7/jPZKiPpB4Az8pEgaFC490EjU2HBq6rWX+VD
8QyfTD6DSo4WgNZmwNswbF01Heioo0Qa2HPJHxpNnRqEw2QnT6+w0qb6oKoyQIb+1gk/2trtpDi4
neCerLlJUCCBd8mMP2v9gzjnlByb+Ylnw1yamIfoZiI3CJ5xvLWnvebKJLjj+EVriyOBR9DrS1PM
HfvfcC35VWD8xF+0Mayjlk7fHqHc6cz/jfVg7XSQlpjuAkK9xxIAhs8e7nyc65yIsEQAn08u6jZj
jJgH6j6hZvPxlsrPfGxKALpWp98y7ToAHJzDy7Bjg5vc3MpC9OR19tOzX0Ij7OybI5ms5TMvHy2o
WRrPMoRofdSlJ8v8+YcUaSTbwWqJoxnXJntbkq+zYNswmHObeIfkcvDRHRY0EeIAhlou9MST8RPR
cLv95PuTW81tGgxgeUEE6Yi6E1bUDI7IaPBRHr95f1ofaeyEIobpG+EVtM4VztddjeanB2XaeXFy
aaysVVQ5J9YVednlWXUZYXMs0btzA1iArj0gaQA8nRP7Q99G/H3GxoDcyrvq8mBtwgZOlRrQvd8Z
OMDgUTdrvHWTEDgT1fNi1JmXtt4n3o+9FTbUjef5ocBYkJb5jgVonsAaGVtlAwpEEwkLn20WHBMl
0ZFOQI57Bk8kfLe1LmO6vFLik0sZmk7Ghhcgf65d0cMnHLs/Fa9ebt0vSm/Ykdsk4o6VZEKRBakJ
cs2pwxJlyyOOrWdBRyUQrLnU/2qigez3kAryTMIj3N28kd9N/9g2Ngs/LzkwsA/c8CRYCNGW4rNW
5rb7hyLp01/zabFpWx+tp2z8k59i5ufdgnvN8yPX3eSJeS8qW3RrG2YFYCy3EC9LUCJnopJ6OHrm
BTwI6V4jMemFemND+gz7B6UXNXu68LgThLYjM8ssKYNNZMN8MSyYNPCRkEe+XGpgl+nnWSHq2y+o
kDM790WKrkTMC9Ocu0EWarpKLckThBjmauLI7bJSl7qKrnu0fclAjk6kffwhkUabbGvI5JqPMHLx
3HS/M9cPr5SQbUlJFDgetStvO0vt8b0Z4omRmVTOlL/DgzuIvuZQiokCxmm10SVFoO+jHa9SEJhD
dsfyLfBCY329TT4AgiY4C5BGn8DHA/z6PPD8tgJp8gihn4roEIt5igHwn3UyjwDv9RytV2phIzJo
G1si+87pFtM1jSRMQW6ylLY8BI7LzilURJ2QAit9JNj/E9jKRstpsup9wCncAy6oI30IPwO5FQI9
tsa8FpBC6ssn7GT440FfEiI7aPiUhsaClTBg75KhM8fmOlL4hP6oIo7avuBMOAsyXfyreWgByi1i
Syp4a5xxQq1tjvfO51ChO5JyMLQ/FaXV6rhmGYljhE9cxH/WTldfRlouTzG6KddwT7DQRiB3gDHE
Dhw0nDeXEubLkiCsr2XNlG4aGj8Lxblb5un6YOfb7GkowNWJgnF5MEBmihESY43hDyexv1aYufRD
hNVdGZX2YylNjcwvK3hpdFRi1oegSYzs0MIJLtj49XgmnH1qQN1fO8spBf7zCKEZBk+VFCVWUhuj
Q5i3eeKciDcKTfcyXomJe8RY6mpsXE8Pm+8rURVizn8L32TJeJuBXDV8xm6lha0ehMISOKteBXgH
Bbs9xJ32tPMLKeuHq2ayi2O+fZ4ye5o7ae2ps4ybo80dGf2+ljAGEVMONwfQYeGq+o+cq/mN1Y2d
9TsV2bYZ2KEjUSIgnQUfSHdcPIk0wIvgNGypd7Y3pybXSbrgnJa/sGFoA0LMAUhDtArOhEIO42ZT
kc6fdPJAQl7RoxVeytSivyM2Ai3ZuVnQmtS2QT4+D7XyFH0L+17G2DSk6k4CwoQ+3aQMutwLUbcb
UddiL2htyyYiiqDjP2YzTgCxk3pLiqDKLQZ09ZyStdLzBiNS/BO0qSsdKrgEZmuWDGY2m6cmkeFS
9trN7763/o7FNWte7RWIV7nqE40G+svD/x3A4GxekuvUX8QCgwbrO12pF+UC3GgHx8RnyWKWuqnN
J0WmVBpVRAxhgOd92y/qrV1y6K83bPqeqiqfP+lPDz+v/YBtOFwtSaPnIFZpkwFIj+Gh/kZoHQd7
f3j0lXzjq5uRkb2ozK2t3Y/MDyql1JYkq/Eq5Ex7P0lO6hvc3w9RT3571/G+bd6XQOc505wc1pdC
5uCvjErd58XTDNSsSokkX9vj2K2mSxXu06Q9H58140Upforf+gFfwsvF64tAWFgmIhXv7eNIdDes
tgBNDgkxO7IIG+ECbgEjBtCWCKNsswjkxzcCG6MZqcdM3ISDGHcN9n8BUHPwMPzoCtjveIX4WkUZ
/hMMJLPNlDRZLj0FW5rvsYGt9dINyfwNTZnte8KyF6x7JJkEZpSl9az02z02Sv0n7Nur66ulM/0S
V/8c59iv5qOSSKO6kY6Yki2OYkgiThy4fw4K8q1rAqWWD4k6j5lpqks8sv/qtiUV4JDTePFnG4XH
FY8TpOCGi4GqAdtS6mvrbw0C2O44KFml0N+B+2Pnq9KT+4jvFvsGKMjwMEMNU1C6EVo6uMlm9ssA
Fj3yF/PERXQJ3WcOwihHim/2BLGynoV9N/ya5gPFDC1dA0v7cavuXgKEOTMPp8Fitx5mCK1mNQjT
dlJ7G4iIF5SaItULxDv8oQbPlwDHij8JKFOmOCgv+8HQCE7PValKPCXwO6EdC5nd+QSNJjl2U6Fq
237erLRINNV13Jd6KK5eWZkML3i/hdV0L0USLZDhaTNoVQp96AbDxkaxgUrubfAdyirCapZa5as9
OWwoKJzMFT1EX8+1/XDc3fIFe+mql/Qo8qz9QVPK20v+RgKlabxdt/7r6TvMDmW2WQ1UfVIj4e+D
66QwSrUdfBuuoMMc0YgVb72xqfn4ws9yh1A/Z3uHOK91R1ebRhZXxftNobXv5I2Gf6lMxdeOHsH3
NhpxC+nvLbvKQFXLsgbN1pKFd+FPeGuRdX6Q+5wGu8qZ5vP6/NjKC1LlyEUAQGvJjvVjKl9vn+dq
l+0aCG6MewIP3SdiquJqJ0got2SL4+gb3uGGFvkezCoyu8vLHFpNzJqn1WI0ZUUbPbR377gwV8J8
Iz51CRVWamR5aqQLMHlZnztgnBW0igNuLfPbvlKKZsdbt7tKGdJlVQwAWTMP/KG2zWMPYgKPdScB
dkA6/0ie8KPnKrXDbNhqp5L0mBVyaFpFa74K7AsovnzVNCzyd8euvx+QNfJz5nlJK/oYYL3HXK68
wq1KCYWxfqHB9mBf2d5U+xVzfCe1XEwnHRnfd2ED2w9v6WAp4XyaGKuQQR3X16W23EIajY5P3idV
4yAVanXD6/t+3IkLUq73+4txjLT1858RLUN6VvQ+ZZn3BmVyyNMAbEJP2EGxau3po1bfaPZCIiwc
IiI3l0HllV+rryaVqlsaizU7KGDtRTQv17TrpybxZSFbZUGo/kdS15+Hswm6OtVk3PXa+peLVXi5
8llxZEFJosOapCXBF6g3SQvzKtRzNommxrjYnkRpk8BATfrY6+RJrKLIu87zNJLexIOs2ogiwG9E
XDIqBgdJErT5pzL4yDRQMHSyyHLEhJ7H7WPH0WVYequzBC08UTDuarlkFyCkN2GPG4MwTn+p/6aS
Z0SZUrsimmPrZQcNxTsTBWV+qQT+gPTzb1s0QPjovm5K/05XKxC3qsFVyblTFaFViTL80lmoCYaq
esci5582E4B7xYxExWYoDzMLM26sL3KVtiz/FiLpbG23YcDg2sYE/lpHPSGC9IWJU/PniVAAzfJr
88M6j7jFU3J9o34lnUmAy5CtkFUU5n1z4XiAnp1PdWetldP81aGctuNC/DnlZmJsa7oFsylebfcX
6WLi+gpTP68M1+u0Rf5MtKP/yOKqX+F4iAUlMK1pjB2Kfl6Og/ZPTqLnBTK64sw2e0K9qkLjAieV
f+uQyWrmcEsH0ZKFT0FbBlQOCoHwQreQC8wsooCfnabnRy5E2yATL+C/mxzGN3n81JLr3SJT1ZSK
NMPpjGBOpIBdzuO+onfCb31wzI16mznCG3+dnD2JFyCMWgodCPVxYfKAFq3lrQngL7hu0HqRWcHZ
D9WzkAm3vbkdweh8aHWkfAg4pIlKHlT9ZKa8TyHNGWGx90noNeL04MkXacbNzBIfzn6JXwilLvqQ
6R0nYQxS7YxlNkgJ1hDfbOPRuyM1Jd6+Xrc9MSNw673wIqJTYiyCpFiXKvMm4RgVaVPLlRHfloHz
xIbWU4FmMn2GSRkXO761X65jcckqMlabN+lRmmMOV69IlUVrMe/8DMDVjgMUg6HXZnegK2BsV5mi
k73IMV4DpWXoXXvaCrQbSS8ypcWTXTsEgWTtiHfVLGEDzP/QLDd5wDitx0yiLldamkGJM5iV+Llm
buVybkqUgXITebcD7FYz/pWpvIf4wo5bNvvNKV7D+ktIjhOPZKvSflOwZXEPPKrrunwYjJJ9+ZUD
ly3Atjde2hWfQYIpLD/KH+3x7HL3fGpMvw1wBpYw6IfjZfNnXwitWrj5zYwELwrq9psqeDhESL5O
V2RGZWq4aV81dx1RJkMfbByNqw09VqgR3+sxXK5LneI7yUlw7TDpDwQJPwYE0Mtx7e5AJoGHX3tF
kAwXSklg5QK1ue+EGVDqMbeaLFD9R86ZanmTdmeTPO/MksMax1P5dhlihCFaBv/ub0MPrKWkrooi
V7AQ89thj4bozL3B0izaoU/WLtfUNVdrv/pMOWYVGYAokdMYbJMRR1Bdg7URax0J/uqS1J7vLaTJ
meAbNgBRTMoZ7+sS+OnjiRuVC6RS46teRT0vEQ8wyOdWjQ0I3RAF1iE/bFrCxxtM5+5mtTsQy8aR
1Rq+idd9VV5lhkBpDUEfoCF+PrSnmFzwUwZP65uoWfsTw1H2M+b9kiuDCPramSs1zHQFcBedcBNU
p3aAgzmHQntVrn3Gy/rad51/a2zMomv6RVRUO37ZY4NYnleWHIa2V0AAQs62trv5whNOPYqfuMyU
6tYtIQZ2JRxqb1oNhFAb/p97PTi6K7cuaFsvAUd452gaPwF76b2EM04XQJXpESPVYEv5RlDT5+RL
RsjcGqj50liATghnnAIZCHXyn4xSOOPkpGK8GqG8jDHOpe6fOrwXcW4eYU/R2hVH+vqHxGFtH38Q
L7x6AVNu5ziYb1zrUkBk83E6TFJPjf68A3xe8WBf2LL0e4eGHbag0VkTF+G0dVkYCVkcuuxVDlZr
At0r6CxmKtupE069iAhwCVd7FpoEjYCw1UkBUjCIDB0WZn2D0KfK9/xFhzpgEVr7j++02vx0KExI
IoWh0gVCq00ysqcUgyDcfpakgJb7hIIFiujmlDxY5NYBaYdAYZAJfYdApSgfR8ReAwvuXLa8kIB5
wa+YHYa4ObWJTEWE3pFyZpJiJ40vKM1B1G0002j9X8LnNsuYW+MJKytDrx1ZNiKNTLTZkMtO4ANV
R/JUgzs3MB+QpYLrL2zRfIn5UcChpJ7CkJkhd4BSxZlxJpsOFfz8r+cz0ixlxKVNQlbveYl5Vo85
4mV/xGO+Aac7dWBYYszB7/54X0/NCrhbF177S/i4Rh6xY2op21muB1sOWFUeexNOyAuiRxNhXD0c
ZP+WAU00z5SA60mlbaW8cV+6e4HXsLUAoz3zNmm8xdpItRju+6YxXw8tY5swhh+mTm+TMSrLQrcl
E0Oac8waAShXPVBmvzbhRebcooom7OaBOHV6fJtkwU3KS4iv2oVj1EY2uoUjsYfVTdth1kPrljvm
3TmphQJ14IUqbZ6TqtXgzVLWQZBuy6oN8sbByGlKPOoZzff1ecK5nhyTan0TjzX7JRG+/mJ+Szfc
3lmUmo/A7/LBdOzPtJ+dXQjmUQzcwlMq1Y90MW4uEhf5u928iAjpU/MWrZzbxDy6GQX9l5GHeN54
zxGRAhY+G2O5MH/HHhNu0IaddmzOaQZHqTs7Qj+X3Ogy8bkfaTmmTePXgSOFRRY7Tt6tQ9S5qBJ7
6zRo8h3jpjYmf2tRbHQLxgt3yJoBDBxOgjBvyxT09hqEzNqe+xuUAlK4ssbGREvVCjnmR2GxIboy
LhFkkjDpr/fa3JnjoAXnGBGk+A8Q54lwh5azifVfZcp0q8UFxg6m0dDOVqcV1pT9oBrOorwLl9b4
uBevWM/+Nv+beTE/g2Wkm7Vdq5J6cQuwMMxF/SViwXdPABxwJJxhPhSrldBINUGKgrg3oFE4HJCL
ItdD4KcQLGGIiEECb/L8VTpM+Utk/6OVg5W0Wzm9AEwaR4LZLz+TtIVe/e3X2FDJnRJeAFloDY6z
NcipRjhd7Iy51oqwp8DrzQBtpqowP4PoZLCvBOAmYRZltE6ZLTXDJzgHgyhDfQlpSmVMh4PeroQc
Jx67mdKcrm5YtMau2jz3BEduuFK8iY3uGEa3/ptddX026PY6yX5EILMBaLDdFZWh9Yw0A7rJwpuI
QD6tAhROFxu0Q8pHZt3XKOW2WmJZ/AeIS0KhFzkx+ZkVut8pBTvVPMNfBwLW/YdSej7DfW/WcoEA
IkZN8qCS/bEEN54kaDqyikHQNvbFUQRRetwfTzSeSz6qwRjSSR5FB2qBXIhM0ax+O18FCVKbyidn
lURSNfBNDtPPGWynXf/bKToqR52/86BuaBcbtSsX1dLgXkmXNMe2QAblc0BsYaccLtJt9yc26IFc
/ZD+cpsm/yMvL2mdBUGLI5zpSPrPnZtr72ANDm1VhEcg+LlBG3hed4cqLJrF58mncVLa1Sp5iDfV
to7VTG2zdUdsS4xKfiYkCnkESQoPW2Fqy/ba0jiOGbKgEGXlhJAdftso31VjU5PPsi/CdxBiIVlP
O1UfQoy6g3YDsnW3i2L6iY+OxZvdfXMiARXsIiZxwkkHyulv9Qu+12rthhqcIKmu286Dhsn2DP5N
FaHzi5I4AxutArXo+CCNZQA15FpD8xCzeGe8DX59bg+wAYnz34k4lmbuNglDRS38B0w16jcsqTIx
fdmszRnjACl+W080CKSzgj4nJEnrOnR3Qh4XVtvcNp8AOuhVAAtMlixOh/PhfUZcqeS+KZBbMwky
SmAdiaIbjJPGL58i4p13P6wDnOGKwrmJUZPn1ncjFUKxQgfQV+4oqcyhNjbrRSlKUz/S8+nEDhEw
WoF+xDszw24uR/k47NVCOLRdeFyYfWa3RkguOVoKjvO7tRswWsFTw/3K0UvLiY1uEcWbXxGrZBHj
JFXrVc753WUWHZTGbUcs/isO7J+M834sSC5Ey+lxpXyoeZWKTv/rNyPTq893TOtYKmQzassCBTpm
hfuPtXxVMhp7XIxx1HqnQIeI5+8qVdWzxh2RfMrI1QCIAvk+dhS2jWHdd2nMdpO1/XkEZtdtn30u
ModP+9NUs3AyjmdtTJcveGUWYSIBosTbMujY7+dl6Q1bqV9MK2+I96aK4C0BWesz17iUrykQMqds
JBlEGyUE25wI70shht6wmScak4Zarngi4xpSfduByYeONdvuxU1cLugKtdWjKH9s8OzsRryvWnjw
Yp1VNe4H2UT3MkmpFpAuc4HDUuIvMMi4LEyogcUpFGC9lLVgvxEkgzBmwctMJBXh4JgB0LFO3QG9
/Y/lqzP15KDqXv+esko5ZzVbBgQO4eQOMW6xUHOr+SfJNNHTzI+SpvNaCIWLusXxc9viYKwrnN+p
9yJWT0ZdZxtjQGfXd5rIlzGEl7M91HocYmF/r/LjELMecdwVdj9WTWdUEeJq9EhPlE6GileC8J84
4TqA2O1maLEmUT4ON9R5UA7EjUmNX2BgK2eEh+fFsVibaeJCXt6QpPzfZPBOEjtR4VxPftpMUshV
EgdnxMA7fimlxidOCDbhgzE9OTJBUiTqv/Ds6Fj3ryZuAKE6vww/L0sICkaV8+SRIuDeOqy1SElt
RrocGwzTsn6Xk19mwRCSncDPiCgTlYxGaOPgvJ6QVa5F4To+9rIglNlA4yPll7tnSpXabOKsYVFL
b76joVrPnd5ZoPEFZhZQIk/Uyb3lvPgiDm693nsqp8mazAdjdNa3PzmQyVIqB4PDU4r4M3C8wvWc
ZFBzRHvZdDt2/irQGZsOeQoRuI+571S/QTa7yD37zDaFWDGP2xmxx34n400Ik5SQNYNgkrg2OHUG
38FtAz9F+1tcy81UlArjok1GGkEdv66SF/z0ENGgbqlvgxloyjXpFs9ydOolZ+V2/AXIBYThMT3u
0RG86mVHp51GGX6zfhVxJLUGpA8C1E4k5tuFbYBWSKWiUwWC5oI2Pppya+p/7xsy0ZDxUaRwdFq2
mp9znrzhjWdhBrZ5SPVQXBhmQXflvUsTLPx2BMifld6bb9dp54LxwOjf9555iOm7EV7RXtmasmEb
ZJKzaUbwXpl7HDLc9PQfb4gFWDA0Blv5ietWLuxCGb8qHTazBMN0aAz4WZ5LLdEGZWy12iBAUETu
LL1QfnOcTioGV7bWxhViKKpzgBnY/cpjrWmV1FPaaX1nE2u5zZ1eWlTyy5ClepfJEJHWFERCI8Qr
ibnU6deKNMnbA6X/t+wXNKZXR9y9gHSAfVtxadaOb7jYp2yEIPL/TX2oT5nGgxOkbf3EBaknw+dc
MLoK+SEzbM7wVQtuMASvm9B9I7TMPXnG/d3voC4yv6sfUNhiT9CFNEMlIuMnKwLr3NjnXf7umxdX
VLEEO8t6aPLxbiL/uQHJdbVQkRdh9ku93RPP/Ak50abxvFlKmvS4UgyLdz8VxPeZFeHbQqiLglFq
fGSAyqgSRVrvkMu3NFWodEMWKwOPbTmJDmPrr0X9MFeY8daPZzP9FkB0hijt+RCGnGSlNPtz+z1A
T/97zarc8nVdz6veqyvvCI55pf8aO+bg4e0OPwkoB5bnOMPZ+5McUsT4n+B6+nC43tr07E5A4flN
JvKXFfBcjUVLb0JENoKuMnXnfT9SBPG/CsvtlE70Ng30G7k+OjeQU5YXhUd/R8XfzBbpdqrFCPKn
khnbcm3YhmbOBsQZURCgdzfglURQKhLXqb2HMJ7VQyk8ifsbgfsyHxsrQC2HFjKMAjYAI4SVcbtx
+VErCPn+Jx350kHsstY70y7gyHk1FZfAgKqrDTIfWw2lJwmJAgcWQQlvgEt+tmd4Xj8TTN1rGjlR
zLkt/Ystn3uFzJxFuzX+u+vyNzTgkl5zaNNgVycRu3POIBexD4T7tuEPdjLJjkQJipYrkL053WJ2
VhEMGH1WzdnS39ldotiztzwVExRRC0t6FRXThBSBgV522RUfwwo/+Z9eJGJFkqU1TyIvlxPc1fQo
3mJubZcOF5UaMx1XhAIFkEkkGqoownnF8wAm3VmlVyj4uNYzzhWHGWotNbVGMfitfrCc5GA3KkOZ
1IllHbj5g8feq4lLJGufbDYnNr0Yif/+cS4h3O/soID6hqei+zHhD7NT+ehEFEqRfKWnT8hVePx8
PKb0aaRRpzsMy9pYgq/51aI/2ADs8j0Df7b+Gd9jBmGIyOlgVR3hSmRFkKnq1g7NW+1kQf1J0Od5
BUAAb5xveOlBe+LhGfn46SF6VKdGAPuyVxoELZuVpTnu/J+BMZ752DYf8HyL8G8IYjrl6jx4AdPF
F6aLObbQ/PCHAYjVNLxuEvWie4mYIv43li55ze2waUwLMGrOK7vr9pxrFgtEe+12gQM/u8Sqg9vF
ioudT967RQoiBwa2cOE1J5HzrPqlDqIoszF+7hJgjfUlHmMDw/Q9IK2c46viAznFFFE/DVbtr+xS
XTF31Z+HbkN8lZ4erKXaVxTjVpfH+q2Zt6ZBNUUoPO9BytoX0HfL8hMmnfyKDXqjfY6nUHVt59cw
addCky40xtMALnP4+1wT6CdK+doscZRwVrhLnbfRNLPOJWkmxQHHEoa+hTqa3pPHjt/T369UQ+5i
LOvR0EorWIxaymz4SozfKaUpEi1hnQh+8V4aO4KCFmOkeIG5H7nqmmMKZ/SINZPjg5+wfqDDfETo
3daoW7kgsLBPxYXgr0BChpARZpXSxkw98gwBkKDPswQ4rReRTLHnN1YfPqRtEPvjbsxUd+KS6J2S
ifky1ZfKjDOC6vdLHNz0Cuxvz11fxCLEMjCcR+qHe4BzUXed5Qjpylb9FoUY1l4tRVJBoE102CXw
pHxTh5SZ0pZJvglUibnw8MNZPv1wVQ9pQKlrOrgXWSf3ZlluYEl/aM70vyhV1I/9ZF0LjAIrRNSM
v/0miwK2sGoFWw4nkF2wtgJW1RtFeMsb2Z3EJgMmP0dLPKrXQYXJ9L7UklZIQ131SVvbx7xyKq13
UtiGcBfo9AHor3P0NZ/4q9FLbzsH3hf83mGthHD0ONa3+qpLo5dGAWhzRbrcK7j1flkkd6p2R/aY
FvYSKcjfE9QowjO5fZWbEyIcsez/t9SdQivd9UARmLMM7dQgA4uAmBcQtLGOkvoS/idIVUB6Jf3u
ht59IXD8cTTq7n1qpgQf58GLSQrka/BjgyM3u85PnoEdiyD2/89YNT/U5g+Od1EZZzTebC8/kUc6
UjHr+r9hqdMVCaSZOQwHBvsnuWdqU2wiKEN+l3lRVi6RsdINQ7Q/xC7JJ3pmTOps4/6dBChlLg5E
FnZYcLujqMpNePtfiw8YPzTHKLdydZxm61zugdhex9yc/nzhU+9KpmZMcydAmLUlOuZ/z3A7s34u
PlGbWxRuFquh7IWgbT0PX7FVWqoqNEPJCQMY7bIyLqiA46ZWV02Opz+mosrBk7zY0N+qk3qn17/6
xv7ZgFZPkhqDZEzZzMJBu/Ur4K9X8spxdVvcu3qXoNDh3GlfkVljYC/pRgi79Yae8hIJzsU0Nfvw
sq7XBxkIp7QfoIv+wDM7AA+23mOx68dHqKRRiA/qSM773gqA82NR0ussZRNvIVOlCsFZNXNvC7W5
NbnJ1RPKr6+iLMWT5zZrm/khmgX9r1vc+TB7JyNpHHnVKd4m+ek71UBwWWaNbYN1iy6+5a3zdsNd
KJL4VyisufwnDD3b1Ow4kMH4RYb6M2CzmqJ5gRk4ZTOI+gwze3nLkU833LC9S8c+SDMlxD5dSBw/
PhsP/W7QcsqLp+psraV5kZTKUZk+xc+IhBi1DmQYm3tpqTXnvYh2hCZVkwlWNyIoGTZx2rnEjowT
R63wbWqnMWomHskADV/y6PRdMBcogRbg5+OnnbpoJArGfOkCiYCXhCjZ0ePz7j71y/7Hi9xFZrnX
82fXQerGuWtTIR1us4u1auKW3YmCe0xBolOp4HMSHs1XKF169s8LZ7m8o5xs72jDpHZWens+5FXK
+imcoxv4C98GSht2o5/Lsac5SGKjtkQVEeR6gkBGBQu4qKD06KaX0aYWmisxmVpirwJwuHK4dfmu
OJN8d+sb/4F7pDe5C3VyvrHzpheeK29aQuau9TPOeuFkl+u0FxwTZDjXMKwfZQpi4jY3f3VjcYd6
JFDmVYLZKia9AoM5fi/RLmxS8CaLbcvTAhZ+UlQMQufFUVZWK+x4jaHGHcxfwcn1wvt0cPjwz+ws
r7C1YghBlv+f7br4yhvt6vuECfqi09WdrPbFWDkYo1xzQnj9qqn5aK33EReg1OjI+WXIcbgzPt8U
QsEaGLJ2KuusKNzlL2Mn1c/srqTItSgL/0H73t1GMlE0YUyJCTM1t4CdeG7TgLuI7OS8jrz+u4OF
bGCiPrXBkqmH9UCJ97j86kQp9I1V0CbPnL8B7FNBkXnj7hhIEXa/uKwy6XzCpjgnrnHQe0Ls8ASa
leZEvb5+7+Uh62jQlZYF1von7Kpzd+KvpkILP89UJdEo8zQtTur1PJD/dDGDif17Fm3RpcPVh1Gx
KdYwSfO0m85V6dExfbYNCy2DPEZqPCLKpTdWeIS+vElsX68ULM1JVe2KbSVrGE0R2JWLr8MePAie
kZu2nx219IVFCZaqgxzBAkYMHXg3a9gj1dKBI0xfFMfrZCYQaS0WImDuAQ06yzEoiFYUgQeIS5M7
VNJ5hj32MKTAA6jI8x3wg0pr2OOQLTvAeb0S6++3j+QbWro3YFs656X7gxLLvtNBOpM4YBmmcn4p
y/zXoHz9yeurK/dblzIPMLFHDRdO/G+GTV1P+b7ZWNALDy2hYz5/jYD5HZr6P/8scsRmBwQseJul
IEa4eZzKSK6DxmRxoebOe4EvH1nF2Q3pIMD5STOSFES2GFJQaR5vlytwsJ6YZ7EjpS5ED4VNnRjN
CfZDStMM8QhhMeBvJa8udJkQROJuyUqcUZfaE482f8b0RUF2MbXKNJY4vh8g+0s/JczwDLsz9JNx
AWqPN2j3I2fCJZ+fqZ6fx9W7ul90zzxTJUtWntHVcYW9vOs+ED7dVT8BtfMUreSrOm5B7KU/5ITk
A7bAAFbDE58gFKWzr7JrZwsuU46B3XRAfNWDqL4XYlo9xWQeLbkqYUCtZrpLqWj8f0BsF31HNkVT
xLVGd0kkb1bm4u3+rtjzcWONudG+kj1ZV4MdVkUIKg8fwVKP/o61f75b0y1MfdiPnnSrIn81J2dR
/s5Up61bYRX9ZyMhX1mkIutkPxPHPf1u7nrGn+itu01knbGIOIZ9zXbPtM1LKv1Ol0J/LfjFc5Be
dfEoTE5B8KzXYHv5hEkK+ZRLZynvbpGEycWGuQoDAqUQzy/Ph/7tKzoaYGF+9F2Im+ZrwfbxCeFi
26lYmdTa41jLK5DIpYCh+eDpsq+0jWcf+11YM1u6nbFbuklmyLmXz1Fczbf8yLklGfI5ZolAmxye
dpAOSq60Gfzwdu7vGMnqJaDXMAmuyXshEZgYF7PhNJYRxA5IODAg6PsnQxZoYPJcD36NOSQ94KOw
leoCy5hc2OHJ23yFAAdjl+QZrO1YMqMSvKGipqz6oHKcjcIrOPIxSO8PDm9HxMIrULDUbqnkGAvW
+RZ+N6xDtyEUUO6k6DucTjStpxHmZTRyjQXtV8pLtF6b7pIpMv0qqBYPB4K4TNpF53/f6xZiYSII
SZCxU9zD9Eccz+GX1CVJhu4Jg4pNg5zWnk4Az1RQI7uEMRLrYNhDazfemU2JkQuVCZ7c3tN+RLRM
XCELv9Tdx1fXR8ccG8VTO6KXGTKxTyhCx66/1Kt+S0FFczTEOWFlse1loMUNZdufB8cQg7nDhLll
VBQRiYjccPLxx7nFgtYUsx41vnBiSfG/hy4IuESmPjlIiiDTLAY1vIQiaY5s3fJRQ3QAk6PcrmSF
zeepIPEtY5jNlCPhesK1LvYXu9U0iSws9UVKkfh4UI5CN+ljYCFlFFX0Ufx2LBYjs5yBKlq3q+O7
OPGijK4bQndoG86s4fYJSj1A/ZCK5N6o8435APpSWA6DULnhHJfganCkHM7YTevTcf00aDR1hV4C
oNMCcMoGEe5EZkC+m3p+OoHA9kQaqJbz2GUFcOgHeS90BrhrCQLHR3rgRG0q6AAkP5UJn3UsyXPN
ccA0szSrcTkdeQKMxQ0yMQwicUfAR8zUXjbZOB34J2CsNOWamIkYfH62Ijn/dMgnrYQWQhr+OYBp
9VWYm75CnYwJhQG4zBfz9LPO612PJIfOKNNAdidb3d18jAzPdsvBCNXgIXm2ZSe/UmrjOOezqBe0
/YH17GThLQFrjva5eylLW2MwyL12ztKP4uB3xXiuT2VU1NAhrRRiT3IARLy6VvDisQZjVl9ZEUx/
FNpN+78/4Nbz5qK3EymW40Kzp5r3V05xmxpNC7cc5T3e1LUcvFVEg4JQ8+9HxuXssGI7wHJo7N2e
KGypr9rFaU6s1q86oJmM6b4q+DVVJWWcFjc/kaPYE2gWBkmL7XtBtERjypV9xzMusXuVh6fKVs5+
XQSMGxhWnDVfB0TwDub6NjLXlNL2KpbaocGFHGPbqDkW/LJhlIKJsTvP1OStxdQThES4SeluGQfI
fIDCop/EcCr0A3io5Z3vGKXkQ4bfELQ8E6HX+/FAEau0nIwApEu531YQqC+efjAiDD5HAEwy9XNT
DDCNQLzlsSJG4Eu4xuzU80H26R9rhrZMLSzEtZDbcq9+zsI52eyhezqb82FHs5krrM+QZ2wl8/LN
wPqd8n1O1zZ2BpXRRVDw6yxJC/PpxA6cRzXuZKTowEeIT5hRkS1Z8nx2tF0uSLkSve+DukmKZgGq
KvdeHewB/Z2kpNzCa1ffCC+TqsMpHuRohBii8vdLbK2wWH+t1Qdr5H4wWaF0tiSJ1tIEOR1G2zS9
Tr4MDmPlZhzxi9V8ZOBpaig7306CDz0vKyRTxyXMm+y25DlqWwWsMgcoYKN39KOTF5K53LPa3BpF
Wh+7cnc+hoowHKL3gzF64H3b5DaR8fkhzbXtFQvZoyG+OeGsy1SuY4P8x1wwg0IRXgRIjOMjIpHK
cHFvHOOicmypzy+Vq/RpVTFlCZ+i2z7YNjxjbfo8E+ez9T8M7oESHtUOq4CICcFFsZKrIyBmN+7i
wBOaTWdNM4GRi9FVfL1v2V15WylDalrNzA6bXi1YhoGHtzT7h9w5Rv5bhN1yJzFhVM2HyWNVxdJ6
w+sN2mZUs4rdkK2WYW3WVaF4vlyqaK7WlXI0uzqE2NtSnLpyB+f0+QA3j4CRg6ucLuPMDXrY7T7z
y/u9dqNFGZv41iJcqymFQjKWDz21AYf2hZesGjEWzHq9E43PLYOd2mKPdCDFvI04qQDp2IhOkcZa
hwrqIMezxQ806p+WdD2j+qNWdyMsGR2ZCZ8rR6SPdjpViWww+ovBsZOoHdr0aJBMjPXLO5sHXUDd
bsRNUJM6HqpeR3693I+ozjvDC3fEqTwPCsGx2KvdYxrjk89LjQ1/wXZBvkKe7/JbPe79OVp/2/JW
xq2kLoKrhTvjamSK7FntYRBio8Gguo57aPkFrjCi8quYFZa5p94VmpmCrnLHxyVeOSpA5Wv10VR2
j4tvkPsGn3+dRfujXyAKrX3k8VRBZAoqLIj80XX+T1K5g3761tbZH5qEUi6wY9pRV4atmnZgZfSz
AxrBdUwGFt79R5Rr9Huc97C2bfWL9ZLMG66LzfsUVzeuJtLTqCzsNd7LoHqS1Vkh/+8B2PPQ0yJc
BvBGc0Ettt9Kj60upEkHFNqpInEyCzC912pSQ+rtunUrQAXo72Qtvf9jgbQAtVbqoccWbrJWva04
ibn/6JtYVjh54sh5UauthIcZ8IvjmbgrS2mx+x3O/WNuOaqqjKemRocPaLxl9c7PhVIoM0gHMcRn
zzgw1908848Jwna8CSmMKWnTnz63ZBFHuud9X2/ASDHFPFZ7Qh8DWe+KTjAitP6tlDlvLXGpRwEv
WLxV2rFaV32hw4BQVy2xwWRe6ba10D4erlNXrL3nB8XlWVOr+vhOVSq72Zx5g3pcWNGJn6OUpMF9
+sbLz3HQLmtaMEWMW6MKKleKAj9LodN3mQMftO9QM5D6rDzi419oPUpXxVeQfETKLxqdk61rIoiY
Q1zkBx9Duz2ZwMOT98/xVikwYgirAbdNf9L7Yd6HPK3G0NqqW9WZ9tPk+IPrF49jKSathJD2uFBE
8zZH4u5gj6kPp3CCBuh/DE/HZZFJ0w36nNMgaqi+bsfGpl9l1/cFJoFsdCgba096xfaXM1fMeptR
vp6iqGkw5gokpPq2TXURkxbVSCW8tpCyPLLtdhvqxEB1puCwatZwj2UAoFZHhuPIvVHp3d84D4Fx
7czqvLmmA2VOxRcFDlyo0TjQjK30AHz7AXI4LIl1yg6ZUkElBlNasOx6xu9KjuNftyE0OBw1xbpF
QknpGMyttwszClIaKdsVDXqfB1gkVbnuayW30K2qfh4no6kRU0ELLuQ8esCIP5YDLxAD/nRPTMwF
boE5mae7/Fvfq0Tp/2F3f4+c6b9tnkIupOPu3LJfju0MTZKNG5yQkiZslaQLACymVrmI4NjMX+cn
RpCVUn0Lz/zlz+UVwgvQhD9VaUCB2oH6eX20jK2Ca1Q9fdwgfI/F0+mcmLXylpwIZGkofJN99Jad
3XJ3mNDnmG9TCDpcNGNkcRJ34iY0jlRNwmtoyHjekdM1gOvnp8IVkiO14tOHva6b2vFEB4GR4Njc
I/EWV92SKqIKpWzAl7z3GmJA19RqgSa/esKeBR5+zQckuEDVjjIpbvQHOy6K8n9BQJN52MWy1pPy
KcLe7QhKwSNv/nFCejuJ6XJuQosRhbxxJ6mwgVbbXDCqwCq3ZWVI8PWnqHJSJMaM17Q8c7ah4Dvt
P5BVmgqJ5HyMCr3NR2N0z+i2jDZNtxcrJ++MlzsBkdOn6rOpyjmywpyDApu6HTjx3nJjr3FPkM37
cu3KbDVZC9s0eHsg6CWw2iBMOXEaBZ9LhReLbw9eXNJ45fvRAWwRpZjhHShy56FM1hU8SJXd3NT6
dz4zI63hBSatPc9ZHTXEL9GUBN1aQRfLfTV11H4n24zH5GfvRx3vGrHF/JRgoSKHRyRWVlt9A63N
N7aVF75a7hJ6ED3+vxA4u9saCIVyVrk1bNHqTuwt8oyl9Z2y6/tkpVw0TL1Q+G3z29Od5uNp/Vw2
SWtcZoXMyybDFLBRfYO+ZvpESM/tQr72alsb/zFc624wti1W3AJnG3eGelVMh2GCeajTNDM/nnQd
REm4e+aE2U4t2L44iSmWT9RCOuCjrcnR0zJAI6IU5Jie4Wlb5Z77iDPnXimSt2kVqPdlVXKQDWAj
PqKqU3XqNAj9ddWIqiJ/jE8Q2zBtN9h9WUm3GXOqJqip7jaDTgyJkoCpRuyPnunT+zsaPnlThH/c
prdPTN0GrgTy1vddu8WKf1thEMTpX+Pt/odbAy9rAefbEhFtxLdu0HMCJZ1q3Fc5g8pFsjvBTxZl
w9/eQnUEj6+Qw7EDQaNviSFgxakmO2T74/HtFSypPzRUQzEWKi/7x4ww7Qy2jWpOWxsYs3gavUYt
QmY3BNe40CwQi3c2lt1QwnJc1X23XITPfVUfG99AVIkc0IOamrtMev1wcqC9YCRT5hVgOQaLh6sc
YWN3z6BO8Vtm7HkKCUwC/uSVyzKLHkYa9n3g7ceVyfACdSoMPRBt1P8LuyAn045wAOWjyX+RNDy/
xXGoaLOdfQZBOB43LCKe3TDUdO+4xwRDzuFRkbjjpAzgZc+4GaZufQ22GnHzfLLOztwogsT68d/R
NdJN3eMFzi2tqrrmeHyv8zzig6dh9bfffJIhzRUpWIsvwUioZ7pVXhfdfET663J8ijSJV2de8q1S
Y34EBByulx+XmofhTOsbwBQ88Ixnoz+RxK6w5NKH2ZgKgEv9vmKQhQ5uGwrWGy5gNuCvqBM+/h1L
EAfktIGyLvcLrhdgidJjlPzzELwnrkWDRHSIrakVMZfSJoaevnDd5rs7ZKSCtCfhzgUPblz+8Lq3
60HisdzLs57ggC7d4cbrwTREwWVUkHY+klrcTL0Pveo3i1EE36RxcL+w2dBwfKSmPqfJIEziF/nC
xEDNb2v+mv5ZzsXDBuq905uo8HTbnQQ7RRjKGLhl+EET0W3h/hdqkJfr+P11rtKJEfrYrwVOi9AC
NwK8x/ZQdJhFCKgZJmX078kzDoX9kOnqO2LI671scRH8cuO3VtbhnvyfhReqzdtfRSKTod1E6U0T
s6BPziIdsWreal/vgcsUxmgxCC4SngFvEd6IkVeOJ/WN/Qiyan223ikCicmu0jMzghJYpBKdFwMX
ds0obxPA4QGcEOTNGcPgf70ldBX3BXjE1TnatusOcmcyG7mb5/WFP+WCodN4jGTI7tl//PpDx7Sy
F9N2bqoHAAWjCPLVJxgBcCK6eJXLfyza1eKK5960jfrnjtWFs8OxBWuDG0JAtEIYKd2ShYgHQMYa
CM4keWlo5gLYlUJ9me0jhkgY4Ej6SnPiqiM8t9p/mPpN5k836836bv25zfqk4QNk8LEAgUE6p8Uh
OVOlnxtMjRtoR9xZQgnm1UhekN5syTVZ50XkRD4Uu3h8LD841pOjI14lj9L2zmaiq+EMug7/nFFy
18Jwzphg049WWnALJ/y/jn+nQ7AbVs5mjiFYGxEWH/XzWXMuDQYxz0PW9hSYI268RsNZ8Ang2eOV
GZXj81mcx19SGnphP1S2gzD6w6A9aZLFVjd18fhUBq+/0Qx3Z7PxeCDx0nHBt+IGYsvnQIjaWoKf
Y13OEWp3K9YZUA3vdM5A5Ko8wpUH8vAdksIr46s2pOl9xIfSdbYhNbIKLoaL4rX2wRQJX3D4wA1N
oPfkQCcxlPjkHGy4sRgm4fzZrIqYVpcX/tOTxqnlFC9Yypi/fUEUR40vkYsoMF3P+LKv7oGVEYHf
xsVUkcIIAXxR+7hbDgHHofA7Hq/Ko1dhMJgLOrXeMGXKaZaFpaD1boKNH/tGqk3YYoOWHxcM4q3V
Cq+ZSA/pdZ/2nlwE+sL4C2MmCx6j/u041os7NBKpk34MbWrLwxjD8Pbb2yDdrVa+FDHotnO3+69H
w43NaqZHDtSUoFuxsImewXeR8hEqKjjbG/eoHDmUpBwy+9RaCplEo3msYiROyfzJz33bURGPaA1r
isgm7RfT5Tow4EzrywfYXn1dwNfA3iTcRl+aWh1Wt6teFFcIQli2/mPndO6Ku1JLx80JqgJJ1z98
NaAerg0TdByD2Xk/NFHKTyuzizp/9xIGv0k37kGAAK5ENapMixxLVLzOsRHZkdd22sc7tQh+XiC1
rUxJk6qcyq+lczlUHnm38iEyKW4ez/URaTYrgwbtYlsznFnA5nYFcIU5ZbXBRFj2pxferLAhKrOH
pO/x02kH+Zs3U71jw1UeqqIxz7VBP4mIKHptDG6mM+D7JHa9CoV3rjUC/9TzebUmcYF3Vg1hpLxW
hJXrzZJTCCh7d7Cq55SgbS2g6n/UGx+31RYZtgL90uTskmkJYUk00n1dyarjznHuHPf8fvHUcx4r
IeJwdL+dtuU9P/CoctF/CXKNvbgUtrtozmr/MiiqVoaX+4z7PuXguZO9NEis8giw6EmmG7ivpBrj
1izBhcheWWuEAeU3iQC7T1DX0WzlzwVZ94rD2BdASFR42ZKC7OyfajMA1Uu7dnsP7kpFDnR3yvlB
b8KraeRe1DMnCAlvO/RX7m2skB3mWUQE9mnkEDAQJ4jvDLFwLw01VH4B6Fq/9DySOq9RIzwFItxz
5UGeEhrGX+/p3T7WixQz0Uq8lEXjgFAynTxAl9DAeiPpdqcwMfkJmHuAAjnnRgKw9MldqbFM2n53
B9P2DcL94c1rScR56Lr1AJyrVOb88/lTcJfPfkuTqzC0Jq5f5OgCopq6WxrJkAoLHMQ7sk7uBZP+
ihZEzpyORZqo0/w9dkgdAt6TKDLsMNRGD9W7IVivsOroMszREw6IMpzJTFC9l4eezB+/qbME4fO0
GGspdOjb/3ue6WkOumT6nWrkUVTGGogu5SIm0uhYbNDVgohPHQOSj2nLAFWiC3g5K//MOAHUH6Wk
bavl2AQHvD7HQ73KVgmROJWxR7SQCSmGzMJHrXpyXIRulB5m/yYnXpwPoQBJpOSL9VjoQOiVJlXU
cIpynNljj/9uKMPHyeFXfQjZTAgIx+D/nHk46jjd9XsCSsjzzVmOwfQ9wQ4nSLYD4tdUdtVNpHTH
2ZFyLfZYmvoExs8P+H9hFMGfMrkPwfiY16JSSCixkUJcaI6I/NRIMgB+ue3OyC+v9eSZKZreBysj
+1xJH2RhwPl7m6BdVkix3vPCnpJrOgAYQCFXaCsPlpRFMRpF7/QuQRbJLvqkBGqaKQmvfPUec/xS
Jy/pm7JMn2zGjVZKvLMhEooD9stPkcVde0B+4IDtCxUqDUWyWF41F/gQyo1IwjYHEPTBDq3mxIit
C8nrfJN4el16pfn++Xbn/C8hwiGM+UQMVsKamclVT7YlezUwqgVtkuJPvUv1HRtgZvSY7ObhDMG2
A2BmqcZlcmyEk/n3NfFLN6oeR7wIXIAo+f9jRR7K9DY15GnehIFKqoc+P8px1bvylFrJV8dpxbfc
ST2ElPurEdhTrsQ8hjg+5v/cB8fzcqNswsrEMLY9QNaZG3HRlHm1tCMy3a6hESkKPy4BTemx43BW
BhcR/6K7n7tLyVUUnbNzAkudLHrMXG5R1yXse6Y8RfpCBDJMxScMs0OHzGNTG1+LK+osmQAZGi7z
Wts1Pw5wgIPhIuT2+GN6uVOorS9OnZlbTzQ+Q98ZMLpAfAPauOCmayXNIalbPobizVGR0pYzVUNV
ZvmiGC+qtGVPwhrVpso2w6Xt6xeyc9UD+TtQwizvwgLbH/lLcVHFV+TR4keANBIbYxxhZYkv8QA0
hA5OV/8ohHjQ6qMcOVWax6xZJcc3lndd3U1wyEdKj3nMQkrp39663I+60NP3rXu3U5eiHF8X6ofF
5BCUUVi7+r2xa+HEStrbXBkUYx+6vVvaWPaEFWslQCsaSVn0kj/qlPDNoTmZ1G1zQPA50ubgolEu
zLM3RTfNlrzovfS0xoX5uRoiYTeXyv9LpMzlOiW3ogVPJWgaSvneZhRIqYv92PZWmpq/sABfdlgA
MFDSLU3tSAtYM4iWLFZqWt7VfCZGdWASRlHlPWA1pOYj4Ms8laStYA8SfNp0YGoWWy9pWTF3MrO4
eUYjIwWY0SVRg0BW4KNvf3kkH+fV542+jhvUbiznHBre4nqYfZOpjTkG4AOyY8UhWHr3KE2u9ypu
yCwl+wvK82kP61QdJh5swtZEhjUDNaJcc8GVhLVci22DjklI1aPMUXk1kAxuk3b8QGCr4Xv3l4Ir
RuKsJbsWlnXGJpK7oEz67kXPE/mYayO9gEqF7NMLYUOEFDQO6H+PHYdU/a/SBfNXJ1I1TDHMAa/e
HnMXIrvSpLOuT/PF6rhKqXOWyVeK6x3xGc0XcIXMkNAPgJz1jHoOhXkQxQ5XkGR2tNpuC4Vvoy6b
tiVr0kVfjP9YVkOXUVg1DKMZBXabu/9urWdhotS0PM7iZCOEMmEmZn6tAgsLbizeDAZNivZStmUQ
pFZjBQuMxj5JFzOsGU2W0muPU7cUyL0VBCC4aUomfNCQz3P3zRQunJZ/CXY2ih/DK9j/0vOeYu3i
ZN9cENtrK0xX0qm4pkRr37tsIp6+Ot592qKT1rJD8Sh+LCocPJAB8OpUy8vH73/iSmO3ZfwsLULF
jLgSQQdHDiAThJTDYywVdzqpmb/Y4DGZ2vHsrLRVyUzB+imtIQlYM8RR9b6w6niDAArUW1+jvPPb
l81uVfsc56p1Z+qemgH/pyEp5qdtgj9676vqHtehcQ64K9qmdknbROhNr/fQd1nRyxgoWMY5iL99
3r9W+vewovdlUu2t2HL2ZoH577oSZmY3MbQjn/HCd9mEv8RMb45AF6C0GIPD6dHc6gPH3y3wICie
mWooetLOwqtAFSPG45Ocu3zCJvjNZ6lp79gNXkUMfRyfD72Ssq9caCvAIV1zki2vjUL9W82Kxcay
EXRyDaFTczPoA7o9iQ+JbN6fyBrpaJIe0izReb0m1AQreJb1jWprcg9eNxfjw//3BCLaL648mDYY
bJXc1P8zlCGzzKaongEV7Z93w7E6fMLZeiUBSImFUyfNk4yNgf4YzIPFSo3SvHN2FspyGt6Sh5d1
3jLdmCkVll+wYDoydgO60U6HO5IT+9rAILmQMkJ1UYn2OW4dv5aqq9EryoPerconwG5UKepn6LQy
/9Mud1iMeRS1+v5DzyFjzPBVGPKUqiZVESYL63xVI4UC/cnApUS3ez2NLWVlpMd9zDyXMFDiwbi+
Xt7aviCvp+f6/OQiyI4NlGZOuYE3qAytpW7278uwk7ZgX3WRPpjhUEhwWs711Xl9/MuIaou6SRU2
soSIYWrKACtbNczPHIh4b+JCBiqL6OCWdK8898iVfo9ecO7o3eZA3BMrhE7BsIHMlRSLnvOp9UFK
COLUW0ZXfglg2ByEMkfdMaF9hgww8PAz7RN6TZh+znIAzk2XN66TX52NY901es5vsFSfOgupkifb
3R4laxbonMi3icWKKQmbHMEJ6IIOAG1Z+/DWaXsTZDL9uqClAaTBTSwn2/NE2vlxabaY0ybx+sSi
Hosnf36SyBn0rxCKw5KYZSzVp2yDf7HSCkbTD3oPBZABe0urh8FJNLskB3/eO5Z/OvXK9Q0C+oKM
bc+Jb41YAvQSh3Kgc8sJQctuDkE6BneZrAycKMv1nMJu0M5dUcwRlAg2mbvtYKJcKVtTvZnTDg3a
cj7kE8Yd++Fa7Rdq0LP9TJkBeVGod31YqlbCWVCD07anDGzYY8Ptqoxi7aBx+1nw/otAx9VZgelT
+W7S+tmA5+yIYHypfpE/gKndLSIC0+HnNlcjSICGoWaECfttXBlMP9NFW8z+DdpbZzxMwZhlz20V
XhiaiKjMrL5GJrc1xc8JHEHlnd+gvlYqkuazFebdo5fy3r+l0PYjh1fPo2uM+s8S0ebnbO+IGyWH
gjjFCOqKhb+ntMiVQnuf4gDU5ZYEdiP5rHbtyo0jUl0YZbEM15REi11gKHHG4JPKkTy0TXZbbPZ8
a3Nru1eH2+NWXwOJMxeGiF0G1INBQV9t3iigsOf515qOsCRE1yQIz6Mk9jbPy58IizL6sAzhsgzl
gYg32njNt4fCzj7Ot7MIHsudpUgOlkdLMVn8MZUmBaKworx96TIDCMi3EllSJdVD63UW5aB0AePL
U0jBQzgw5snnkU4i3TOv0CR/NZqkTrMtpYyRlwKgskjzituW1xqVOCJNsdwRORtTSY21zIG1xfA7
YD75nlDLx0LHqr/48xfBnR20qOLS3jIbikkVbGmxv0HKJVwAA54nCc5n1X7E3vt9+DhRfUizNv4E
FsAh+kwqeEmRLNe8PUEDtIT8jtv51f/6WWBni6lGPC7WAET39TidPZlz/gdxF4K+dJyiUN+0pivA
Jtr+iL7qeRjSM/zR9pNnVW2wQAhpguBh4qcdnDJ29rsD5u4vyjyNoKbzenxfb4+vcjXM/964xga6
KSEB/sClXuyP+65748yt1SXBqTbnHrq50r7wEKjdSpw6UAmLbiQRPpTbtjSRLgGVA56WgqLs7htT
q+7IDl7QX0/2gi5cJc9Y/fuUB+TSaaYBXybP1ptXTheWgBps/oOMFX/AiUbkO1zNh6X/vOjVJHAD
HLHRk6wV4olTSNe7ri02eZaX0kIPq6nAyV2Zsowu/MTOCNrSsRekxpLGQTP6UFyWlqK6E1BXK2Lc
aKvPFNngXT+yf6UD+JMZdu6oP/E+5PzgI4vHk2OV5ktWcVsVU1uO4yEKM2Rv5I32OGv5Jik9KbTr
LqcnMTOa45IjHeyIYF/bkrbi4tPwpf0ltssbw7Xq3xlsIghlzMKatsDZejk66Ocfmul7Kt074tYI
YxAS4fFZlpDnWb8H++1fFk5HpWLb0wS/JOy0gI0YevDYKZ6VHteRt8ckN71AJl5y/o2d2qy39j49
vLU73ms0ZCk0wIu5ehqe42biwuKWT2KDKg1VAv3Nc2u7E4+RWF/jrDzFjS5V5PSfv4uPnAvULHma
/1S+CFJQTuReTjIRjLp3+hxSSUiQKYj5LPnpn3IPa0cN3nrrpDhUvvD3v7kjKv5M/ovRbN8naeLM
Q69sr8Lczk+qxs6iAMNqzdPnaeaijCYe+cfdvukm8kgkNRIKG8q4jeBRkXvvo3HBru3eT1zROs3P
ge/nQJUwXkUfA5PkcT7cP/Dh5Z00XNBM6SucVNBCrk7w0mh1ATEZ2PX4gAsHsqhq/xh5wNCpNSs5
nC7Bv4tDE1vMG3l0/tIiIihFfB69VyktSZnUmO0985lHhWNmXMNHsfmKxiDJQSk/SeL5O0xUNY8+
YbFbLJkIWdXodoy2dVUnVE/dD4xABuss9IrkK9MW6e4/NinjJMVJqKxXw/fnn60JQglD594NHhVL
FjtR/PsG7KxSy5HUSo4r4rTp4yr/WsG4MVdZzZmStr8Y2zsebmHS076QVaDjr/pIXN6DnGB89jf8
dqDQDRgL/e/Hf5rXZKppMKoGh2vbDJLpapQnLrjYrefCzEHSaJVK3KjNciw2VXqYK6hWaugE98CK
9bxbLfLtBK8PdG+V2mY/tE16xLFBEzcdhAFjKs+8qJkqHjcRc8hlLhBMzOhxs1QZRRLcbkEvhglg
MeXgQEv0pUciEOwsiYRjoTpdiclTOvF/PWfflkiJ5rycxxaEVB1EsjEJm7eX43+/5L88cFC8udXG
i1rDE3UK1fCvL8fngOJp2nC9Hr4DXTNjWWeCKDdnad4C/iWYrWKHoK68i+l2w6+STO29ktrNXo+7
SPViZiODnrtvtN5uPcPm+r8muEjG1+OiOF/tL4k5aJNFjFf3lO+mxMQRR53hF/HfPQQPXGuB76FF
gbBqNctI6N/C4wlao8nkIvok3RSys/u8DG005V6bmLEhynNsx5raxd+t5HBAhwchfJNMw3ShHMWR
BbwI3pn3CDgQEYqXS0hBQXPuhvdsHIGtngpe1K36s6RUsstDYCBnpxXbdJNV7vyp10e7P7z6DHW+
4ymbC3KDQ9hX4/PV20NIVBId2d4Bl/o4tSNKP5AMKlrojBZpLIhu0ZnOCiomUIHJWjFaW5TPZXaW
5y3RL4UrbQLpTJx0pg0NuWrRwIZYklKVfwiKeFlRdUH2YR1nTuYr6lnMjEzdIKFn+8rMjk+A/mPh
e7LK/X1Yj3Lg2W9o12f6XTKQzGCn85wFi5FJ5l3u/XJgahdIf2F9ot7yYHT18UKecoJmUU1e8uD8
juJXneMiephFQ4YJTVh38iUG9rk7nEEp2J+VugYtpKUZhjBHmmsz6Lm74NFPaQg1lqOcJoEh0OIZ
vLSy3Qa6gwNxXmAmTyMXfqU25h+s1QIcwNWGMZFitR/uCeWPIR2ttK6TQoylZJbIrms83eLDsuBH
tKXxbUNgU2OgMFU9vhx2TM3nk4ZaNnZLKiuQq9/3LzdQH1PbcxqCtLX9p76EzxLRPWpBCJgGFrSw
NvNQl2naLBt5MG8Qn3K1keNQDrgSHdEbOWPF0OCsuIxaVxLEgHsvhlUKqkhPnuHcXW1CUQLZEFHx
vD+Qp8fQxwzMM1Nwec211QXIEDuBMOSB0Vfygzj2i+NfeFgKO1frd8e4Qse6CsWkXakQXuBwArKd
HgEYNS+EMu4wKjQ93IZrpiXyiDJZ5md6XdwLIfVHKrZX1yB9z1cJYazzNg9e3CcMKd53NX061qgf
jbDjvDLmdqsw4JCPC7yCWL10EsswbPF1vUf+oXSstNJ2jUm+bdws/8RbManC+l1sS3PrR7OGzuCo
vLLJyEH9q59yxGjjEsQ+u1FunP2QKJRmb2leBuHodw9L27A7XQ0y7Z3AGlNDRSC6qaVoC64kYVFz
PHTx+1GbxE6bGxehbrUOTck48Jxcu2zKTVoBpCDpzMeyqMusy7lSYQXf/FI6VM+l+kE7rSDM2r5O
cHr87OIGXXpK7vRqWmnatiMkOdxQCrb3BzjQkVOIlgx2oIe8hKwlXgVogVPLW/FfKgseHrmVtnkc
x514ZLU2PU+gyjMCagTovDqW7yENfcnK3Zmer6IyJ2SwPV+37dGJZQzSxC0RefHgFeuklpuOJ1Vc
ydvJvZ4NTGAMSGEvRU6eYWIwbbH+TKyPjNdlCmNFA4TolVKSXQ1djhttf0AsIObtLrKvrm5JiPW2
+VdVxL4dl1wDmz+IUThNXkGyp2RKFgaXbi487Y9p76BDJiCdOEz0h0X9ecNtPqEi14xOt6wWqusD
XneWnDkZq5tLTCKQ0Ei2XyJ2CIpifXOcHjou6Xe4Fkq2EqhAhTn/biRYoLBynlF3Ze5QY+AUa7T4
lvYCUdDXGeTP3FGOmrJw9k7vOO3Ba78DlmQeNo8oGnuQzZqrj1waBRLt1Hh0FMPUEJwF0/y04v6V
uWiaOyCcL74c3eBa4YuZ+JiWoYTP/lOQA5kEBnyE2iB4zxMkg1zHJm/qKgkzD6hnHDtSaA1aXsh7
dtHcyTNf7AoIROOGHCHoyN2dCW9t9jYcqANkcnKX+4LPavKC04usyEmoEbbhT25lLCSOrN69/C5p
29sTdnu8ysaq0p+6jVXN9RaTNkm/kooM5+Q5TOX6zRi5j3lxEDyRpXWHxk4zJc5XiLiFaT245Glo
1vMBRBaNjgULisaOOzJ+NyNgh2tfPjewuuJ0t0gPY4V4Trnb/6kVkRJQ1oY8lB1z80qLbqEJSP+7
ZLjgKoQmuK52MzlXkOY4mOzGWLYFI7ol9RTazaLtIV6C7bCJOyHnVuAcR4WW7lgK+eitEallCgN6
KT3ogWBXFu1ZOELDZmUUaXLVeq1mWkSt2V4Uh+ug/oLIsemfNNBn0PaCLUG2kqtXK0pGy6OJ491e
1vlSaFHNeZe4XDOV03AMTFQOKPlUBoqwChc05qdYS0YBDXXAG1RC0545KxGUWpaRlrNE3tGVvvly
H2Dn9d3AeJzuTFg6xpWY5HnzsvbrUNb2Y4lhb+mn7x3Wg+Z+NAh1GgtnNHjrNfl5jArb97PL7EqC
fFsPpXx8VBNRZC1qFco2QY85X7nJW/cSuMVxLNd+Htceq360VuvggzMKGf4RC59yhgFTJJIqNAfu
9hhyQK+x8R+YaIlldOY340u7liyCM2MozlEMBvMKul5MZEUJveXvU6EFKa2aa7YFfWll8t0VBidl
9czDC7RqZMakXW9EQf55lJKewBxV9VFDgsUOf9MxdG/2Cesjf3HayTJWmCEqaYL1KRLmyH3sesUm
IPpC87LHbGYzzNAAIMqBhiuRgJi+f1ZewVbgG5tAONlKL7BSlvDlreqBTk3GktpfcVfsVd0NGo0b
HcEauGSSlmV+417D3ctlvHgtJKFvX9Mw1JBKPrxowJwedWyJCDYgGA4f+KKplZuTjqws/IWg5K4A
LGHrhumYF8SihYKHqZiYGhq4G1VPBzZrM3tt5BbPa5aI6288oYZKjsLvD7V0crhktxzn95WFqF2a
n0phtU8Z5pkZhFJmwtHG4bIi0cEp5ckOxkZ2VynSnWd7YqkqIckpzkEE8NHcWFqLnoYmjEEsefiT
8DHlSCHwLwsEjdvkoLmnz+0MMKcSiLg5GoS3Xm2SnWxIUJfQZICqakyeLMTZLcr/BAlpvZZNySoA
vIJRByc2TfQDc1PmB+NCGja38/ruFr4+tL7h3FzIL+ZH8In0Rndo+XZqMoUtf8qVAnPMzqIofmOE
5VBEadohxZM+fMHUDwuDMyajSqaLMExF8Sz1vvOoT1hRKA7nMJvzigAwVEO6cunmB7xcdkAMFkVo
3zoDnv3nuw0KGaVS5EEWCyU1vWMU7L3GdqK1hfhNE6kkdQIiFTXKUUhFzoZOfyWdvh8zxzcgKHB0
Psl97asPIPfczHURrgFh2RaCP5ai96dfoD0o4saukd0+MyfTnvRFwbGIhMJAKiLyjHOy9dBf13BC
w71PaXgTZ22ugYmqWq7SajZYSno/XMDurtXJzbYSLvYSwhYG8XZXprZ+B7q0Y8rAbbckXT4HRvG9
5f9GlAgC0QaBuvImVL3Q26jRiZafYkG77eZLB55zHhUgvthDOS5DfoYco52PX2UhtW7hOz/QUqEg
8DfyC2xrry2fqhFtYOtm6pzlYiJxn53rg/Rg4SI4pRWkaMbkwVi0hKG7pIWkgmZgfAW5FPOC0nsH
GCWjrgJ4g8/pRaCkH2mHMSRK83bQblVjlE5Zpp8iI5My1/x17O7yLeWAlQJnWE+vZ0JHMeBevGFv
HR3qt8Psp55S1/XKpEV3r1H8MfPlP+khBVKsVYS2vrcGlNV3DuN5U/SXVTbuTPtbSbf5y5OAAkIb
UPeHt5btQE+E1ST899l5o/M2AdGKVDXyhriB5DKm9tybHbmDIJFPeVfcCkMSBQ88CNo15mcn+Maz
NWuQ0/vuQcdc2488G6y7hB5Ptg6GvbgS1ObGMm05WP06L7MU1FfBT1MSTLtiXhYDZZUeVSUhCJja
GVEt4OiCGpqV5ksmCCiLTRMAuIl52xF2KvbmZ9UPb+Y7OJEDFvsW9KAW5asqqhFph8weE3jtaDWZ
b6ikaNYGFNEDpB3xOBXkY6QFPB11atN3fKNjCTGJpqJrzn8Z3pTMfNEJpOdBOSIBgkWOOBtPhRlC
irpuqWbY9NxfLH/UPIkJr48vJRDvzUeFPBlBAdtrptqDrasb/ZlarVdRhWp7Qf0TCMKNyN9QnHPO
EM9xG78OfsVNFQGVLpqt041rchr6xp/PesMtAAD5JK2FsKw5v79CoSONi7rHjGbS6xbr+5MjVblb
xhUQ8BOq8J3S8MgZj+dc8Vou/3fuD7EvrCRwMLxlJKKHpy3Gz0MlAEjWwX6bc8Qtaj2BQ2WaytYb
R3vCI7OTCNrXXVLI6wkEQtNYS18sLYB2EYILakIBfgU+nDb+d57e1M2edzn2vsFbC9DS1JK+RI3g
g2JlQ0WtYRcXGeXAiX9oIegNXC2y/Ts8mYKUrFZkdJx2Zt5o5B8kDY0PbXEPyVrp8akU2+AOmZSb
8plV1z+W46hlM++l0gYucRO2gQkw8kkDFWVV1jZWXbjiA6tfPXNcm5eFKb8uNn5tAyVYPvciUeMl
oOCnL9YgqyqL1Dh5ZXuLCygWh7tRVAg744wP09n1dK6fdOgJV/WHlx7t9LwMnPZwGh42pgcPx0fV
Kh7zqJFKWIeqDbxKuQGNk2/KmLdgVyQmOuqsttxyCSISPMptxfOnrcdl0tBU9SpCte/VQABW0E/4
Az19iiBaTiugYdF74zavvzPCZh83Riszg7JekB0jDfcm/N5ryncKVKkU+0acjmx+hWNmY9zQP8z/
p9gZLQNeJdI5jfVBiZYRLiNV2FhbeOMjsUU5fOl2TUQFCjUYuAx83pa+WOQtsubWaWXQsnzHTfAk
qObW5FKEx0Fo5XJSdl0p5PT7JF1RuOHxJZGxfJ2onSUL4uZlawyCUsVqXMyMzVOoa7pifjq7uSdZ
O3G40lxYy500+aLcIs51wOgSQJqlg//EO0TS3vr366IB5RXC1jBvRI9PMjq/k6xjO1SUm3JEMzVV
c4vSydy06SeBXPg+h7gf5hIDFkQVKSRir4duNcXxUcnuaZL4qMfnJz8oEd4fDsn9DPyfIlTjGsZZ
7Y+yHDpJa3U1puDn2GfRygdL3dw0cD6EKD1SOGSYStivWJN9tUFWhRAWnO0D0x5iym8Dc2fozzTy
gFqRnOfQl23xKpKZtaB+HGrRkvMRmqaOanGE5LcysqScAf0KGyRtz4HofWoyjwkmgMJRhuytIsAW
Kl+brhI5l2b2zbvHU/QkJg/yiX3DPOBJMvQC4KDjJ1ulpPmNw1ghJ7Bry2mOWL6TVk+au99U79xa
ltuEMdjub+GqtZiQyZRq1AtOTRwfQkiDQNzqGuwQn/6XwJnGWfx1/L65+BnSKUEP85JdS73cJBBW
wm2LRuz7mVR7mWA421IFEDvth37sKcdlqUKQB9p+qQCeKyo03aqr6RrRwtMH5GVJ54RnInq0jjFP
TTqKp8vlOJAbdL0uSaaYPkydzRHNYgUcdy76WY5eapxn1mrFVHyLfC9D+BxXsugy6KFfBWTa9Jsb
LKNhNVFWDfn4sNSahhEvWIfNMR8/wi7ZXCPKdbGrvmeq0nGWoJxzcZHB4o/u2pRX3fVU5fq3fS+Q
5u09UJUJQ2TjvDkh59Meqkt8rj/Cudrd0cFOcEHuuTBmq+7epGFRA41cKhEB3/bEYhH438YpBvAk
+jc9Tw5YkJKObRS9zXLeoZpmPaplHAz6ARQ4xvybqwP3c6yJNiA2x8KQzx1gpfFTFFSCFnIN/yoU
tTnGIKAZlXVCYcDxk91l8INShFhCpsGQ+SdOmZQL6Bc8DLYAhAr+cahNytRf0RL4XaNLGPNT0v+4
HA4q9GAGXI4yh7QrvhQqORRQccM8YM7YvhWFizvkLlu+31RzUaaZTTnsgBxawdbLeujgTVbu2zsw
2PaD6QM3LMRp8I3eHM4DpqTcJgNVZI6qlS5snoewGoddUPxUrtxY2OouQatqfftj6wumeVe/MF3z
nP8FI2nGjcGCUE3VFEPmZWQ3ziQLBCRMykX58NAJvrc1D8wGDVs+QnWE82GiJVMxG96pM7vm+wF3
Lg8PKFMisAeJslhvFVjtbLzM2HClzLhnaf39BKitiGlaY802AgDkEnl7DTLZU6w7Yrfp50idljhW
+azheD9VC5eTz2Q4obW3KOkIpoE0SfRVYf5icjueVEUn44f42Y78Qt5d6lucWbRCWowNdSc2wVbC
vL84tEpYgTotDAtO9ziAnZ7b6Y2+qxH0gTM2ObHD5eCfOHVdMjE7KUYeqgVe12TxhHsgwUNA9bka
SZparMhy2Vbu2RoEczeE+OiY0VwB9zstH6BZuxtC+NPD9W9LL/Z4jv62lndRNnLIefxHwbVU8r7W
vvuHSTXWQEoxfucnoaD45tEbfUmtCt8CUw/CWhViBDegyuXg7YvU6aQlaOYig6OtakLp6t1uZ+Cd
PwK6hum/0tbNRqy6V6W9yUJqFjPfzqOKMvCjmYZwUT0f0IX+IAUqwtbFkFNORxy2qc4VKNQsTSpA
oOOQNUfMdKiwmW1QVtcqbHc4h8PciS0Jh7aRSzHBd/pEbbOW1Jn65lPxKkYfGVcnd1MpJzyapr+r
nZjTZ3AfB3Pre6bjvErHBMedr+4VBE6D1Vq3SVElp3WHd+gERDpew8q22Iaaqi+92uzYOrQp18+3
7qO/jGy3GJZwU9oTS0uwFiVv8TS6wymY/EAkAW/3mI+kp9/kGFi+CJuaBTEA1GQqsC3KkcQ25qD8
0BtV5KAKCDJhpinnqGPoFpuLmcAqPLwNZgnXfGw6UxezaOk4gBLkgbDU6LY9OU49Dlb1XxTMNn+R
4g7+UuTIdKdEaNKP2sXZ4TT8LpeRa7PrzoaMdKzkf6xG+eyOtJRFLvlp1xRndTCCmEFHg1Nc976k
eOGs03JPDtQR0ykJEOSZBjj2xfckIOBWGO7guu6ntA==
`protect end_protected
