`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
QcFiMlLsVeWOASQqcVNGvhIRoITK0S61ty/hO9Gd+oLo5iE6FCWjpC1sCOYmbWF0OI/4bWYmY8bB
OeczFZbitQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hOYkxy3vlHN154rcyqzY7SSitfoFZC0ZpAN3mHGvGxbJFVMG1OZ4ojjc/j4OxWio8oqFpsfz0pcU
J1I2T5kjIwR6vGuenYgBLQOm4e+zrJvBKHRXwB/VjEKnzNwB/rkH9n2ql7/Tc5LWJvg5qtCJMjfT
6PdW6eSNtJ9kndZ8rVs=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QHOsKXuQ+/A/odkTX6QwQcTY/UqT1x3w4GymXDd/5si2QTIvVXd4y8Psx9+yew3gUeDvFrismHG/
Ii/rHNUCZzr7cRmTS8J+O1KQD+8Y3OaDoQMEGpi/3WLYFVeRNLi3EiU9+IEU71AV9J3g9+krVFe7
DQ8Xku1TQXhEVPaHhMAoTFgHhaAenv1b5hbODVT4eGKbKNCDGw5hCAr2NojrdlHE5Hr0RK8Gd89j
Y5EHiCEpOI5hpQDN7dsMzAFzeTxlrW9p/MfPmwrCExZnnn6hwiQqOEz34MPJGvDbjmQj++AUBQ4j
1DAmY237Ha71Bm9E8wYEAeZWGT1JDkbI88T6xA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yr3XPS6SBLtiRNjZt1RYliEYeV8iMrByLbLqF+fCNTuDd2fBQqGYKPZmSJILcTeCb5Xr2hqobH2I
h5nHvymBRYsvWypR9ydObJ79EBIMxiWlzWCkYz1O72FEn2+MPVG1hnabAGwTKc+B/BdKgisWdOF5
Tv0LFOZ7766crueQHVg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pE8ebDdnE1YcVVFyDIb7mFBNhdm5Cg1ba+sHx8GQSOVq/kUXEnauBzcGSEp8LvzyPAS++Igs5G/x
4vsIuBM/etAupLg6cudrIHE5TsxUPZmD3i0MuNyZ5xViuUVfI1RL6Of+eaSyTMzRTfwMcahyWpek
/560YQCYqqxbivcMxWDsmZcSxsf+BJqx0bCjAm4L2f9yMsDImrHOuGQl2SO2aK9c6MvUyK12xRKW
INIupv+Sj509ZkXecYmb04lC3HPxS7u4KwKhVKEE2Ge+LVOxZonwTiBFwdL0dNBZNW4/uBVGPeTc
/dnZsOsh5UhFvPx4CHQCmzxBqbg2t7SMPX6WSA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9952)
`protect data_block
gpU90XKm7M0hrsMNPo1Zu33BKIqiuTUqLTkmvlsdRnteUSyCMVXoy+j4S07PYKRUHjELjy6g1JsK
DGGH9Wwul9Xps1jeIhGLlPCqsHwGo93oATT67+oO+KQoY1G8fiRbxXrNdgx/mxVUZOR9bDusXkAp
yDYUmWQ91zkgAUpZyeyhd4WkbmDAaIsgDqO5txIXd45tE/pZ9o1r7yTccEjxPHLQZAUBzbDtQDFf
PJh6uM3ZAw6jLfrow8qXWA1MV8jAmqqGWX6eyYAhgqHR185xZWnpicnz+KXpvngeAjzuPYLiCYXu
6aZ/0DNL2iQNZpF+qjpoDpJg2ndkJAcvQZ4V4BulL23nI5dI+PDK58EHItX7nlyMZenYaNXSXSX4
SqcrVQfPt64CiZn0mLyjJlwNfSsEMu2O+q9l0sFRaahtf2t/76uGn1SfkoNXlLI4gnCf9uhStnQn
YbcZE4qutZyRSEMYCXfTNcnskDIaWXCQwRRFDCnJUBRZetJvU1k1p/ojl02SId1v7G2eqxK+EgqR
JWuVvKbBSYLA6L413eUZL4NBikqfKE4VffJOYGH4kR8yZ7XdA+LLhggaBP3jAXDvK84Wx8cDvhmi
QhMFIkEweb6JFGpWlbduqhPZ/DqqCQ0xIsrsAaJSs4WQz6268+I/gwcGkJj6EYnr3a9+IXevliA8
FXLJ3dyhGymxiRWgHcJUkROHZKgj5GLTZwY5qHCo2sRSxjLi8XFQgn2PcGau5uRx8RQWAgSzp7eJ
b/I27tRzmIXySk0S3pyI+V75Muz6XZcluSFeype8sLrfCOBPruaKa7fPyk2+mRFYdnNv5nf2wJLL
J0Y46tZvt+PycC0/GToNlXMXCjGUgSUvQ2c58xSu12+aNAG9MK9lSYSzQ3LXH611/HxwUlVGt27/
vCMnpho5XSUZ7OvVbKhQFqY6yWtSOY+aRXfNzrtc0cZx2svUEfZQRHmzR9ODlo0POB8R+ECDhg57
r4So3FPwAOsIHeUya3Q14zW987qQLFR6qGsW4tesfs8kayAgSEoA6uX4EMuPHln4gHsrt5WMx4LC
fjV3YcSlDW7TzGJSAwlXwc3zBpNII2IXePEseJ6FPWG157ZrsNLoQZkCWhpd67THGsKBGIGuk1MV
KEawRTym5dZSNNZS9ApbxGQqRTpAaS0Q5ESU0hT89+oTtKFJ3EeR0MSJzBqNomaEKVKl1UMp7NkB
GCGupWtRtITohprZosGK+pOFQTfmbwETSHlq997I8ibIIb3s6LRpkCC+lqJkd4hrwieRnUXklaIu
NFrnkLF9vyfYbn88KoC3hZ//xWJZmNRnAr8ofHVDvabYscniGQj4KR9NpE2JPtD9zHTExqCM26h+
AVdsV9TecPp5Runn26D2Js62PRTclPfrZb1VK/vLrXLucQ8HGvnmkhdDFeuaIV76ouYOtTDi7k5D
sDsjkf2m7bjbc9pUsiu7gj328eVAoLPbBzoGUKM2c75+SfvsbH/Hjjd1uQtwjHjNzb5F54GJznAC
HI2pTCVJXidUEprKXTVvZiKBZQU+agtuxcKOuku+sG+29mWWCoW4zJvmvVRGDQkad7QNUADxiF3f
HUf6XSx1DiMs95GvwWBTxJUFvtp2vP7qOrMZDvXaRsX2Y7PU4RKhibqgLzgaekaoMDSSrT3kWf5c
KbugyDGvSWdEhulsCWyqzD98Evg4/tftJ42mvNPdoZrYr7nj53voHDG9zi1wTWCMkXVKTmpoNSvD
MwFQDV2Q+mQnwIMkNhl2ylI38DHd2yniztKdBFyWvIE6faPJJfsevYHIiXPrbbld4Ry2N15pS1JH
65gVXLqj7h9OGrRPouQnH6yQKmczECxKhy9ywoGfAH6Ag5rc7ktsvVIQpPI3AaXLh+Af0GmheFEB
us1d0HdoGu8BivWM/Tab6V4jt+qIGuRpi4eyzt+gfSBXqYQay6K2+ePCihQAacytDWHJvHoUETJM
VUDvehmODL3eHhe4zMqUmU/8rVpBR/njQ8/nEpn3/aRfW2032l+CwF1FcmvMD2Idw3ws+UjwrjmJ
Re4NpVYqCGZa6KAon49ZUpRmEVl9iKFIM8ISc74oFHRTzudn/bgyyES+XSPDL4a65y+L/wpeZ0uT
Uef/ioCLPNL1uGf3dBZ4HGAWpnX1uxCVQsrpvCpglb8IN9mB5rn3/7Fkgh5y9tIXZKGvJ7jMH28r
fqlU8H7pX74fyHx22j90TitFc5XVlcoSjVXsOc+qrJFr7nrY+TlB5wBfVxGPmJSfCoxZxUoai+5p
JCvN9tpey77vqjnzZ4+hYBTAgWLM+li/NgdXHKS+PnoB25SMehJjRmqipp0Z7aRtlsyDVyOkar4e
Aohfy7IPbAJPYdnlBZtMcWozawuG7SVKSE/MAXVKP9py0SBCrvQOvsnYx5RNpoA6MvLz8R3Q2PK+
4otPEZ5Dvh86JQRDPY2t2OJdT6RllHAJcGQgKJcd7vYjFJVZDuNcU17qKfTHozM4imj3mBup/Rex
MePUzA3YjZl79oP557YgcpV5kyfFwxWXo/E6oOauOYcrq0dqJrAIDcnIeQ5IKbrUOrS6MirvuZL2
qSV8ls6ssWWAnoXKTvC3HxgYfyjAveVC5R8zgvK+ei2E3poP62envHvJ8s7/s3OglFFy+O/oZAUz
Xw1cgFE8gLBvCcfFc9ABcDZCbGNd4beMoucqZsanorCwbU4VPaHmYueMHeIhWgybSwNNrcmy4qnj
1vryH1AdrKN/SV12VzEL2hoBV2x/L+5FgTYIXb5xHRtinSbnkEb/17ffX+6OIeva/zYGgo48M1lD
VAGwYJ3UBtCBMxFQcxVE+YmBJr51ycZiDrAHOJHHkJB9DnPWlER0uJe+2Hwz1RK8dCKHUC8aSE9Z
FoJRfeL7o9IkWpBFFpnLYGAg6cx1jV67APZkkoO55YeJE34QAvAekO5Jo2dHMXxcdHmgipVm8DTZ
ppH5AZrQGPaTLtyMP3Po5gRN/Ioqwz/BqTAB6r4euj+wiz51DcV2HWTYnM0w2t7k099sm/PUqFdN
5UVwXzhOQIrrfvMcb4Et7B6tYKIvr46tjHYfuALgNJi2PsILEBTU36zRbJpO6Pyi7jQePHOwybkt
+/XJ9C5Kuot26pX1xBUgMPWMSDUKezmRxv+v3eyKSkazp8/UyjoJv9ZMv7lozinzoGjUXoMLlMQ8
dG2Bo1tI5YpZ6h4ynQ4MDNBtw5/Ob5gmXKKq3ptc7lLzqsPhTBoguTDBXZZRjdjHpN4BSY4mw0W0
hATmkXBfzKwOPeA1GGzNFeHhmgoAHzW8RfuZZ5fEHI4yab/mv5I2EeUZUGgUaZCOuEQS2JiIFZKa
sV28OubgOrsGyVNJxBTVJqptzTd7lWunuUiuKbmNmXBqMqkD83VWBpBmyJqS96O2fWWzYE3vRmtH
lA/N2D0y8yB/pnAW6VysJ1c6B35S2bvGOs0QrWa09hlOaqevrntffJMBGJr68HeY301bpDATaEoX
BTNTzTnTswz6w50blUvk1hR7AyDtcliMAwW7e3EZ3tv4AyFN1PNGpjMJbZIcfRji3cktXHO6PVd1
Uz9rCgvmzDW3gXgMhJA7I0LEPmK1JBcNRDdn1ku1SfbCiI10vM+jSC3Y4PgTbDR1eULz94R0tuMl
5k65VbZ2Mreo/ogpReAsWfQ0tyYB3UUOZkPaaXSWkveV3AyoSD2WvjqF5mxyX9Rcmc/tjDFbbwcw
ww3T5mLCnMibiIQs4NMZvsCNq1PFaCjPMQUZ/HIxpkLCDbH8nhtc4uxQB4MzEwocf8lyDD5rdL9t
TwwfR7qQpKxmW7HC3quxE7Jnkv4T58ZHc4efdpSx18ndIT3jCJDIpEVEufuPVCLieODHYsAzM6TR
1sNDNVFeg018oJ7nWS2zcsdSZ90dYw3kM3PEPeubaf+ASa3tMevXwwD8AGGHyZQ410YAFbda3VhZ
wW7CScKTc2Uw7+BgJ6jjsuRtaudxqn6Ezm+QT+KeLeIy7gjjiYTfagxkFhZb8SR/wT3hTIS/m3TG
EcSiXGoKEVTuVIUvblAXtVzHN8w9JcTua0RPKfqeBshWLikEUV1UioACBy0zPaWA6x5OE2dp8Nhs
oYYugH/ZUmgJOEpTSgPZFbd0Rnrqd42ZZQNos1Ei/qUuZjEYLMKT2jSf6iZKix+rlAQ5DJBhI7Or
DeD9AswqZv4aBemoIeuH9rIj9i+F2ynarObOE56snLSUlGnNPxNnF+9jZF6L4Dmh5b5gnprY06/C
uAsrUvLTJAhujSWwZFTLUbDSr3kKq0OJSz7FM7cL398PdRo7o8sWhAngiL5QefWOrtTzX8yjfe3n
rFlkomXjCnxP3Uyt8CTOfNxzXXdc9xnUXo2+gIH2wr3Wl/vt6KLw56IHp2zWksPmtOtRzclx/efm
grdTnquy6/1VqxsyMVh+A3L3Khm/juBHzlsJ7KWsl//qgN4TGvqEAi51E7XSeq62x6FT0DcTrwZj
KvPw+0T3gUNmPaoz81mVbs9YZxuCZ+out5G/xy3lKjBMZBCCMuaiHZJlPf91xJLJI4+twrA2fuZi
ZvS7vSzcQWYuD/ATmb+I8APjMpG1YDFQSouBzmJLISuj+tNZ4uimlgXPFONXHO5bmwn6vroTFfTH
npJoKpJ6xfu4h69+aOQK1TCZPJpsCVIQe2hQQX3O46nzhxwdbUrpHJZvct9Xhcwb+kUNwIBuHg1K
ApFufkyNFONdC0aFpqKaCx7SaCkib2RiV8zzwgmNLNzsiKlvjT09XARZ6ljlZhxT7+Kv85NWhl7Z
ABoGO8XHHonNxl1s9o5UaogfbU5JtalyQ7MkBchbbwY7Gv1IlUfuFnoVBU4s/c4sZ8NB3jFx7qNE
9aDTRE1dGFQf7236hbLQkH1CrxKF7HctuZLVmwV1TFj6CZ/HJh3tqoAK7DCQjkLOi1mef+meemDt
dHcocjc8kkm0CK1A5BOgc7MEgmfUtHBLUgagpPMCODTYjz4PogI63Zx2jD+JXpGxU4hX+G3Tn0kF
MPx8KF+AVEt2Esl7p8XW4dkzYC8l+byR+K3s2ZbTuajM5aWC9G6Yz+s41dDDLRAaIf1D3NeYfjB6
z+10z6ssesF0B/OdiAZPTk2asQrai96sLXuDxquiLIJvDPpwyhfjcFvnG3R3OjL7ld7TwzL+gmzW
0as5D93Jgxj54PMpEq8OEFIZ6OPUN0wdLxpMrW4w5ADgIrxjwKEZUCvM4YPNZzL4jV2KJ7xXo6zV
SzGT35OHrAGZd8joqrEaU/U3+hRyMH5S7uvUc+FylU8Asrv3OBPCHG+MEGe5nUi7tyAUEhwJXPn8
xRX3gM5xGzlu051hpGVEDNDwmiFdK8ROQvF6j3X5lDL1WGjwvZGrkBVuFGIp6VkXBvTMy4qSFoWe
Rdf9S+HCvalwBHR3s7ctOk5lpOdpH8aJBQNlo51oUu08SfExDevR+MDwa3VPDyPqcyC3Vew0l17L
Z1URcaCO0G8oYHaSK31clLwU21spPg1Jd1DmWu/fPpeppLlGiOh8Sh8z3WsU0GLKIvwVxU55o7dX
GRhr/F1H9lhH+5hjwa0y+ZFl8CYtuHJ5pg5I9Qg14r4N/mtHA/vVXOkfDpFqtovQYQ1x9HRxdk9K
JSvNdoADfmGHaK9hIJVV7MmEUIu5c7F4dcEmgEn4rpZOknU1zZ0Ij9yIt9w0lHxQpJ6SdCYqQHuH
Ihiwx3nNmPiLCUxDOrnOIh3zqVW+IplUmy45KYb3h/2jlxLJONVn6odvQP+FHJYWGeyjGHsI94Ly
XvlqbgqdrfK4hJoiQUFqQQPaierLo+RNOvaXE8YaVIqDNuUwnhS5S/DH+GkXQm1VkCNwRlmqqHb3
itCXLYI5gryVxbLdw9d0wxl68nQkuWSStcif4ZQiCYxltnF4KAjAMycPLu6mtFYDLgqg3YyG3MAi
/K96+00Ikcy4CKJd+TOa1CfxP5tGFre2PltPngwupvlmexqGUlJJHzitjB7VrHSrW+dJiOZpJE+w
uqFOouvx/yQI8vDbiEqDExCP7qtqVs7hXTQ8ReDAHG4EAipAaLafrT11QiNq+Fe53nUgIYwpk7Yy
zlXxNa2VSp0uSJAzwzpGlXbkYSkV70zup3WKgeDy2NS8vj8wQxmbgaMa++pSIfD41BjyR2QmKNRO
b7Zliurci6ZPjo8xznAxGWJkDU3yJfhPJFy4na/OX8pRN2y93BQNjpGHWTgXkogBJe48/LZXcUVW
CTzsSyEmQt51FYxYeE6geJd7uJfqVZDB3GbE3qIIaTN2OSuDt8ccXecthtiyHa4TTqDgkhLDFFA8
RyTgqmShkJjFy4tJ7PO6Cy0ZawsLKTvCQqtJp8lnxWsJ+wSL8EVzGxqdIcsgMUEr7lnlqL4Gc/0w
qLzuAswa2yO+Y4+sntI7qweb1YsVf0yYXGamHvFA0rojjJSMjK2Gm9p6dyiUqCZpVppJOTUAaJGO
BL1sjASUru8GCgRGWLEyK/ztq4XJN+qVeGCqMWyJyaY2y8e5M0xeYbcjDYeDQRBt3Tz5NCYSJ2k7
WBXeEGBM67JLpQiPvbtVQSErsO5Y/GEAk1wuP8753D1jja5lE5gRAYlkPhf7N8XgFY5953asAocp
gzAu0tYfUN8QzJyVaOERnBjPC/NM5Gj9GTacizu3h5knNVwsl/crDghD7XpLdAUN7PB1H+vq+3mX
Df/ruIZFz42MV75tWVL7/HFK20OtUsTMRW4tXLcf0hiqMI5yZPR588sjK9V6rNOPuy7M4xgNU/Tr
iTVkTKKMRyesE74FC2rj9nHrLqu8j4JDsUrcvNHXH/Am/ptJaOk4VePMPE6GPUSkzfPezejBwr+k
CgzoOVLT+lB0sBrGnwdqcaapxOcYn+jHb5/McmWyITDhgTM6zEskiyr+EcJRxFFr3pvDFYEi+Joy
PPsIwZqWSa8P8PpwTNFaw76ajqCeYNEDxcoyJJ1Wk/Wdz0I9bsVGpB/V8N1Jz6j0zIDwrAjdEsis
frk91sPHfVHe8yhTuobtkpxBp7g89EKCVSBGfhCEIyTkELO78RIVfCYw8xcIigbAp8vdWF8YaP7x
lUi8L0GaVyBbFZgi+CLQrfjQHx3bQxsC6DtOYCaYXvL0JIjbT9gHjQ6t5iEW3oMhAk+OCZg4+X+L
rJkh8R1uLA8B1A5TZ7uaFZlB8RxmBJd0DbLlMa6c4Ncj8pe0VmmPE3w1gc88PLPl7XdfhhS7ANN+
GVtPXhBty1x7btyQoo62FMqJN/j9ZpUIQqWI/HalDdHMYCX91CNBRsTOS8lIhvHJcIppEkqjKW1t
LFphxlMCVawZMGuPjH2WGu8sy3xvsBaUpsIfXzeER/BbcjxAGHMovBBi2bVAQ7xJRJVw1i+LKq+L
T8A/HDuQdnKDaZFvZ/HzyTJka4x3PSdPSIkPuFEmQqhxaEvDzs1NEFVv9BS23B+JRSoXOeGmX0Vt
5kZfyDHmeN5chuB8G67bn4rfzJxLbILgaUTc1PJYnyFZVWCEfiwgJpY+gqYqfCopa1YNUgfra5iw
VfzP/WBet3GBSfWRjsHKtw5p7b/Ibmo7H1AQ6q1LVu2I8xbeh4vQV/I52ByOKkHJA97nm4o+P/Fe
/GiIWqfUtpc0O4i6zJLl2UVAYdt5zp2dQqZy0sk+PyUmg9fZULa1lF/2mp5Xjfzhliw+5RQs/Lh1
YqPQ5xb7e4+OT+q7SW0BNy+9ox5ZYziFHJpFN3of1cPKk1nwhDt2KF25AHJdyaiTQDX4VCu14EUM
FMUsnMD8kWnx2gES5Og2D1JJfjAAEFF5BNxmhJu04b/C94j1UR8cVLweXehffKmCvehbmmRtp5/f
Bq51xWW9XB3iqA5vIJZ/oZd3q7HBVpBSHeyhgFmQq9qd5+GPqEbvaM5gEMPceu8DHx4uDmsOWjUu
MJY7zmTfpS7XMiVc7l8ezKFdIPH9RLpEnOBOQrJh3JuX7PwbkNfRIlQEjIjwueCjQL85WRpsEz0t
Vqe1jBw1kWiwUuAYa7o0KhCvscq7VedAtuU5A90CSThbDIeO7lZf1zABqzR4F5cgrvPIYp0nrdrd
E/ZQhlyMKRwZWEM6yEqRdcFbg07kj1Rf7NtMKJyeu7I4fqK7ccYMNQxqKodIKi2hZAFzmXRJOfky
x0b7NUTC71mm1O2/MG0jmThSWoMQPWS9gGU54XvBnyWQa9gYDRNrXd1M+oNGFR/QhPscIPhsPwze
uCXTaMRTar16Fv03H9ZJpU+Stes/6Clu87kSuboYOEY3D7fca5vl76TuOZV7/SHwBpRsyXL5bfkq
gQvYkFgGuFoxGZKSEdG+uuTHZ9lJLkimicNXo0Tqhipe1imEe4McPvf9NymVHSksCD1YhlNfh5D8
fgUriL6Wy5ECSnqNs3XDsvDuDiciUFYq94oLmDtzrkgJcfwS6VC8/3e9y+/sotOCZJnryUOaJ1R0
Otvmp6N/765mNATRCxuQk9KOr5J3fCeNXlqf536yYVmi6k+S4MihkBPoe/m7TWTiYvcKbEmIHTt9
thES/e1WpWtnRIUZS6j6+yhWiNvcfkjhKyO9aZTP+43oDN15K046y0mGRJoBdIiTKgWeVolTd0GD
eawcSgF9/aXYoAHBDRBLcqNihqjXZ3tZ920oCYKKno/hhVdKyT+Hj0fs+MqCvEDlSqhkGQjO6mr8
kEKCBk/79bObhfz/2A0yvuOYFDzv9aPmvpJtISXcFPStsJFQ4zQ/H+9HKIhFmiHuIOVCYfo67Z9J
/TE94f2D4JtkQTnc+5Xk5S8E/EU7uaw1H+ovmiXiXspKVqH+qYXuwiVH/tqGCa+H62FKYIXXmzbq
7+KXGU5jg1K9AWeq3uc9mvn45dL0DzMN/ISGVD4KREzvWcmqBnsEmZCWT5B6Qc+VP6ANQqrRYHGR
ujZ7pYWi1CmZWAi7gavPT7MHV02BcWyZ8id05UZyDmInIyP5LbonYWGK4HS9S2dNjqTnQFcbIt/q
8Ib/NFgKwbU9bg7JZjMxnUbINKLJgnWyWD1Fq0xqscje2PpWn9QQQS7H1PRsoLr79lB0Rx10/8g5
wc60Ko2p+tfAq9mS+DURv6MlYElKVIkFJBKVi9zqrGJQmWiVAhZz44hkuEk6WHfWfgHjdJmcRO2O
L41NaS1cg6kI88fjU/pTVbPIcCg5sYsYHbjPhroxhKkCTWRqjiukfqwQza5Fl/tn9XQwi23mPk7v
iXP1232xM/5vAhHampCf3bmxUQ0tYe6YjSYCaTBxQMCCUT0NbYjtXIkuPZMBJYWqQYPmAxnVYlpw
kqehtLcXb40u86QVqr3MvqHrsFNFmioE/AzYo62mPGebL5qwhqgtGgrAidZtUtoe9uXFrtR4AY6q
IKIlJ7Kv87OfQC9YTB13VS8FJyGdpaOWKTIisgaeABaeWrpjU0GK5/Nu5oWpM7VMbAC+iGe3ALU6
gE+jxhM6frbZaqEJ1XLrQIARxjq01kihbTTJ9TzpMDUYvcmpxNbZV/xVVMYErsACvnfoa/UXzTnK
pTae3XpHMP48krynxJmeCU7uSnxOt1a0VTvQRapOoa26ajwY4mWNFzxy6y0isA1Soi8ySDpH45aA
Aln2Qemn0Xb4mmZIehnH8pAKh3b/GVQKD0AX7j3tOm6xTc7ET6XFZmhmZ1KWJarlisseiEZQHmPl
BD/eZXxEzptkckjphNOQygJEYOQ2sJRYGTeWDIET94kIRvq+05OR6WfWLxuRvjnUsRniBLD1gwuf
m3bYdlSrdGdBe4Co54H4IDOmJ3cMobxYa/SsKCWr6SkZLlVwZ+Ug3Bfb0hjd7T+Ry+sZRy0JNwWc
faiXLeg29OXLmAgUV3Z+qxJ3TUcPplZDMy5vX7npKnxZTSLh/3mHVgOpEKvpEymU6lubuOtN6M/W
RO3crMTJzdQtHRl/wxuXQC5toxdv/i0GfAPYBQD/vv22TRf94/x85b5Xu2PpHXoeoAP2JDZLFi7K
VA8/jrCD1/EpfnhE4oMoVLds1a2bgEO2s6bumIgfvAxzlfJOZph4eLZTNbB85zP/31mHlcR8eUiU
5yqSeikdcBZ/QUql3+ebqrLhsIBpJgpONMMKwF2kPpVbPnuNzQetvXs87WpqpW2Z0fFfc11IgPBS
iI9c1ORkXau7/kBkpOFX1GtFzaMPAyjo10uoyQyfhH9euirtb5lDIA+3R62kBfhQuX/XvHkz0wEo
F4tFVUvtqQTd/z2ni0RG1bsvvaf9YJuULup0Vws9ctNG9yBdHjMn6bICHc1LbssCcbS9T8lLRZ6X
5pSmUXhHqA6JtBiwoqjkeB05kc9cwKSTbLaBO8n7bv2HTjOgQ1//jpzHMjngrH/VFC/AOSzu0vIz
xo6CzG8IZkNRLihGk/XzXEyBwVT7Zlk9K/A9cehHegBcgLxpgiPxdVC4QBTHQs8Jtc+dznrRdG75
V7dJuDhFscOVz+zzBo7o0JQKDbjx0ZXWh83xwF+rLKnttfoJa2Xy2a8uCuJLtP90jhjvsi83qRjC
sm4JIE8I3w0AIJVcXBre8eXAHbbkEVG79QD/LK50SlJsOFPFmQMepWfytodp+grzVhaneQMqbhxL
qWXjsqHU9RJOzyiWyf+6rdAXPpAignCLY0qGLbhDib9LvYhEGt+qPBJ8W7O1tX2yZWQO778On4Sx
3EUW+t/pNeXCnPeMy6dHRmJ6UyIZeJ61DcOMiXEl7LPrK8/bCA4eWvWJcJe1spQuM2MNNKnu1TY5
BHsJtyzpBRnsAemjbi3miczVRuObTYOtevg9mKtA6dT690hJN7ex6QpK0kTjDt6KSUHBmFvCMvaG
pX5qOBmP1qyrABZ1DyQL1BHa/eq+0jhCAw9YP7mvBCTqXWaiByy+gbFCpusTnWupbeDNpFbKrVU1
LfHSt8nzGzND0FPKTCLp/NuIELvLo2WBiQwhYuMdKSjbosggaXU7IW3wh6NTxZrpX2jjOBTkc1Rz
IPYP8Gk03YJ7zAUbtCDJLEsLq7w9IlKKhwNVP5me3XQ0JzlGQZkZo7LWYGBMrHewjhp83hbE1n+f
W2MAB+Vp7JJ4DoorjfJQE4I3EPJlwico0+tORDiOLXwtI2yA1qrRECBQywIjI21qyP65qHpyPm9c
lvaaMfEtRDsErD3C/rkOMUbbraJZnzwQFQNKS2wZXdi+vRp5zOsREN9oVX7JdRo7gm3uMmk9b1nn
FkdlV+IwkIBSC3h1rvj9A2MG3tHz5ebKRrLAEO8BtNMZOY74Mrrs/OeXHUl9ACSZe9ibdmP45NMq
oiofGfyZE6cBvp4ZgDY9d5Pf4iKWbBqkuB5WE+wrie50Z86Pl8kz0ybcEEkg4S3sAaJvrBp1H+21
vN9kMdRys5Y6BQV0Gw80DiGiQD9gLQ/3bUjbmyDttBUpOF0Lhe4nu/x2HrBPejxvRUQA5L2pHRjf
8wRd+T/hpzxG8i8XQjQLqdGz3kvSZlKi96+Zm2R1u0wSC+BnbPEcE3gpghhLs1g1Xjy9PhfqoSoW
+GJhRAlHEG9zz1qlNTRkGBq2ku+psNIXyK2+B8xkiVLy4DxOB3sUMV/tKB7ZSMwA/4TENc42tBWW
MJjif4/MnUztsBBilQWhWMJcOdF+EQGUr8CfuneObzHDzoRHToq2FXFe/yDu1xvFKFshhc7xc4Hz
hzAjz5O9ZxMkqkbgUmcDSw38vWa+79WPvm3OGbHGq0QMxd+CeIqg/XYvaM4MhXHRgDkR0ZrmFsVV
qh4RMlsAuoP0xI1o7R2VjkSVQZWn6/62Hw9PhztR2HBO+ZyuQfgI2e5Pf+3OiOnA953kOYVdDgvB
yaHArcP9zYZOnFkaRoocMwkRXofTS7hcxcDmZTaPE2fcluVBjiTiKHkgw7IDmdrnHFYoOU9/7y6V
HFIOeNE9M/Kr7MB7al0qgAcumQRYbWS7TkFp2WL6qSLPHulTgI0l+Dt3C8GfSM2eT18CfpgkNxcW
3MUUZkEgEBwqn4J9uv1cWNdegHhRPbHvoxJf36L5PK4iy4BHOQ986D9sxs8/KE+Gxte+pKpJXJR1
w3MIfbTkGEvXsiM6YyOdYtFttMC52itzz5qo2E+Jp6BsfwqsBC/gQ1jdXBl1u1t6xK0OZLHM5PCR
0tt0LRrJRm/ESUL4xs85lK3fzy1EivR5qveF1ypUNseMiTJRnE3P/8vDE2ebq7aahmGwg9lOJLV0
NAB61tq03I2VuF1RadGyNFSRf2/o4OiHh1SRVMf7fUE6groFH3LvxhXe725rmcYNcG8nS3I/Fiiy
RuuTCrX+Y/kIXmXUKYQ73z5IL4x/5+3pAYMJfPzU3+kEyfjPNxamWxdu6oOm3fSxH7MTIlz2NTd4
CHPNj08xaStmC1J4tcPL6otRZCYBsIEWU8X1wAtE4agHtM8T+gYVn8qzJtxXHxWnGOPZhkV0dF61
03tOyyJzik+WW+qlCaUi+WL4ONxSBCUJa4iwWUW7VgYTSTvUkLAjdjvQ726M945JjhXuR2aJQLwy
yC2Y3Yb4lrPJ0bLOxXlUn0obDhUcj8R63IcKlq2l3OJ4V9umR1gO7vR8jCtvvSVddCQBo3Foiz9p
CVAX7u0P7Yeccx0iBOxKRiG20YwouoqSTld52TtgIywkzCJeMhsRdUSumRRV/beDIp/vTmigzH6y
AvFJH8U190DYvUNLZH8LEgDL+XFQvaXZhsETZZOg6cHL/w+K9UN7fI6aq5YgfFk44cvSKs0CxzvM
1T5uUCpkKevfcJlMsqSnZVt9KxCwDYgxt8Um3zWdxJrmGGrbCnzYKylB8IasfWekcsA+YT5A4Bz/
1xN8QkwI0zzeO+X3Udm2UYes0smy2jLqc4Ij0zlPo+mb1hfC3WRN/gfdNS9S4dsN2Rr1YGBmcZJy
EvYnbXDRzMqRkWAAfd2Y+sT+lYw0w6Pb03jD22ij4Nn8BnHxm3XPfy0Q/g+Zi71ubLeRBZ+TLt2W
I7jGEB3tkriyrA6LBvLCy+oWnL2k9YSNn3Jysw0pf9KEhYEbswl4CgrFd8GX2PQd9va3gHmmEnv2
pegLwl5rzBJOLVGcUU0+KgDGxi8iXOxcIC2txM0iOo7m+dsSnMFj8YOMvh82P/UQ940xQv+orIKq
K0661sBK5inXvDsXyv50+F0cumpnht8cc/2mjqZblRaayGY85s8VBXW0nk356qDuEowy6vuIDLKw
9RY4N+B/bWqY1nFCH54IZm/4fxPbFBm85IyaR5FlldoRBfEesD1w0FlrixAcmnkuD/RYPobVZx+1
94mhXh+LlKA8v8+JAfNltDdYH08qWrmqbMYwTwcczguZvg==
`protect end_protected
