`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MWbeGS5GHztkzJH8Bj6JDnj4HZJjf4+Nzir1V/R+uj14MoycfzzuWOJUKwWvqaHc9n24ZbKzjSl0
GpQ6OEOz4g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KRqkUxz5VKfYBpP8PAruePs/r2d+U+52d0/GbcvW7eqweca3eo5YZeAQn3Fvb9cqkYtjaVQr9XTj
4nXCD3i2TOtqlOheTpliFhg29UXpdk0N1OAaBYwZgfXRXOV+QgMJ7BTqr2Z+XqC4mJMEpAdv/NR6
xn3Oimtm4QIzCWsTh3g=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
n24gyLxDzNhH08HAS2S35alqrhj9OK5eSVtHgB8riM7xW34gYJOQsi/IHUn2K+tU/XaUZG5d7DrR
hsZt0xuORZnw3zCwebGbQ8Zbjx1F1rARutk26AqatWXzNErWrfFCY1rTsw65YutWKPiiNYcj2E16
iGukX5oNAGVT56IcqgEomXckOPChlxhfVWxSSNG0qLVlAgiMxPL0qIqICbObaBAc46ViTq77+TyM
2euSWtPnGGzNnOAEcaOOIqZqgYcE7P+yySENcUJqcVsmJigkO2yqOLEaEeISDQlIjUjjQ5waJSTo
XaxMpDHOHpIh8uTk78t1gBcra2hTUrV8G0nc7w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YA1jSNB4LThkIcXsqhmt2InUL/Y6tFhXnUyZOpdTwYe5/Z0o0FpjiiHvn6h0IrfTMO35lvXdSn/g
zBGdmxb3c+lEsd+Z28+8eF+jpPb/LKZwrG9wYQqfJEQdM7mTCWm8O/iwdUWotCXuceWEfsIqdUqy
V6Bd7xfkXV8NOvyWXgQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jPyYrXjJ1/WswCy2abk7qjkLc7kyaRAZFUZW1yyOiSnyhXzwThBhyZCYtTPaLEdWBrGYQBdD1SX3
ZKJbbSbeBvEeL339fLroFUVwWytX5M1hz0pxa3ErdKUjI3L7wuR7RPEhBp0QylraTFeapMuT+b9i
o2cI3By+LO8RBpjdwoiM1seEYozTBctZMzVaBOxJ5ne5cRuo9FgbfUi0kLusW9io0AM0uP30Ktnd
t5axgJ3dclQXtLWE33I8wR89FbTLvw3XvFBiklUtxHHbChDZP/SPkFXT7RW8wp5WoMz3tfzlZVk4
0tw74CiM0uNRlbYA9Gaw5ay/xC9FIlgHqLvcJA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5472)
`protect data_block
qYlXyFIMoqOcdxrvFhlMYgWqUrS30hdrp/aPpkstBRM9S2eBsT3tciEVB64b5Qg3bIH/+/pW79xn
JVTFbDvOuLGu72GhYKNWE6S3YA/y6Vo87GJLO5nzzSW1Lm57lxKDgDt+h9a0ZYvNvBsFni9ClZYv
+dhYlWOsHCVu6G1VOnogyHWHBpFgqdbKmpX+yPT1PcbboAHfBkl8R41k3nkAgs7MSUc/nR1y8APO
wOIXSMZz2by/Q68YfogcY8lhb+AkymntgXz+AKlR95sY0zXr8GqUDS20hzDYWlG4Hkeh4N4xNt1b
CiS8Cv8g5i8NsGU4zekHeIKUDXGflFoP0PkTD11ySwXE4e4ViO2dRDFIHiASaBTPEL3xorzlN3yV
n9NRpHfZ9Y7qDBmVnbSRiHIukG9uC1ctBrmCgtA1GpB6Y/hHLnjZfUmshUBveIvbYaruP8+1KUKg
Gii1RGtViy9loU8omletJjmBnIxxYkNgCMsXB2TJXNjau5581ECo8ls13OmvmTGFICgxNrPyCuAu
I8IKRfKSG/1eEHyDWvIwCT1z0rICPQZV29rqW0JJBPL+NXb3PrHc6hKI9wwJvJPPrIOeen1h3RFl
kIj/WF5/8sseMGQIfInpoq04oNIxehBHB8cPVfgI4koB4gF53NKBXD2V03IzG6ZohQBl4r2xI8FK
ps0T8cVVd0cvPabgajLd3OZm1SnN6YRuLgCpfgB5RSlGg4sMC1hQlzNAqLDX+Z9pSzuGWtiKP2oa
jHgdVuhryQ3joHRk1d/mMa0uaDg5vSRtTJjZKTfAgVfF2cWHnrGMgWrzBgHPx3vid+utwYlsvT+g
kHv7I/DPcnBtmXfeb6mtfiipaFw+zs7eO0NrUsN3joURowB2hlq+NuA83373eNd8IWWo++ewgMrR
B4hNT2YUj3MS6xT7ARhqAK4Iflmd9OVKWmkuflk4/efJvKRUGPrGp2Je8BQQ2oLUJFbUevCdNBf/
vC/5eWg13l/zfCahleM7qCGHpWWhgvOVWLzRNTaKMRw47MgJqp5EZLAVRPvo85NV3DPEOkVBaKd4
uCa6ndr8KQn42yDL5H3HGU2xV7LSHW6u6+iNZKTv/Bm0sg+yS90gtl4Y5gkXZhVcylpQqAqmSF1l
5U3y4dbbJeuhBRVIn+mYVduX1L1RRESu/JKyNDUDojmbe2hiQDXeC7ZA4axA0VNBNG1fFRgxe4Xh
lbWrHSg9F+WEWOpvDrCqlsjd289F1/yX6zwxldxjRifJyb00xI+aFOSos8hq5hIVROT4p/vYMC2X
9PgPNsqCuj6VhYjgWQp0rInsUtODWiS2bemPgdZkOr+oZPBJcNhtRX9DGxUZvfarVNEDftNj4OM7
x1dEjYSnI6/O65OL/rjUXiIk2T4OFP68DQ3+FT1zaOMQ4qxjqmYDf04Qh+78En7DN4nz5xBJmf0X
W3wwbDfF2tqXueh4Xh535a7r/Xupk11X+JL/9Mpi6WwEgtAqbIuLNqJTQygbd3JB18tLfDahcmfI
yG0i43oq6SYIdnKxsqktv6dcgaWZFC3Cm7Hor9Tpaaj8D/h916ehncWIp5tSnD42qUb00FV+D6n5
i9VC9oGca2Hx3svfpoV5ZtuW/0KgPBQ+oY0zoTvFdbsxeA8muaqBPGCP25lUPBeOWQP2Rsduzjxy
R1gcS2oLzLHuck3F2MXlIXC4Q+AqAWB7VnWk/PK+h+Z2MMwr9B1SFKMZQqIuunEDlg46+zMC2hf7
d1ZWtF3n4JXyZ+b0K9K+syYvFQpZOO/6rfDuLZdmyBdD02+IkH7yF1vS+/p9QsCXNJ4mcPi40ClC
1/FYOgd75fgNIpfSu/Kv4EF3EyUYQD/p7lMa5hEv3qc75g04jN4jyVhtOQuLqJ6S7fo8L9bLQvlz
tbHQPlg4TF4akxposxVMqjdi8xoseUJivDN1P2FE+BhyCgKWHww3KIwZzoTxRvROhL3xX4mxToyq
tNmoTd8OkUj2RRwQYgp39mrlnjQorN+Fju3qaZP/ybNL+qNYv6gV7DXz488xPQ+WD+bbsTsAGP3M
bz+MEwn+jAw+DcSpE7D6NkpwLMhwHFO5cKGprhTdbH/INARjJHlTE5ZWaTfhE16pilZrpV02owER
UgPwvN6WyujjuAnshmd5wQV+BFSMHhOETKUrB+BrQ/d4yK+UNEcoKRnYfM09v1G4fXtzqJGHpRWR
TCGAPupcHdl1MjAZhdqiCoPovJxYWQthU53Yq/qCSLxVqcy3EvNqT8urDp/HG2kssiRennENdmsR
BPc3bgR00zmajKbEhSDf9JIuvrV9w5FpOl/JxKCN/wZ6OKUW2FvMz2sKJjAcEf2e7uuxKB6ICdX0
n8LxOZaCvcMVxquTxHF6EXSOagdIOBR4MOTeXtRhYsjwCQ8XRbSZIS+6ziJbz3s/AV/UaAO0MBnc
tfwjcDPKXQhKMY7FtdWNkQUwGEKv5DIfPrvYc9tfrEjEoXWKw9yd2VHjUHpR4hxG5N1swuQfUAQD
cQAArlJcoC+FdsEfjTFLp2NIrP7wluSw9zicEHvi2Cmq53JjQf2QtgQfuv1UKZvKF/3VqW5pQCAg
yd/h6bdTLo3a/iSV5OtSLZbApoqM8Exg1caPhUgmqMyFG6/PknK0HE3a3WWaIy8WXUiP/ODLXkwl
ojHTuQPCLL7uMnCu7bJUK7yUdmF0FEtuxPVvj1JHYHsJbsYzpFC6WDGn5AerDeons42jXRTlCRZX
uCr5OjCKdcptMcvPFo6BnwqIpecdsQZhSutJIQQEmTik2jJBlslXHlOnVyEPx5ELePyQxXkC+FOy
DBlMpa7DIKkXlyGl8FObwyOPT0uMtsDY6zNBDgloa6zmj/grwhMGsic9feFg1nYH2Tbj8cdWL4cA
UOgi67KnUW1Kcidy+PMQ2cNTd9klIqo/K5rahAdUobwVqu9RoZTIc1bpgPHivXqpBMOCMDtIX+En
4vKWxsbWVAc31SQeCft+sVehHAsC8cKZQlAc5dJJHT5/ypbGUT4Ys9c9vKxi1wnmd/BIxm+DPgO7
y3W87u8kkKq5MyPr3H5KW3+ePfZpdSAiQRU8pfd6cLPXng5QYbF1Uw3fb6MemJtPm27NMeaAzjCH
tD5ez5kCxRsibHN7q1Tc6sb02i83oZSAogYz8t1P4hOBEsS2dkLmiuuijJ+0sO40GhRUQCcOkfKP
8s14LglMjSr1mVtzueaOy03qj2QITXZJ5QfLriCUn3r/zV34ifwpGnZxYtSESMxRNmKpZqxfkR3h
U7WepaKicqr7AIC8CU4n8XYlY6tVbr8LBPITetTc0Yu4bkXFsI/BB47hW0Wi0WbyuRmlMnnYT55T
bDHyXk1WMu9mA2EdWVAnxTX0ypoV8BBHgi527MUQJEyDIIconAUUYojZGOVQQthSFWWxHFB4PenW
gX2ZDsGSirJaQU1Nn+YcepM800AQ6pV2HzlpVXqhwDT+gAPahqTexTN4T/Rog6dGNr9LIyIBoepl
7VcxqZ+gOb/FfwcRJrxgtdGCKL4+FKzdRp+L/8dWw9JjsOlIhuakzlQC0CcNXTmtBJeA4eDqnALn
3yvO860H6oiNsppymZirVsM/cquamTbke9FyDHft3IsNYfvFRkjuHk2d8J4yx3t0pbZGDoL5z/+Y
XLYJS/zAvkVlZvZz0hY0hJbGyXa4VX8Dork7JAAOg+pomMyR5Ws784ggzDxnL36cH27bFll2sTCO
8klNQlDr2WhAtmiJcg0LAESnmDUtKqWnN6L5cr46T6pgBiJ5VNJeWMY2Lw3dBiTxDNlX6reIzeSK
/OnqhMXktO7IYaL6UEKYGqkqHN8/sigbvEkXMDFwu1EsYNNqikv2qUjoGy3rQzOG1xDrVUqo0eYH
avvMAzqL0yYuWGOi1yxrY3YYu+ohYGfUKA9ZZ+ew1PEIm+WMG8osJ2TPKY87rZunFiGY3slNVSvk
9dqre5pXBbXsjUmo+IF3Y4SK2n0S1a8HfbH4QCmVTguVPYNIMCnqbIrzHroWT5gc2L4MkaxUtpB1
QEeJa7IvRV9FqtsQtaAzkzkVEzfyKm/Ckhq23wI3c4UN/mppQcZfbpcoayl4mloHMsUc5fGAxdYb
7wQR1FBXqFoHT70aOdl42As+LX3mYaGg8JOUD7WivzEtbHq59FeyEqYrWuOBhnlfxzPywaI8mrzr
3ZqxZE8VpWET7N4pLa7+fwOF5PgD7bijQ9lBwwnKsTdReRJEjOk6QgZwYyYpju68Lja8RoXP+Xjb
cBzwl1Zq2V2GYV+OnDR39HP4RrRI1YGVZidmdSPAmSLpBL7ucfo/nHLnoKrgrqBqD82ekDv9/V7+
VGkjhYSW5yuwxL2/DQ/ZIvWVGqIPUogSGmGFZh7eSI1wxSkz0SOAyC8skWxNduTEaux7NbhDyGSX
d5ObhwmduR2yM4pXUTci1l/lrU6ah4DuqWOCXc+WDrD/3l3Ka0ZgIUeHBIqhKXlStqQJMsFkdeY/
osknxx9clWfN2UIyaF2zkKDcILDwcBc8ym/o5GeuOh6Y+/lNx20f4dnGo3xwQOYBNTTonxQNH+TY
a3itngw2/DDAX/bQAVmZvwBkoLBiHxxy83zJG5UGYoF7znabyrKigYz97l0zjtngDY0UierT2pUV
Ced3RuosPg5RPYhgzx/6nC8otb5qP623gaiLA87E7nMcevT7p2PT9WLww2s/JVxEogofhwuJdLMQ
QQT/OpXoJD7tPfY26fN/Fu/d+p+nK+zPqPG4W116J44ufgSanDdkbwu4SH54JLakT1g0q6OsqQqy
3+VZTEUj0rhaHorFKhwrMTtARi6fYUUa3wc0s1GgLdLw1NruKkJBC80xQN71/HaadkUMF0CYfM73
HjeQyzAxPAeWPs6Dpnlq5slG/QSMjKtkmlv/uXEbbGMOUaatcOSzdikI+eXdx0M7ApV58n+9YKtw
Ws8fMXoQd38iwym/fQaZpljb6OgB1+YL5KueNMNVZjogpDo4sBRKutMv9StYTVJgd6L7h8ntXuib
VY3aJ5tt7GWfcOgG/8MBe0W9M5k++hQ7XZDtEUvYHixCA0TWAL96ziqr5EckPevy+OeGYxbDCEQG
zjbA746dN1OLiPEaG6lBh/gMZQnO3Yub/pIOkfEafuPdgqqwWQxARU9Fk6PtoGJoK5Fj51+5uBOV
H/ZiEXzN7zQs4jQuGZgYNyHGECtoL2lgqqjkYr9jrd6Kij1kBEmo1MYkVeug6OXl3bjo6ffOLjA6
SXlzO/6ZjKkCAVEdSCUzIVwGWFuyqGFxNms8giMf0YdkGwuec9dbJe9ms6d89LCdiXIk+Tr3BQAD
ytQDm2+1iey4OlOIqcdURYoDtTlTU9e5GGWqJzwhfXY2apel5t9BvvISnY06gcDLIqfDj2BhT6+M
UQFJY/g/i+hNCv99CN9DNIkuJ2zK/6Me9i3p4b8OwrdncS2JtEX4qoBAvqrAXGuLETTlEJPOEkak
mPIGdv2Y46ebXfyEhuE72t8KMASP54ZvkS3p5T/RI8D8pfyEBtZVKsov2gfGoLzklTEK8Hf81t5s
Dti0OwEh7HGT42KJCvZ0/eXyn9c0B9pW84ArYAbxmS/vluiB7tv7OVK8q0b0C0v/R3TNVvUR9bzt
g95hp180u213owaDLr2Yp/43zE+UHBv3WTuK9uPsUjH2/2t3p3BZ1/4QmrxpSwq5FxPYB1aHDTmp
jEnMzE0vp3bKlULWfz3ymQ/eHDUVkyW7yGQ+UXHZs75YONpR0geAnDRwZAgw0gCLQ2KaWEHYis+t
dMJGQXuE+s7JqAY7cZJq3JlqkRjTQFztSSxWbv5Y0q7/UdQ8TqpJ1lQ1oom4eVWwkI1ZPGtolb5g
ld7K2kDsIXg4I/QZkejumn/ZrQVgkKqcbsSCHzWn4ExH9Gl3DUopA2+1jpEfrfJxZUUxUCdrg4/m
jT7BIYwgysJtEeYTe1AMsBSiRTUmsS5r/IuMAE/LlkLjiqHMXY/+69lKf42hdVSuqoKW/sxfm1Gb
x3we/26zN1SX/HRgk7DRH8I8qJQw4IQOBrH24HdaeiNx0bTUBcbAson7ndvUitl/IEbB7AT3CjXh
isZWvhs2OkGPHRJBdLUvctKMHnb+gP3mbuFJnKZHOk3FMYg4GkSpnufKsv+UivgPvYIBtGyP3+F8
jnXOO69wbvFnfBeQ4AMHKIZD/ZBuNCT7gDeFZKZig3KlGg3rXXrmYmvPKb1qkXU64QZPNkD0uqxj
jOOWLL9Sdxv+hOuF65fWSnWbtFdHF8aOjFyuWU9slyJm6MdXWK2cVxiXM/OgzmC+zlF2yvE8a7HY
cIUO7Tk1C8nXNiDcThbPdKs3j1z2YBsSJ37kde662HrYBV0laG8TkgjozQhqjBOloDT+SU4lJYe2
cyZgg576Q9YqZtvUhWDqckb8FLuQIxAocRk7J3N6h1Wt3S+or1TmXrZjs2N0POfhFd/qTIniOfNs
qhapZK2DBfg7da8bKZqgvgMNeUiCWAuXzzuzp4iCHYt8Aaee0ks06qF2gvaDB93execHTjCt/dx5
pjBEJSMNOCPA/QePWZ8IBk8kmA6hwZU9/7adKiGvuhxhkM+CNvXdD57k9LHTgWHD7+TYr1naDHVP
YnKsdwfQ3K+faP5cXH+odgw5NKzrbxS8XcT555JyEAz1HK5Q4EUvLASJueVhwV+5+dzxreo9fcLx
OcEV02U2Lm5y2UIa5FWNHzubHewC4tViloh5Rro2ZIR7/drrTU3H1icOmCVFF5K04Ggt28ddcHw6
dA+ANhQ717HwE4uVn/CphbJ0CNM+U5/yj594POyLz+5C/Et8Yy45CYU2C7/nf8UkduukaQrbqrfb
FuoGVBE+I7cWjldSYXY9bxVBgPSljdHXcs6Hd1JpvP+mdxxfkiUIGvGI3RVYMN9rKMwMWKsPkG39
Y4hCoy6tlgbAQpaGNLpk/UPvcWLIkx1mbFheH6EKY77hXqBkl3cVoEg31oTqLsHugl6ecwm5yRri
bqg9Lbd5pAjFMF0nxL6SWLa9O0cPc0hiFxw41dXYhNS0Ru3xO7vMdR7WFkOBUPOcYGDtD+DUFCBY
UXEZFqc2UA8iThpeRuxVg5YwRzzWlEHcAMrH+hJy+f3DoIEDSRXBpgk9lwAkvIlcC90ut3d5Lcz6
U4hfMUQwnJpI1dY2zzP5SvWtIbGMN2tR7314QXIqmZ2rsesp6OG9U8cY9wTL7DJUosl4tnAq13no
jOfKGqoCZ/Gmp62+MWf/MboxqUAA55Rwi7HpDI6q9FxqpqPKAcT1paIiHE88PaI31KLk/wOEGO0k
`protect end_protected
