`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NRS3DPXartUDU+iZHQDisAOqHrOKFXwuDgLVh4L80bbA8lfCQPL7g+5y5Dp1zyBN4zr+e2hrBAow
uS1NyoFR2w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BeQTx0EpjGx09KANltTxwfiL18AItjnwdOxN/7qujRiVSuHatL0RPsY89R5bHUxxn4RGyOnCprcQ
R61CRVx6Jny9AilBHJwk9mf0cyeE/j/H+fPHa6TkzCuTKbL0A4LOqev5Rhr/bWF5XO7GwsRtsp6u
XFgqdZpQmZ44oWjCfgg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DdhGkDMxHglc5PApnjiMFQ0No88ipaCF27PS3b8FL7IwZRgHwiQ2kqJxfXqdlF68g/Qr3+sgP3+9
a2g59PsiW5vvOX9pyljXU0INuBpU3kfcz1xnx+PUuKYwDvPDC9c4Jus/DpFgcwcz1dxP3gHzMPeJ
MpHBMAFTETEllyjov2FOjiqC7pBMBVjyvlQTp1RNHklSjfmxBqqKaLXbQsFz5r5gu0bjQRl79Q1r
ESp3H+TeVflcDzZwCQDRsZWOPYgLfIkcrPA3PKe8yBmdrnrMT9gqs60tE1He6ywAzbFZA9L7rMFr
aUOO5YxCrlehBGqHPAbpnO/3xpkXnY0PofQ2ZQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ofmGOY6xZsFFWTKkNpr3PfpNxAGLwC4eBHWwyVY0PhuMtESSYHqsnp1BwoV6BxSz4iGzfupWBG48
En3V4t6FQvSwFIUKQcoQL0kznfZOOlp15Bzd7R5wcBPl2Q4kEsoZC3hEOoPFg1iGeTNBxdItV5rv
hNQgJWJL5LVWSG+Mxww=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iPXc86sHm2HuZowIe0d6YPB6NxXETDpsaOzf7rsoRp0ch5fcbMk1uPZkFCzjUAz0YRb1paPEjheY
/orr8JJJjbrHizeu1wQ8AUYoVPV6NiLGZ1a2tCktEghzKNQkAr4SAcNSy5Jn+nK4O2BtI8c6PuI0
b3lgSsM3tgYDawciXa6VU0XokyaefwSxxBh89Z2u5O7Ew/fn4P6Gcr4IdsCSG5HNKb9pgg+iTTJ5
/4BLg+sTa2VxLih4XxPH4pWsh4Z0EEnpVqI2Bz5Rti9xFgecgarU0gqjU6OGX+KrtVaWlZPqYuYc
dqss0vJS5GeHzF/uRTRtXkB6114rzCqoEQJo/w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5616)
`protect data_block
ub4pWMLtkSZVL1+zikFsABqciSxTcG7Kz9apqUp2+mySMsET8IT2UHdvg89BHWqI/3aviCnR4+ef
6HOnR8wAlaztN0J5JST6daXOvHvwaYJYiYu/uQOpmCsQgFdWjv1DFUuVRexLT+WTsrvXEkFZG2OM
CI7l91U2clHmoF+yuXO0QquJPj09x9rZr/A3G71HjlHq/wknD512WexNLWq0G7Y1Ph8FnO3w6CwU
WoktbCYhon2B4KAj6yPFi+42JKwVTR/mEhutRQBXEjLcUlZOaJARk+WqLdNbeT7IP4M1nX6g87ZX
SIeUn0WlBjffEZDiZ7Xj9bu328EuyXrXbVBUMZxVWsYxdWazpOPEGQKPFwhhF5s7CAXAH3i/K+1C
7RpoVysO0Byo+yFSjcN5CL14nlzgxr1MmPNN8rsWAiwWZpzCe2fe9suK1rvgBOcY2iyJ/ZNu69I5
lVuh/pX4GmZXqI0gLGTCeYhtvMwSXD9BcSKPPvdc42HBv1UlReaYWq6jgO9PZqXyJVVC5gBJJI/7
2TtjDfjdg4isfpHPK/tmfuWxjGH8DEahMzkchYnd9EGMDZ4UR+zmJw7KKwmmfAA3a1BPKkDq8Q7P
HBtwTL3I45zds2ElJC1BenEbpVGIo8a/uePwUeZz3Bpq6mIbB62Z4QrfRPbqwmC2dWryykCqXhEo
cQLJVDBCRMVIYINRKiP4GEmKxt9C3z/pQa/8Jc7KaNWG1ZTWZVjwgzR3cxFXVGaQ5ZWLQV8el/BS
lY0So0TbZ3hcnM6cOUeKKR7+qxuxWPQYwEaWSMDoj35jt+Ct1hCMdDeP3jxk8dYNd91SlVOj/ejT
fC6a4KypIfPdP53h4zRHpR0LxH7wLOijrsIElMomO9VIxhDGQ1seX0iE+a4yAODyMXjAMY7C6OUf
IH64vrGvZ+sJCf27JoohGe6XqOYahUFO1FKcTEa12D1Cv2rjQxRJ4z1zZo8MuxDAKkCGJvoy6KVV
Mut4ZaUOLDysiRcJwQYq5AKB5E3rLZy15r4j/IF5ZyyA26tgUkB49Rx0YmK8qjkiQKU4jrtbIi05
JztMTtF5DaERdkz1ymZL7pAQCVIsBUOuci4BndpShZAd24fqUztQoyr9GnLgxuP0D7R9SmVeYbT7
OkkvV8+TBaE63MwxDLQNcuzgZoXnoS4X/UXKB5GCCli4XotAsnq6E3C4w8uuJ++ehMBZKBtDJhph
ychRZ34PReb7Gx/HvrONvUIp6Rka6F4V8aWC9Vw6Nw/z0y5J8SmkR2W5CfRq5Kmsb3zcB7pCf+Qz
3MXfIs5BXzxMZ4JpKitJgSQSrUmrEYyBJ2rNjE9ht8TdA3L2aYWYjN2DXA8PbUJHWke6jmI4Wo06
Yjoh4bxUUO9owwKq2A2A6jPYwkSMzMeET/zjq/ID3wbVrYmTH16wm1TG1h8KbSxuNDRHK1ErYAzU
hmY4ghTbz0Dw6GnBxEaKjNt3AGtcBNo95IbrWKZwqDuvUY54Cq5KrcTy/PobsOW+6HxSLND4kHCp
HO1opSprYHOYcnZemPMqLdrL9KFvOM/2Z6GZsFKR0nTFo2qDQLnu0UDdo5PQth9Y/jB+FmpD1pCe
iHECTTjEahNI3pe/LNcUItY8wtvamyYz2ETMukTSo3fxkkoRLDhF1cH5V1w6aEjedMmBCj2vv0OF
nZCtsuGeJ0+zj8fm7/c6g1j7SGnuR1nQMytAwh+2g4qFK9OFFg6dRkDHCO4F4hfRh4+OA20oYDnM
Pad3wjD0ErW1MgQFS2jM2X4x/A1hInlskqqYnQnSnenE7GMlxSaOtVUTzULhMSxf/ToiyqTwBX05
BLe5wxMvMuRE74NliNTjGSJ8ingPHIHFyyqxWIc6/y0RNJvNnBrj7BA9goqscOgPAiPnA/gDIsWP
1vmwuLi4nO3aPsueZhjnMhSvK1EQ2a0ylwWv9Ktq0U/TQizXwvMAA4RC7Rj/2AAcvMSEQi6mxS3t
LOBJV3Mo/Km2G6KGZ6nVmPvDxqsQB8bQVmP0L2RZpqTNqiZZTTRQXhcNR0Hwcf52PFduMa4qwxSL
qA05ndQAbsmCi/HXUoRJV0qNhzAdNolwyzpGOUTbgXcqa21VDCvdbcZdBNJgkMKpqnH9I0+sA37v
n9o622X3YbyYRc7kDZ9xTELFmecE11vrW/+iJ1SuDtSoKC4eZ/7maCqwEqFZP8VqzbSGx+duGdIk
5UrswstrniHcAJmCuFZzzys3m3yGMyhKryt7VSS52L9ygX69S9BFhkOGZqUkCCMn70E/TQk786l4
vdplqF1knVdAHQAa2zdEcJ1ZjKVdGHMRKXzvPL1TFiny9VkZAur+UmMlkFa14WMb6wWHYjWOGwjk
d6CJizi8oM/J6mHFBSw/5d3dsgS0zs2SUO5+tLdlOzu2ZFk063j7c3gblGUkr5Mol2k8CcsuhX2x
dShVmozZ6x8hMSHN7q1K6JOKHkuWVTsG+cfl1P9AjJdqHFzEw3P2fe0OWOtomeO8Psin5ZNSQvnj
O6uTRwuRBRLmEJuSVb0upWMJU2reCsW7WZqUtAJtozG12x8QaMTqZKIRONkPjTNw4rVI1Uv0JJ7e
IxJCrPaorX71Or+T+SyIcbBs9fBWNx1bjlTRkkEtfepi8kxIGZ68sr7Rb7Nrao5qvDdPiJcU7lV+
+60/OBbfw9rYBLt7KvH7hX9JbEiAZsI8je5Ynfd+4gPEaMsBlcqv3DGG/tyACPRAd/Il89gKzle6
9ShZMs32nu4CMWEulRaEl8w/rZ9gYzvujoAwbc4L570N85mmlnJWnfrsBZbG+GOLb1slNhJMZcpb
1ff33L259VGDXz19JPLnzTZfSW8wSZ4ZN8Y9UGIAvxQwsA+QtfHHw1bsxbBYLnexoDsvQcy+xdvS
+KYt8SfqrK63qtN9F5bMWpzz/7w/yOQ3z1i0exufqu6TKF96TLL6IxORBav9z+1P3aOi4Cxy2xvs
SkhGKpzYqEbRiMAiEhSAi3bt6bXu5Te+PczVI8uprbaj7NAv6Wzcx9wPH5TXx0gCUjIHG3G5nDKx
M1sZo1A+CIXqOd/XUkfCXjegNDChQOoJ0GxwqgIap2VAt2Ge6NJHbR7GTo99CK0vxZZrsdJxoEem
th+TExrp/FSjUixgVb5JjQNA0JRx11W5JujPRlwUH7PRmc0GQymcQt5cguQhu2p2UgFynOP6Av3F
mo7Q+REuFP0CZNb/tqI7TdqE21iWFiIrQaJF2G0CRBTaa/5zrJ2NzQ8kozEIq00YO1R6Sw3BaLio
8qQT/HZ7ZmuFO5kLuHZrTzGyeSJuc80fAJ4/1Z7tvEb4e+MVFIpsx6FSVzvh/zPoROFKh2qYy5DU
B3p+7nxUR1kWazmZ/DY0E7YwmBa0bqfPNDbBnjRspSn/bo2WRE2IZ/CJ4EYcnUuFjqXthJtjXUV4
SM+mFha1INXA3xx8EhvtGy6XksCg8wm3pfF0r6TYHxkQW0J7/Vx+8ckvkks6luaP7RarXiV7MK09
ApLo/210m1rxILlI71Wg9UGUJtF0AinAtvCo8LU9toKVaCBnlHthu3pT6D9z3hCmbpqHF9hAnFXe
sj5oCsB/i7ZHz1IJnx2cnUu43gAxVovNFy6QsyDn2RjqlL3E1GFfXZqtggcMTWZn+OwRdmoKNqM8
X5uRezfeegJs9keMNUmx2ud+uNfEk4w+9GcMkKQENHg1A+27lsdTtjSjTfuaHAroarprDFJ3Urdu
Hu9sFPWQcAtPpFOqcQYkziHlnYvWHHhpP/uQ57Re0Y6mYBiRSggHaEichCP07eOm/wyMJNmS6/TB
XKryKygjfa8LWg6e20wveTIAj/ysnmu6zchMuolrLbuSkCyyqit8cFYJtntmhNlr6kpfQL+acE0k
UBTZjrPIYnKzUXKFcDis/dByioEm8f5XuZCOuDb+Q8fEd+0pmxged2HX9gE+5O+s669JiSDYZNsU
bMxSi8blcY31lCze1xd1WC6bfLQN+K+RfgoNErBQRwts7VkiArtrLc/kuDP3JB5lnckHmLGAfhht
U5jt0R1ArhpMFYkbGkcfTpk7OMa03cQQeBXOVEqpa5GlagvMlrsV2/QU8qNfdGd4Xm/sKEBVnvtK
UnWmKKPeD+avTreSEjWsXeqrUig6TFcBktvoX5MsLze4aKX/hKpvpVIP5n4qShAif0N8mfF59D4+
LjjHCnV0/epMAfKMuDmbxfgp8kCwMIk7NiRwHOHnPY4SAOELi38tdyR2tVhbegb7Nh/ez8Og7E9Q
fHccOWKfsZe0fqEK/IMd1a6BPRlo2nQL1Pfse31jS+Dud4SO4nJ2sEpgpKDsTUrHkm57Uk21FsvJ
IuGB35bTpnSzaK6r9ZOIfDgaeGTWcLiLc6LK+wQymJ9M35X1qdWZJPg4nRwQmqhUJ83jX8MeEQFe
zJoqhc2JMRcexZ/LSRH3d6b5BZ54ZJ8ahKWM1eqGQ9SQSK6ufrFUJonJhJijZlK4oaPnLa5EYFSe
+GV//3D7FDPaIEZARsBo5mb2thFwZsyPRRqxKdph0mwtIqb5wGG6T9qzOT2yEQs0pYgXerOUDCCf
d2MbZVo9Zo/nShPdP9au0gTQ2OUFuLeaLRCuNOraDCOhLs5cuIGU4jom2+9l9NbxiOdrH3DTFN9j
b8oWnUwc+r4gk9K/fvVwF0xHQt38AprHQHVRta55lKU6nAd10jEuUpVVQTQ2PIEV5V7rvMjLonTN
+SJyKXwfb6yKgCjloTvOV34AewiBqbwNz9Vp5/7LjsvWWob3peRvWf+cUF3JyYTtPBvUOWreT6y5
C71erCtB6pJ5BDeslMTyZd7l2F1KBxUOMGJR6DWLEhPNfCCMqQq9hOgEjkBiCwpBmJXzI3YPULJM
8D31eWq/PT53FJ90r8ZsadoZddKtnNErQSW5XV8W0JXhooxjj496DDym92qtuqI8he7zoxU7HTC3
CmTAwLte0BflxvOpdNGOh3CvAGahwnbO0ZkWiX+zscune1kM08WNMQMPVbEKsxIpOJ7tVWpn63ed
0ZSjNb3XmKUN1lZ5Y3fqu7RqBuDBxBFNQGVkwFndgvawB4zeM4JfJzoTewAi/deVUwNsvGKzBr8U
c8953qmSzxLMy1lBWJg4mHZ+cgP4q5G2UD8/sY6JDDvSoE5tVC6hvWBiWJ0D/pMkhVGBg2NnPODo
GxmOFG2/ZEGHohNgDYCbEEkrx9MqsK7jPiWcfNSMGf5eiVchiZEhXPIps3+x71/fr3Q/2soi0yFC
K6Gn07Ph5UBeYNhEWVkTObZARK6kpPOORjZZpggZeOa6mEZ7t25JMT3nOxQGEDiJBZew8Z+3Ae9p
PYbqOOesGvWBJ6z7ADl4iJ8AfZzXlat2D6CyncUdmjd9wGwsw7LxEVnVqI58TGZN24x7fnZjmDGO
mZwnPPTm/US4vDRPRvvO4Uvvju06Z34kPRun6Jy56uss/pgqiNw3dRqJBvnMUwZ5QpO/yj70XQ44
PYbiPxjPTA7ZIojUMMnzjeRVV2xNkYs5OWcFbQCryabMc4KzwVjtZUq1smj+9X7y2KD40m0Mif3z
rJIKYDtFrgnULtKYSn0C0KbOsh+O98LFh59W3Ojk5kyL3onsWy2g/bmss5/BxFLlMsxy0P1jGRik
oMzKcF9JIlvIQj2SjX4dsetZQ/KDt7c6s79ESnwKnJo5YjByAH1z4i4/ljYmwSM9NHisQgAya4JL
DlJ6j0gQFd8sHyT2lFNlwNf7S/r+lbVCpw14B8Uf6tb1HE1dXyDQylgKJa0g+/aHHNo0deQxkMnB
pmV7LG7fO1pj2tEdgPIxcTqybTSk8d61HfSuQITsLcqPo2C7NfQqSHQrTckY6Y6SIB6LF3hSD519
UxORpR4eALurJKG/+25TMGI1yYvZ+B/PKLWJsqAzemqhkQ2mKOqrnJ335cRCVJhurqLkeYvhta2Z
eFWI+C1T/154ZCMfePWdZONchPKzGh9sY1uxGPobCDDwoZeaykKCPDezQITugyZiJ42MV1xRfL4x
j5Z60Fspe+MDvNXrOjQteFIGdbdMAdBJome02KE7oNKw+I5vo/soiWzLq5cfmYHXn4HsUQAFtwAO
iYRVRK1LCpeucLQ2c2ene/6B3/Yz1cMwLmNOxdYlbZNhtvhdj0gOLgFOkxsY8P8cOcASrRRYXnd/
E7tjwdn9ZJA0FDkrnkyvrr9vrVjYty5rFr5dAi0YiVxpLoO72NSmFHRPdkCrZsmJhFRCkeDELs/s
wrRMMOraizLD1jiVHtXdesiiH7P72c1zXMWdRLQ/udn5uI++HH1vy4NeNxpfqUnmsF9I1AjinIpJ
d89Gg16ycGPIOr9PAqozzacqwacOULwKv7O4Knfx6LKXMJKfRBCRLuelv1QpWzUgvOhKZQ10EKXq
p7ha9h3ur1NA0TnQoTK0hrIisL+EcNAfOtS/2+kgvSKjc98u1RMc1+4C6HkmXuxg/+zGJTDaxnJN
NphWeqZvnoGeLST6bKavFIna6R8g20MKwwtTQSjhaeuaxXQc5HXppSDNTfHrmDri3s2JXCqv05ow
lmDkLW0pfFMfYJEEpR+Xc2lIhSQ/2Wf2IS0/bcq5O8fYqbg1f9gl/gw05h8FpzlTw3sEPYB21Hm6
ResnCQJBe3IIy0zS9Wt69OoIm9IPft4EM+ayr8fgAvjN0AsLdjiBQr8f68etR5ZIUQ3ozQQpWeI8
NGci0jzPaH0vuu6v85MSiCuzXn1902D2sYXE1V2lp4dICWG2lgK9mpGzGm3koqG2SWhPNFeSATZG
mgWWKOErh6sGoKer7E3TQjz/JgkDRBa2i8LMTkilpFcvmTZisVJgThMfmgxOHHE9DtPqxR1EDQYv
q0AOlSO2osX82wdQB979pptfst4kFgD10T0Fk/PG/ttX3La3WZhSMaZMBziD6CkUwEMxM4ta58/q
iX2TvmtRAuobhM5x3b5V8KFpQbZa6slinTwq85sjUEJ1aANO45bbkfeULMUTz2FwasZ3QW5vXIZM
12zmCDAhs9TV7bIpk3BQY073qsERXCfonQC0bW3HoLlHkWqbvKYi1i4755VaTwlzpdeCKnkrMt2k
81DEcePw+wG6+As3Wd1969MlKotglegqVE4uGpmVzJhosOTKQ+H/Ndaysg+02r9PdjhcMqNGwD70
9txpv5cXZNVQ+oFCikvxWSJodQiR5Nh/7B5YyIk1gjUDgrbYcK8ovzOGlgxAJXjFO+gohgPTZUQc
OuVXIolfmBQI0/UxgXObV4nmLvfUzAkn0x8E6mGjhzygrzm6CkhwAIhrNha0gDVybconoJ+U9xTm
wNg7f3yzpxmkSqCfwntl8LeiXdGqXQ2nrQ0Z+IJu1LlpEg6YU2FiHUJsqXZGXVT+YN8RUMFzimmu
PC2IdysGLBs33zgbW1RLXscrebh6F48rWedSSPY0Ek3bTqCTkD5RyTdlzREtdzDpt7A0dp6e1jCK
RUbGIXtrEV5jTAOiK4wAnsQZvSkucdlCYRql0va+
`protect end_protected
