`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Bd8MSgQR/XPHDbB3PF5sPKutlr+/c9/i4CLlCSabuZLZL62g45+Uk6g0xRrISr7Bw6sqlQ3U4BE3
llmn+zgZYQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
c1ZCWoH+srVT2mmQXN+E5PGMBoMQnPW4tU//hhv28z79rX5UbFn+I3rTKRv2K+wtd51qnICLQpFX
ub45XA9T8p5VXq0H8ICqHNYh/v3MwkmO2yEWWgqnzRoeNxPfvg2oBVfI60fXP61b0kKR97h7hsUx
5/HzZE99Z3IDjrHScXw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VkOj3vI5Tm9ndpUhhcumlaMml10WvVW92l3FRMoCWb0mQyRMYwhSgktN3+qQhK07VHhMYq9MErmb
iSqeFNWdk/q2el67hbY47R1MfvRORmQ/iGDVXjHLfSlsNhYv7DcKkZxKB0sQRDjUwi7OBHX26yBd
/5ZWgMDYmN0kqGtMpIhGxObvS1uN9cywnZb3wPtaKIGOdsAY3hPGSH8IZXqzgOZQtoj1Xm/qjQk1
GBO16jaozALRIvuXZrZqQplECaL3YJPH441w8XGGJx3iFEqzfHhw7TNewIULbhAZw3br7UoBKdTZ
vSiZOd7b/7FPHReXbBhIaEhsXavLpyKWaqH3Vw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wtzqZvzpvHDsooUxvWnOfSX8v7+RJ6Y8Jhy2BSWGcSQMumoBPqwQ1xadmJQ/pGK6M3OKsTMBdr7i
NKJXc1Klf8ZG0hXEBISZIUZkIg8xjGip2KhrjQgXzG6STI7rqOdeHnk7ABtRNhEaO2PyI5lbztO9
oG0BAnHrZQrbRMZNVrE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rcYLK3ltYgsN5nBw+3OWoyp6RBDEcyS6edNP3tCS53rOqaST672epztJn7XRWf6zue/f8mYjnaAD
sS7+xn4tCfnkRYGKF5uX+lbyx3tF9UX69u8UNPTdaWCX4qn0106MBSKIbXEaYOCw6A+WCcECw2bU
AyD0c/+JAi+zu+jh43Ell9Of8huR3bY4+NAg/q+E1zhnzm7qdwGqZ26XBLWM1FjNNQqlpaGsNi9n
g+xyC+p9VydMYlj+76DSZl/woMYQvifmHKEXlm/FqW4XtpDARgbNRtCeHuqRdzy2vFQrELoVgcla
bIhLm/iiFYvlAfNC1GcYuuf494s6qHR6Y1H06Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3248)
`protect data_block
yssl2r+Hshkb0/k9xZdC//AK/amyqZb0qTsXK8Mh+0G1RV2NYRM51xzvSuT0PiCfc/eEKMbVqVM4
CIztlUvknQCze2dV4POpeS5n1EgqIQ3rcBKy8vYDDfwjnw6W1q+B9m8BwIblrkc/NI1pS9O7HyEs
ZZnAuB8D+7wCIfw68Y+ZHNS5P2wt7jHCLXGEjZ7cRyUosqejUK/pSLPEgNGqVCzZ4sukDxrY46dV
RcdtqtvU//SXi+yMjYFXoD73iPv1pbPzypnyoUab7o8UtCl6rimrNFvqf1bJ7DVuiT1n++GaraVg
I+9lRlotUj/w4zpOK8FtscGgKZowQ3EIj6vtMq5PXxo5r2A6f3m9pxraIkPxAy82TwbmDiP2UnC7
EzaKqn9WbXzviNIP05pVZp7msWQs5WVjlAAl1tSGW6Kh1fnnQ4o+EoBxlmLme3v8A+tPG6fKMr7m
k1GkLkmI5NrqCloiu9aVYFkB4TYLKJ2W2XsUIkUsgwyVCs/CK+kzIEqySbNvuvP7bhjQ/YWXHz6/
IlApGxnf73Q+E/iL6drxXa9TYMSpkz16J76uQe9USWOUwAc4QWGGk/nbu4WxjbIGk8TJ4i2c+YgN
k+xqmMjYcUpIkPw5e8IkhCQfpVd1qoGwg4O78YMWXqSXbeI/kn4C9OlU1xYs3qVUwHE7Q0M4mnaQ
e8Zlb0kk4ap7Z7Bc5HYLfOXMvXutBHuBwlTZM+GxgX24l7V59K7o9o+5YdxjC+2tpltM70QzCqHl
tEplh5rSVfWvK8g9yA49S25W/gjh0QxbQMADl2gaT1uEkxIne+Oqx6xRXBODwkbmPA+xnMj0yrwR
ypT90Hth4LlRRSuVKFN6ZS9SdJLnfv8fJ2Qs/HdQrD/5fREwgLMhcBNHBaffDtP1AnvOxXsIzxkf
XVOh2VEmIgHt5QiaeDDSTsDDbXs91EcJf6LtUWb/8tpdWtQ4RnxbfMyQHp4LSOsfjOch+NpLanLw
TjSNXHUE2I+xL85A6DTzwlMIrH70YMWndwxxXYpyP7t24E2+yWDb0pVUXsP0moseQ7KarHF/ToWQ
LMeP/3uZJWG7UrfAF2BCQvOgJgzwRRF+ixewViusXcbfil9eY72NQ/DWjGhhF3QdKgTDtbKuUzxH
CiW5TpaD3WszooCIR4D5tqbISUl/HRjuEQ2eorboC1oxDQooeJXjoHfMEN2KGQ+99v8bCAeEMBIT
NnJ/QH8PyA2SytFrsv27u5lISIBw9+f8z+7YOKbwV5zsvjyq9iLUr1He8ZvQUJtUSJ3tRxqKbhPI
j4Zxb49yC8BzfbaTLfyPdOY7EKrRCBvN3POgUvcaMRPXKZKBTTF8DZcs0wv+mkUWs7JGMPa5nmka
iQljC7FHWOzbv7EwzUdCVrcoYdxlNui1gABqyYpzQ89ysGpHj5tMddeu0GYq7XWROyEt/Vlh/4EI
wDgpnHR7dDIMLwKEUwrV4klQg1Z08GKwRgeLK59BFMdAQtjJuBdbSG7CmYD1LLeIZJIxk3vHlbNW
LFkLUlWmRfSYgqTJvHePjKSvCdAHsBHiGR4kzg64BPgZC/tLqS7QXrbVyOqKakU2z72jlRmR5tyv
5r7m7DBIHpGmBsFbwhgc7fgohgzXFsL7WaJZVrNHf4PVSTyEOTsLjmWA/UzpFs7h24me+Cy8+WmL
q3r+nai6KU3aBSwWXw6X7M0vZWKb+doZDzrKHXqBAblKDCADC1cGwIFUlDQFmGBlex1bfAXqes9+
2MdQ0vqIH0JdsghaLbOnfDWvPu/sW3Nvxdzk4botSjxcHMC5EV6gpjm0hprl/ianj0mdbdx3/R8e
bOd0vErFSNFLS+fCo59NCZrtDZC9bJjS6RA7CuF6lT8Og+ngtlg0MxldeA8CeemzF1ZdgZ2Wfnqe
f+08c/SW8RfFWknysEA5qlMqjeAtUyIB0K4beT5Ix6pgjxe2VKBLnNeBvoOMAra99sf5y7SCAP1H
NEhmu0zbWOIyuyzByVrZfGvbEDrn7iQvhDx+v0A7XBHBvDlZADmTjAKtyamqTLfoDa1JjX81mAYw
dYjaoFonVYnZKkcfqm4GMNWIQ/Uxe3loc0TnsqqQhbn5h7pRi7x2Y2lVnNGWT0OLCYvVQ/08MKgG
NsymrnDuyunmsWIxWndf/qdbDGKs0Pt8vEbJPuqjxF4QfXl3tzg6oxVuKw0X4dHIdapvS0ydPG/n
EGdsQDOZWc83XyIGloYX328fL+tAdDkKsJmEYKAsH5ws8jeTg+YxWMqawmah/5FMmBdvwf5Pj19W
18fTXTKSoAnY+FnIiYd3MHnOPaOz0N3P1wyGKZOZk4RCOMflCKI922CH5dluAhX4PKzf/NggHg4t
y0sTwbEQzX0zUPJywSzoUiUF6oyTKsTytWxxl1Bf0wcrOMMS2SQrVfFgLEGYvxH43Q2GLojgln68
aJWqvpRwlyRWbbrFHlZGFjYyMq9vKkPeDut3Ql/bYsNyMoiBHy59q6RXeexdBPR2iFZH82BdIle+
pQ1OZed8m5RNJti8Zu/mp5J8lGkqfVdbWA1fRWNiQ654ijarb1yg9HkUMPmwBwgDUq96q0xfks9t
F48kcs6HYcKv04KyFPhp3kltN0X3tnRwYxBAJS0S+xOVzKGQGApg8Zso0QWwQD7helFgp8n7n8mF
WeS2qN7Kk6561CRW1h/TovQwF+EPQZgp0rHsa9BaIkyxwqZwxbApQGAu0ZoJbVNNLRmZL+1bI6qs
FmtPVna1PimmUrUj8fD1CP2fODtxgUX9r/fLoCdo8NRqN3ACnThDKjQpvArJ1K3XDDW+oK+w/xH9
2dqf6jhLf/8jFlyAdxpesoj8Tj9LrUPRUa/U90eFrWE3LKtq6advz2ubB8ypp3FGsOtTmHzGHMuv
qOcrIi4/TjVjWGeIM36A14fu5wltoh2yIoTb7l+N9jGhVInkpyddXqkzwdvm/CClENfJLynNm+gS
LV0r/ZAlYV2nhz/WD8FCr4d3zjqmBi9vgMsSnPw/mgCBIGtEF3wdU0vZ2Ub55pi5dS5iMT0jQ4t6
LQ36ZAK3ISUy4l8zwxy6ji4PzyCZ0650bnXb9WWj+qBj/jh636m4Ezq7O3q1QlmnAWOsmgfuZjdY
RAcWjr7O3thH5MFG6YTrltFaWk9+mR0QXSk+98EZlfk3O1ocAzxT5eRYXpbbjudSx3yy5ngglU4w
XLyxUHXosIh8V/mjgAevGMS0du0s84Oc0K7+QlRQpKUEhep4BpIu5y17bCnwsasu5CS8c9yEgzB5
/la/Wq4B11lNUIWjt2+jiFFjUWVOmtGUNVSJSDym1dkcFMwrSL5ygh12wUbS3ysDcrTdDijB+azb
MN6UIKpM+Kg68wDeo5ZJxk5RXarXJGEtaoJy1w9oBFZ7gRPBQRRfGxgNMIzFfWSrIj3CrIwvBTmx
GCTSGoYYiB4td9zRiM9dRjynpF2RVvWi6zDKhkJkKKW1N4dj5PnUBHKf8NEyMdvR3LDdV9oF0hpI
BsoV/K+GjdoOhSoSjtoQ5+3t7VCvE0ogH3TwGwuJXmNqVQHLt39ymnhHjHgkS/2IwqhI+jY3NvX1
Xg2jdTtlIXMDvPGdjzQyUe2sNFKfil3Mf7Zyds9fC8VDbpts7JbqTAA+UxZmJ+fhUBhgJLnasGK1
128W4sViw89+urNsCKK90DCY3iuoLZRuiSn2z/fSIeyhP8m+X6bghGCdKeCO2UlLLWpHRmDfz50P
9k+p0t1oGy1m+mnjeKOb6iiKkMBm/tSkQkupb3iO7iZDbj43QRWUSr5G/rKQqYDkQARaXW50KPAE
iSF68g8Efi5nJ492BD1JJVw71VObDYURwCKogV+p8CCSexyapuFGLnG0q5lMZajsENyU3++2gb3g
3jbe2fEfJAepmjXLrkUJuoZ3M74Wm0Si2x78r4JnQ/j0QNRLmsn5+6lLUsvOX1Z0C/dPb+Lhi7bK
cPZSLFcLm1jJXd14YXJEccjgPM2SXRO5LQxwjlYzdRXR/lEtCScb0XHppYRG/smhHoaF+PGB7jxI
SewBT/tf1DOi4FCM2jjnYZHyQpnf1QkXW/ABzRAVn5p0MXifXPBsXYgL2Qa+Jgl6e6NN7RAZYojF
DZo5kMrw7CzdNGJxHVl58hSob54SeC8hQ9l38MxFEplAtik9YGPOeikxKezMnJTtqyVUQub3uwgM
pFwY9WwC9+XIgBEStlokO/XjeLe9Nzbq5bgp//haii2PYZyvHXrnXG2YCJIkZz5WqbWIKvLBUz+I
EasUgf5V6J7dbePH2CfGQdMKTebdwazx1nfaQzB0ITiIKxskI6hM2l57lwNSCxtwBey2uDjCuM4=
`protect end_protected
