`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fHwnat1q2UM+waeDfU4bELJ/BSa0urwgWiPCsDHOP5MqNgfSeflMlseOK/ZrzslrZ1riBx/PO5tT
H4QVkW9BLg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NSrO31Xr5NhLS4JU+QjgBRO6jfbsOmudWTGFb7C+Qm/NHUcAhOFLhuALhx39ihHm6swUodhMArfP
IngvKAEw3AZ64NpTReM7lahCtgxxNkYRm0JlmBB+qjgqJ2fyak2m+3P90BfE4rnCnJtQZeeyRtlI
H0RP6977FhVUHmMAx7A=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YcYnCRtAcoZg58QbzCFwHqGnmiKFglP7FblMBLA+hnSGXmDTdJvB3lVAGKK/e4s+GFe42kb5gjNh
GjpwIjrGP/9IOaaEgSnmUFFXgWznJzPO3xt5hGekMR9VRh4MX6T4o27jrpd9pc5FNe99/jJs1cV5
3A4UJoz9CvoPxC9N+1JZyNsXlFSG4k0edbNTYrq/k/no0P+1C2HssS6zl3nb84MjTk1cOGTx+4n7
PIfjqAxMmju3WV3Qn8jtsNFAkytVutwNNr02EZI1EXfDYa8YsD3OjE5E3r0qZ34GCCVxR38bAmN6
ngmPcNDUWlU2znOG4tSygHltIMUe7NHUSZOjWg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KtMr20mQKC6f6IxvUTv/aIC4W6NKrmmsaPz+HcRrD3N2Sus2oxcE6RzHcwBTZ/RWlVbHB7HSvr7Y
nKMqGLTe4Lh1/vO2rTztX37XyX8GtxJB78cluBoOeEsvS08thc4i40JvnUrzu6tZcQjJE9clutwV
iqKuz1NwVLTzVyktoTg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LqNXuZCn1Rm7Q3yGzPJiE+/oNPMocLegeKbCsa2WEGmAQF4rxR8vG4Gvo07vPH5NtckIS+QZKZnE
e1GVVcQCYVBL0ipecqsB3m5Q7Sxh9om638rsI+QaS8cwRwSdB2IWLzE7ZuCA44cuSdQlHD/4DQyw
T1X8XzYgOp3GgL9ppU1JPjFAndMezJytgRBBVdy1p0Zrc4VfQ9MUhtZDZikYWVXeYuMNNFTikBbI
Rscypn39y7xqmV0cQJ2dATrIHNW66x0bVCicfbWr4N6PI7/6cu4YN2AAZSBHO3kku3nMam10xn5q
dOK5kA+QfRtskl9R2aQnpeC7uZ6x+4IKs/kPMQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 28320)
`protect data_block
OxJ/A/pxK+k+3xJkAm71yaBReofwFTRGqZNvgfTj0B9yFu1Vle62peEsORDRaNc6DYDf17ZzZtF9
j4EAvyvSMEHNGYxLs579wnDwqy6w/sY3Kr3l0dPQvRcs89pQtIQv45duuIX8mZvEInPflgyXZ6v2
zipymQsiz7TBfOnoRswrUysJXA1tQTF1larPZJJSmCSxnfbighhska8K3A4AD3haWhYxLbUqtgj6
K1TpmlgZtBQI0QX5Q5ZMBAFjnVoP8YgLcrgMKrBGM/6wFvhTrkn5Z6roNg4a6arriv3Wu0G1Diy8
tihvRUJCJ3QEBUrTtMGN8n/eFE7ecrRYSxXZfZSNFXKhFP2rd5b83j4XonXDkhYOhX7sXf7C6gxJ
tgjpQofS3gkMDJIBXTIhHOZzBYjE/WShL1bI0ibI/COzU8voNDBQtIET/u71fUcKCDE/V1FcHPpt
i+N7C6TvjICyMBeK6vC2W22sV95aTwbEXtGHillxcQP89McGH7XNgXzJpDiwMmg6ZWPLnwsiO4Qj
h9hpJ8lTz/vjlhLTdjzsf7tMJz9QKOqmZMZPXdEPktGgONrmt0bFONMXDuj0QYsizJsqF/v27I/q
DXBZnNPdXhbRWUquOU8cdgyQXDou0UUFgCgqrM1mva+qDORspJfd+rNL5qfKZJmzqIfEltEg0W/f
59RbqMEBnBGIhfDNMJRyYyuI2yMJ9WrmkX9EOgCDj0Etwjz6EPDi9TD7xgAoTb8CDjf4a5aa0X1Z
m97ihoUncQyUabVurs9icBHsRtSMBjoWnkIOMGoaBYorHm1MjPfbIyz7DYac13nRc7MpGfVp5PnZ
NCwo7ycxhbbD/II8zJvgyxF8FYg+5ysE6Pb28nHlckMm1qw3xd0TN7rE9NS5wvXg/ZLi16PyjoXe
3LojKJQEaCu4E8ztaDWxEWRKiesG2EvMtBzpV36ub/mgOEHV77FEw42o3D9aMbtknU26Ehy1IPqm
WwPiWjKf+/nYJeM+nVaiTnzMLHfRvHNQLe0S34Qitqe2RyXM0zTWF+o0CD6ywcM0MW/WSdXvKZJJ
FO0xjDlZ/vaIL7l6hxMb1jOyt/8aE44X6j8kAdIKPbJMdIjVOm4+VjhE9XHJ5rKecuUaP0shLInf
OI+UOgSbgUVEvE3kF1TElVQrW5ZeiyEq49fV4ON1qnXrYjiFJjo69ciqqOrvmAgpt0VctUiYPz+k
ZIBMDnj3mWbjku5B2Ckhr4FBaiQaAPmd2oI7cWvio/8H1ZKdJ/EUR2uA778H4iF/6+Iz/xSXXjRU
2VyK9dRAi/Q9IZTLmzwITFeebg4jAzBb9JlyVffG5Ec1ew8mge5Oi2Yj/sPW7Kjto3vX5cjMiUrv
VLdpLyUiFKEH4NaxSHAzz3ASK1Q4nBZWfimDrjNHPapBkXqNUrUmGCHSZcSAw3vIiMEdi0pqH2KQ
4Pv/EIPG/g6+76n3z0zrsrim73SG6+rb/vUE/zlF76jygo3/bD/t5dcjW24PEim35k1FumnPNe7q
4lmbO8c1ytRbPiZW2VIWJ3KdKc+bHLdEn0EppfvYC0UatQYLGqCdwhqSq231zHA9fN+IzAriEcSm
bQ9BPwS003NtndwSXGzcBJbmX98XNOyhW4jQOrMTyMlxavAHWlKyyt479Io5+qlNVWCDyjsNex9n
rkMUHnn8SoNMiWsN/QoIe5OQbUHbx9r6TPCdan0vl2SfJ492/L8W/4hBrlvPUSc8mCj45qcH3C+G
h2eeeF0BPeM0O1ikYTfXD1Ui2cRMgXTYmxXwi3S7TXPZkZKl4SFbObGBg+4UXW8kSow7DmyHsYa5
z+gS80jIaJtkFH4yKK0fRIMs1x/gjp0gkhKeCaK5PnCKNIJCs+JfoOh0OFW/b4n81Qrge22JauWo
+FikgK/zeKS+Q4UaotS42FPMaqEgHdohay2ar6KmeRnJoRUlrsQkMN8HMFSkd0h4+NHg9AQ9lXBc
JQVJKijvO4727GrPlAynPUWq8TSa0v3RkIRF2cVCmLj5KH8GzBUxxi60OepP6xA+oBOkVCJhIUw7
ZesLf23XE0R9QCezaMpKvjhpEZqpV86rWWJCfXUNmYS6k3t13q7fojz8iWCP9uCzL3HAOBXP8/V+
6SRgBTKZ8cSh+vM/kE/FKXzEqIUv1+jeWmwtL2TMJ1FyonGtSE3JBONPfNvNJevwcAtcG8v83BGd
u9wsXdSOVcPwWKPjxqhZRBBc6vTxuZpD8G3FTGodsXRbYZVin3lIaNJgr7dryw54jJWsOjWZGk6l
m2LGLAC9lm2GcKNH+Hb4VzmI6t8mkJ2U2hlleP/pCcqGwkO8+8LMHHbdDPvBIcVOGh8lmyORohL4
YD5S/E0WppJY0VXIBG1lHnzP2z3O8b7luWsNDhPkYaWn/0dOXw2UEirQQBzqmfNU0+PK1u+IMLKG
wBS7JSGxTyE1mmBj44fXWRmEhsSqKx1JLStphERDIeLugaAxQ7C7vFBFr7tchbERGvd9UAchGrO1
Jee6WBH7n9+ohjJ+GkS5tjeat7GywZZqT0h7IPqzF3tstfN488rwzViWB7IRXgRhib6kw0CrRZ0d
n8izhvZCzyChYO6rAm5yB9H55ntOM8BpguM6GPkcMPL20FCYjQsRQUlUDrZZpaZIsij83IGbCVTV
bi47LOYA70ANrcoFAOBZiCv9S0iBSVNrKyRRMdPX9F+vBnrIdJ2TDK++zlBjax7rkj982x0kmSGl
gQNVemVx2OhQ9j+hyV9xqh7cl8hec1vnfNf7YVCSSBHgj6CYPD7s9YiETyDomjFdQsLY4p9U5dVu
QGlT2IFKMNBQVWYsoMKlx8NUIYuI8c34SkLZozwyhzMlgWh6cVHwsv3Cp3UZkh0l3irOw+LEQa2I
c+5UfyzVIwhb9X6owl31vqLsxPrNtdEZZFEyZbK5JfhvOfiJUWZMoEyag3h2gQoJ6cv7joyN/5PX
tlE68LHGYfmjhooGwfHYuLQAs3QjeBp1hQop2/BGmxXzVOTfFKFBXep5Mg+9RTeY+bY0UgBpvQpu
baUpDqpDsEPsAXCBqK7oM3IWoJDMajhRec9XUNRBdAqJBhR+YLCxwtNweihfDZZJ3nkDIw95Qwgh
FuEwgVJ48aSE4A/trkAAytV9OBDZXVojcALksXh6PQqAkwnXBsZVx0kXjejbqmwslxsgC//mb0M5
AIyRB3ANPEpeLJekhl9K69ISP5Jv2E2W5F8DPy8GINRPn2HWNasxCp5a64+l4WILQ0MZcYj//G62
IqTKIskIOgCeGR17sA+qh04dzkHjkWQpF2J5Iu2cLPSgMfnGJv40WAH5oMQnX6DGA+tSG7nn8pPO
++Dq+xzCQFAq8Clu3Dhc1z7Z6qiHiR6zBdahn+yi1D7jt53p2Qpr6aKYVaOrt2Pv0pwVbqoNmZCn
8zZD3AUwgkLn6bGdMeHyqXA7h+SpQO07fpY7vttX1kP/GY8io0R4gfdwTiLmbvmdIvkpQYCYcH2q
uFDCthH2CeAMaWd7zvZtQ1f4fWzIWC8+sDBNN1eD7wEQndgTWui71F5eb7GEMHllMXM0CKIsZXPz
DXtPCZ+WK0ILxQ16ORdBGlNpv6UiNDRjTzWwv1EsBVUJ5nL3bUWDy8GWNdsJQulez19wNx63FLUq
6a8NkmKdsJvO6grXpFvIpQwATFgvd0QsdNqjjjz1sVF2ynm5vF1ioK5aEXpWg+eh2JT1XvWx5Su8
M2Dud6+T4zdPfYSbqOEBZ09j9PH6C+5p5wJj9ZsznRj+YYEmpZFLvZ8bZqIcClMmuhFrboCn2oou
+gWYl5q3P04Ue3qqe9MhpiSCsHbFJhUMg/D13ZJBzrKeuhEn+CyFPW77yFb835Wv/AGIg1HonMvD
s496UdrHoSk+ab+sM02fGEeT1XxxpV5X7rO/uGWQbRdH3HSZ+NAfImxaYMhS4yPmbqVi5AslcWH0
11xjvcMlAA0UYgeWJlNeJTh8t33cORJcVL4EA+dr6s16G7tT7QEcbn1q5XlX2SZV4S2FifzvAwF5
WCwhkZZJYMoQDX7myWUWytG0wjTyYn+KTXPrALscFJUmz13veE3zMOEUqA+D2tgwG7Gr7+hQm1la
MSBZFQx7Orikw3HB6JeM2VxEvYgUbquE7Z5M3fR2e+r7QvJUWdeJBX5+ek7y4U6he7ZRnjtQFIkX
6ZZBm84ATmCIP9GKKTfHErHFgynzhLad6V2LrO0coPZx20x77uHjEIWA3sp3nl9zg/gHvRYUogeE
KMWFN4wYyNnOWDCmJVNjph4D2EerUcXZbtyqwS3fjHzVfGWC+26k7t+YD0mbBGn+r3xoRWOo/4Iz
BRmFGbVkWuRuxNfNR7ZpHU3v0/08JOC9yzvBWk5892cNCm+3bY+moTLBrk02g8RXSLj6ntwaaAD1
v3ubHoj2m/3rLIGGJYC9Mm01/Uc8rWBPT5udbqZBqGork+oc0Hp6HGku/r+RpTI2hKdrOpCBfKy3
XmT3/orgvxOqnUhI84itKIKrOS394KW3BCRiaRPGghpsr6Q0O2LoNgEibOeM5mL9iyNsnNJijW0f
JL5ce6LHXLgyVhreBvwbFy0N6CNBR3HjDO/cQT7GjOn1ZOMePu9alLFVWAtlxiAbd4fnqd+yr0y5
o/2QQlwQAfkislct3xuAz6a6wJpnVS1y+mHY9p8qlJ7b3SlzlefvD7a8M4Daq1eFXfaVVm3R0K88
6A6hEuUpj3b0ZxdelrgDelh3ut2XtX9Avbpbx6R5Wjv4lt309gGGHQI6oGa1TSlSAM59YbqSuqzd
7cDElX34Wt/98rm25Q6Lhz58/DSFFdAEBRxoq2gmMtdl5T6dSAoX4yNlQs9Uw7kYSu1u478fAN2x
d1Zi8fs7yCee0n2fq6dK/xO213g5t88pIdxwJrwhk672sr0LaxopC2HOqDgBrc5euh/nmhlNCNO3
Ft7TgSDdGscsZLT35PAO/PmNiMgmtNoITMJYn0sq1aZYx2alY1BZtKyCT0OCnD0qdDWD6UZXTdhN
5EOZ6lMZokfwS6+q3j2KEkfDKeWLwY+iXeoNGy1ooWEMQyjtzTjL9HzXlvXKrGv2lJ+JTU3b+nvO
PN/X6WQfVYgmSR3ueTapGRRi+UsSrI4qj+AZnKDRqfl2WAeJy5Z+STC1wbYR3et3keKVp4ROYMsT
m/hWXicvY0RueUdOoN8uYQspgJpSp5kxu4HJ65s3UjjREeTCMewCE3tAr/07mvjirMR7y8jUbU5w
MF16qseZ2mK3arovwHvktu/Ho05vUCJBKX04RzTZZAdCmXGia2eW1y7pidDJI4gXr/88fg7UcCDm
jOqAmSKKpoFQc5H41tNXeq98FVOOCqL448NyewcQWm5eAAJfbGx/wbpcTA87a1dih3xwdhbdyorQ
Hx9AS0toNM27/mGLvWZ7+mAaAz0o70PbwIS8tqBwCOUvnzSBIvEQ3sa9QhJiIDcvF3Zq1x8o10nn
tdzBjveKu74D6TsOyaaRyqjsjPOZ8iYrLVQc+gF9uokGMcis7Rny6i5hPikByJTr6Ebzq1y3TQiF
dqHBMlsenT2hOmL5gDU+KzzLP+cqygZvmoyZ3tNlHXGBgNpEc3/zwpfmnz1WLDY2XHooHU1zjKc6
7muBLw2gSDT6fu77kj/50OuMVVlRbMNWWkZjd4X1RbqxI13rdl03ImpWtuRitP3hMs4//54+ckVh
y8/ZWDx0CZCROG243QaGKy5QVojVgljjfr/Ugdan1UBpdSfJFRjKaF+lLGzQVqADoeghssaUedq5
/sXzta0WlTnLLqslu/nvK2DdMkrxjn3xl6UnhyrsqdyjOV2ERb0u9s3bbw0+H2V4HhyBKKBfe99S
Q0ikqvVQmg43a2S6f5TBx5NaOZtdkUGn5ytCuxVVrd9G7tcc6IPeXaSbbKt02LYTaktHXTxuwIKB
VBZUdor6YNDeFBTNww3UThsIb66R1mR3AqDj/4DXTQIhHvDHrFhlNth9VE0QcohV5VOg8LaxnZG3
RCmQ3S81nGLYhBa61DF/gBzU760CymLYqpqHeAbVyv9XP6XjN64ysIRTc3fF7G3P/pE0zjgpzbD/
bc3c2MnOXdilcImiXkSLrW9PxTzYQ33NuqexpMRbUPeNS9tgZu0Ma21SOooPrVtVDC7KP8v9llMg
sOWG6SGt3HudcITfxzH+RuQjubP0toPlfMkmULZ/mQrmqdvoZnIiRnyNvDmYsWIIlLAYTulZBY7y
yqx4xv6ukzWQxzQ7ttGHswTwjnMONW9WGYbMytaJFpfEMV4o0pQZo3CHCrXzlVpFg8Fh1DZ597bB
SnoEwA3tOZmCVdUE/MpOkNfWRlU17DARPtvk9aETw4LBi+VlNHf5UHqR6bgP6qm03j2ygTX2msmC
Iyf+No464c6L/Uvgz75QAwn28qtVq0fbAWGduoAnInV2F8P6veKlks7/b3omPOxsxaJ1aWD2aUhG
8J1e7gK6YpmaEL83GZ/0pHrLHR1Kk79bRrvZB9wh3PpJpjd9aAfSkiCyIDI5ERDpsH6PqsiXmeSt
M3c/OCwtoigR50fT1qxo47F+0ZW1w41lu9kUlsMkc23kn6LlT0fZiLL+kpvlXq8ryHDmszooME07
F1VJZtvY/15tsKOfLiaKeiqucCD+mSf9TU+DTDfCkkp1vgEl05o4yV8ZpKeuTh838/4wpLhDwAw0
OAzmfZofephiJZh7MeAVbKdRc4jQnmYjJoUGalfAqU6tCyU0Deq8Guli4zlVU/lyiiQUXJF3pxJ5
54BkV3dRQiTFofJYVWXM0FBETeLH/idSvi4dGRTf9XDKm2Q+ivdl2h51Gnf/5bGyr8Myg4rNylW/
hXAJKtwyQRxdcCOmfB0lTnHRMUvdViidAROkEekr+ccTmYncbiO/MfixPP3jM0ZcUSyPQHesUUzB
82jS1HfJXOtdhUBzyOt2u2XJyt95XMHRR+XDH97gUZv0AoZVr1xkLDNLU/2Tjfjd+sZFwuLWYmSd
dwJiAe+dO2SE5ER6W/2cys5hIV8c9v+KrCZ59Nzx/BlO4DDeRrAAu0GTFdJdwK6Iw7JL99zv8TiQ
AcEWKxVS4/CJJwD+qlHd7dznGWZ9B2ZEySpoYZfdroEWHRLFAbo/DK1hugmdK7wYlqQKlf/AHtlx
ddABqHivpi8Ic8fb6h8LBvu0/JF+ox9RrKd4llqD+5MlqZ8ObLW+tVc+bT5E7NUekE7sIj2VaCkF
9p+E+R7x9VFofsnJVKvQNH3spgPmpf8AZgk1IfqoZ0ZeTWP7OVhWS9fqBKByd/ACBOhj7Kih7eyS
nUonnamqlqsmnZs2pu43B9K6CkAfOkcgahgTzRwcV1Udl4LfOmegGsi82YA/40f+3zhHiiOXsC3O
hTV604oz0++t+8fQrFG3/GsEbGmPoWIJoHgfWp3JhVQx/zKb7hH3HAQk4g4BDYaSnn+XpUNx6tJq
izQVaAmhEmyFPMwkUHwep6N3PAxdWaLg+MvItLiEt5HfnF59aaTgn6CJvPEp/uAA2xKmcG0pVdkI
NeEDhwpTG9F9TMo8EI6U+unacqLVnYlOMcXCOHOi+RQQ9Y6D9IvIAmEB48uyHtueDP9GiGTr54Zm
EK9HPPJIF+LXxfSrYMOOVuMTmyh7Cae2O9pDMHO+AxHmQpDuoMMX93kwqDtGlOrZVewRzOEjxxAH
EQs4i5F+gyb+vQGXR2yIAYXaAIizjHtsxwoFVevDbSl+FnJfj4zt4j6bdJwQNXog+iIdg0S0jc23
ReF/9WS+jUDkkjOGlrBTxCg4AKFxZcgizb9Zwe4WijK7ddPK/w8W8gJHUZk7JF3NwdvMr2bqRjF1
cyiTcPyaMS3+5n/NEOgG88hyZSL4MGqLeQ0mhRfyk7u5XhgQl2DbBRo52ltM4cAa5/iUYfsES1Ts
SAp0wCl5MM2MTz1u+twbLEKth4G/eeUt9kYqm/TOE6ZZmE7/vvEMkEULdaNhVe6CCp2vuOvR8Sko
OltG7kvSm6bzU2NBh7dw4B7Z+T7EfIDexS73bpvuklSue2PeNESzWHxu66w63UBq7bol2jFmpAiv
NfVF64V37EGhBFL0f5ehMV03Moxk6qs32bdwR3S6hOHbZZLhPc7nj4ZpWDXAFmC6tplj2VNSBJSC
YrI9wF3OpkUVNUIsy0IjK6WpT/wN7Z1BFmSEybjM18HBxg4WMFeMfAc7EZkntmSEN7u991OA0s7l
MErIV4XaUaL0PbvsCy8uuIpUO+P8KqNzqiiVvwwicvmL2U/4+7M5NheZkD1YQhdDv2i8gKkd7zIM
wV+UZKMOcflPE7foEIUoAp59gpxacdk5zDFn11slDJiiLPWxiB0YhIUSCqQLAia5IBHh/IWyBo7f
MtdzMlHxxSJJqrEt7U77sg7QbFVWFht9TRxOYTO5jvHgzLgG/dlNNaBeZ/4soR6Tc2Iwx42mx2Ik
VH+ervtkXEBO0rYPLvt7Gow5WhQAkPhrHhlqryrB/UjOluoaV6YHdTG+aS/CmwiX5TQML58suN9V
y9sEmf9gd80/0xQX4JytG1+rrnHU1PyyhBzwqoISLqXzjkSbp32/tDptCQ6kfMfP9Z75qq4Y9GhF
vWFEr40VhPXkfdWzqOfkuvLW/4++jSFe6pkGOfFyq9HygqDfpqSc9cJS9TcuJRiYwXftj/YrIHP6
e+gECW2nWSLqixNxTaRZmjmcy7s7fuT/eKiiDB6fZgfUcEU0qH6VkUi4STYMCo9cOUyEHOypYzWx
pCQsdDlSFE7OqFjJ5/XmY2rDUlMG/2uxyOsc3CqQNy5oVHvHP7odPDPbIWdu/V91cOy9EYBz04KP
xHkK9u/1ijP3i4WsL/XTokhE9gKauUEFB36tHL8e8ECq7tk2y8Ar+a/4W23GPtQ87zzei0VeXbrM
XvEujuxZgcgn0a7b5QQy7HRNs1vZ/AVjKrMjHU13tV+pQ3VZSVcdvoL2VBhuLWQiTSQRdYy8DFQm
rp01I4J5et5bU8ZKmBWog2PNHeJ9u5BGUjEOHCuJcoIWIxqJ4oZZOigg/V9ZqnxCLUGAgz6Pc7CN
uBQyVvQsBYhJGnHSZgvi3nLxw0ss69gKIiMV/PIE3oD0S8sOYs043fxqiJjivJNSbgVMbMEypIIC
hLWVJOcaruVH8w46ZNCV5rN835cyeNhSh3ymwIEsNsetpqrfrjQM8PN/T6C0h/1VkOM+pTzwB39L
qE3WURSLpy/vDZ1xglskE9VedELRkvkUkWcWlfHhJ4spDgzud/n93hOCq2T/h3eFczZT9AhHZl/g
GFVe2DpRdCyv/OSQH1PkDoGp96nB7VkN4gPR6MZAGnkKHW9JgbVCtqAEUEhSHKVqMFgNxcYfVjQm
Jkq8T9qMpZbiIPTqmBrF5x2BlIyuI1k+y7yce6zT0Tf7tsFpwVajtRfyxgg2d9VK7CaZRkeOk12q
iXjPJ24aRkksbt6ndhe7GFSnXEtgKn0M3u88USKK7IOQVLlYeQzMAzyaTUwTBEXCeP7fPnyFloe+
pcTvj+simj22zsx+jdLi3zXYHNCvVC/iRR3DAoFITxLZ2eszEpR1xHPq3TmFv0jd7r+22kX56cqe
LlF55J5AwLH8u6j0BRYlzKb4OGPYjCCHrYheOdmgz4YwrluSwCMa2leNYJp8HPhb8a4f6s5SIWdK
KFxdAMMD7I/EZyWQRnZ5CBomuL+YzBb8rZWss3sOWRrMC8VorInHa5zUblRTHdbul6bQBcx45Cht
hvKSdSBwod/TjZ2Wc1rEBEfwejJ+BD5ZnQ1RV9vQNprYHZpsjAsOSHWaPVJBm17igbhYZniT3mnJ
kf3Z9S1hVLieUMmuZCKn0kZ3xzO+Vm0XQaRrUcgeACt90pIN4t9ZTy5R2FY3abIbubJ8DdY1Fimq
YSAFNwe+Uh0hLzAfhQuGG/qDA7KjNpgFhJZB6zkMzaqX7+KXiCBlkh4vgOvfs8dAFQFmovKq7Jhv
jnTlQVZ+3NhbaZB/K5l0f5/3yEJdvWOmG6SycwXKBFrM0kTrUnCeQnRkV/dGS8OI5si6R728MBv2
g4QtLjlVSSD6XMapCHnCVHduVjcX1ClAVffWOm568bYtYwf/WfNoPCcdQ1cTnH4Ql3eJv6C0X5OP
XOBIPnRXGegyns9U6Ph7stTbdVvWMQ2jOHfDiNWzCxb0hHyeimBV1Gi1kJI7Wabb4im4s/rptFDA
I4HMKLqgLjYlp2zPak9h9WkcU/rJXzreyX4EI5/7JxP/9oTetBHyGolHoqsWjDE5lyrSMyMhRio6
ERdwrFnhUye/JelPMyw/z5hAGcL8BQXQdRqZwmaj2KuzsKKno6JSU8HKI4FhKUcmNyxePDE5ynf9
1/nMwq1vSk7v0lHWihOjKTlRLToehYdK8kpm40/4s97ayWYsmOPIGYglOtNhZRk0JrQwGeAAnC+4
dWTVq6KIfOgzDBVxCgRvLVIPlQRBjT7cc4YPwMA4z09a2cnlCd5SxO+WyeNUKVQDa5sQqzmdH0ww
LzrD42rgzLQmmOzZdvlekGcONAKZ3c2cvYdjpbAvtJhmjGdpOGeN3MqIFR6VcVQXv0MwzO/QjF8e
tNWLLIKZIw8kP6vwGurMjdugA7Zw3HQ0x+VGqeAr0H0i/9RUImltwpBwRhKoYMN6jGB7dS9YtbYy
UJBPlkcy4WA1/eHwT05ZE8no/rXE9JgvrRuxmW+/+B3wAO5ARDPV+TKoZMeszKqjKFnLTMyq2Sgp
gvz+T1jEUNnClEGVOMHg/gN4f2dl3+A2a2RjipCa7RqmNPNlzbQF4M1Glt4YXNZ+fdyt+UMgzWQv
yUMhZJzjKcf1q9zI6/QGUz2h4CQTJXB4CqUWybVY/TnSvLqN6sciI8YjmUwo3CMktmzjHaZUZ00X
Ge7J2M4jhAnLkbHBlMWYIm7XgV5qPwWFZL5xAGvLmxYq7ywnk/4qTJbdIjNKae6inVPWolkOdU1y
/xL3R7ULAKzEVjsZhUzxUgtqsyL+VXJDRUpv/K/aQj6X9FoIB2QrO9Pym7kRTSjYirSBj4YuNVSz
mBzaYPIEIwfz4MKP0/uQ+1pRY+NAXp1GNqGj5z6ZIPV+DdfFKuh0t0lw1Hhrv/VrN+hgjQ1Rm4dt
8UMNb7LDx8LZyKpTblQj9c3LduTiwXekzZ2/qM/E3H3yFZagiDV+X8T3yvrGIHPSR2UMPFkrgmpU
txTYi8vQ/NQ2SWd/b/+L+HvYwSxe682IetdokPmJllQvRPtGgWZ5j3QX3BRtEZ/oK8/BbLagm3qL
RX/+gPe9p82EiKi+qTu74quPrprF2IGbKt+LOQrhykfsvv4bIOzA9zY6NLYwAvBjwzgXNK2fspe+
0JzT9frtKitGLsvI9MqWbQj7mRTTRD1y++g0+kQSmNAMTMNj+gy8pU+4BAQVg8QcMDqbIVqiVtKb
b3up1h5x8I5EcD8Lkw63TdoY++yEHlVVSMOHtfWWSndK74nJqND536gk87JJjpmOIvtdTmyxad1t
ep3AEAt69TRd/HPwzSaZaJKxZlNE7I+TCkKAh2xNa6YTphuQn+nOUVO6mZtofC7YvJm+IqoJksOr
cnvIFXYzGKBzoDYgMjiXhCDY8yWJMRaUyt8tmsW+f76Q1PuBeug64uOYmgIKOAiG0LeM/Pt9aYhN
/6uzfpvpgXscEcU3f//WAVrIqbuZFFaloaxIeCAnGUYCfFgeXtYwX3TX8fh+hyHcARyiHCTKn5wF
wL/aujJRBG9qonk7Efa4Uly4MIjuDdUpi5Me8h+zCR6pIjAzMkIfffVLmbsiYi7ihEBxnD8PjUOd
ftHd0v1j559XyHBxqiYvdHzjNpX+JZE4fHdd4Norb/0EnIXCqT9/UM+KYXv7LXbBjgGjaN/3I3Xi
nihgcscMlGj3ODunQgUQKkUyx5Kakv239BpfMWzlERBJ4KGbYdFX2xB+9Li9SDOXzcKmfm3KQynr
S7gqYgZS4TBLKLNlDd1CicnxtKfNX7ghHcJiLG0oG8aeqfmRdHonlvvmERlfoH6aeaD2g4EXKGFS
5qmCxncQq3z1jXYCm/RIzlZPYMsqAi9O18qJBp4I4NyfsOZAvUuUFlxrZHUrn+k5aCbbizWy2k5l
qnQLhEmFyjDLELe8Rpn5Exy4bmRpp3fIawXZuO36OEwll1PHVhwE8bHoyOCNgcEcvfocPzVUUkSM
vWTB9wcgI8YNLcrHEM/0VXx5AEej2UZAZAScp48of0MlLp/oAdCw8dTjaMT8/o3Xq3tKBhYcizn/
UqBjxmv//yEJh0GHhFEjHkD0fhee44mEBXkppiqspg5ErH6cHTKgXkhuhLcc0NOvm617fCHbFKc+
aqldU5RIF04TqRISpH8D6Yq1W9zsyoOdDkaLEc/OxacUV3Zt1MPpKKb7x6PIGpHHsuXeCw5m3wjW
t7p3S+wSrHBJlScbJTJ0FbxAKjOKqq+M4+2nVu5FgJ+6193b130aaURLXeoptHH/jSW0B4oUuP4n
1kRLsKFg4/zaDp9rYu/iGGOLycPnNDeQ1aOdcIHfSDnKr74GImi7gymlOWpjoBaFTCz/375WJnvl
XeuV4C8XOfU0W+6aHEr4GAfMa6YbWzmwqEs11eN0XyJc6oBbL5V31Tnps9OIAJtHwF+VjGOxqroS
jTUFfmMd9uJxXMBagw9osvgsjTSU2uZgTOGm/gX6v0D8DPl1AKpt18MFeEPtwjGWnZI5Du4EUDBv
ivsEQd7pEldMFALaijHRNjHpiZjwagFwf1RkHXx5ArhjI+iFHo6lvJdK+iRbmjCqr+u0K3Yfsq6d
PwsKchhmIQDaqojxJswjGST30BDdj+rqta/G14WKdgViXvRbleVS6nGYAru+b7uboRw9r5uEcywj
lME8ahirwCXoJkWYeZ169HS6gxmjmk3P1vF1B2nvnlRSb+rQQWyeP1PBDSQLeXk14lFOkO7bIPow
oRHW6wWZnrrdX7ivNOtgqxo7ps1q+DprWjbOitnMF5AHn5TCMhF+gfwsRp29D99m/zQAAAq24Bam
Ltii8/LBMr2k2/tP4+v362wvb+UH4xzW9rhMqitYhdv1sjRm7U7IOr5rY6iwnIhykfUcucylxHcC
p9oUqyKtFkGf7lWSTAvdA2C9yGPWnJu9IoaHah3ozHcPT3hJnr0ImGwA6xHDBKDYPJevRUGNmFEc
BhegCNdUn1WM34hP2BLRoE8sPzgGHgUGpMTN/NRj1H/DNuQCfTus0JBNJXByNkJHL1SSE3xyMI7W
dTBYhySrk2qa65KoCcsf0Y2uLjZhi3jRVimDLxFCGXADPm7im/uSXglJR0EuEHHR6bex0NSKpVm6
T8EIsNZDle8My/JO0iCFK862Jy8TM5J1oFoFB7faYUi0SFPZC5/xFXfVZO1dRE+WNop2273eN5cW
57Sh7efBic9y6o47xu1zzQsP1PyT7g0SQjaJv6sJJvHC7Ux7MaBNAxamNfQWdwp0sEJQFK8FOWYj
3pQZ8v2jxpkWlVTCv4h6GUarJhDNertrMNosrkPvDouGWj/+6t//2FgoCaR86ZsvHhNpZEmBgT/W
x2+ZkN2Gu3W1/vSzQ8xYpXIRdWC5Ng8EDGEAT3sFtVQzWDYY7V+zZBN3aYsQORfRrJX0oLsp302B
YdNEAD2YHCOOVGqSXxHamj6NOEirwiER4bYKKktCtV8vHdWjF0A0LelsbZO3Ai4D/QSzz30Ec4Zw
fa+umwITV9qt1If6B2/OQfQykLBxBnJjF+fF7kwicHO5FxWvtydKyQ/fD+UakiSGbipppuO4A++a
DucIyyiP0z7yDI2jCrucC5p8dHCCJ8MRBEqqOazkGUk2tEK6g8t0NCZeSEckg/vQIn2VL9AKIqs6
YVSNTndhQcQfmKCTyqPyN4f4e/v6IZblKpDrr9IOeWhTklu4OlFXaOxLU/ofY2BZfFbQnyPyBl4v
SI+DWi7H3Qt0mKhsP51/7M0MSj12HAGl2FU5m88R3ZKASmxlHOfLoOEGgd4bMb0VTYAJ6c7+IKC2
zxEpcQTDVfRzh2z6k7nqv/haN0K5w1bkdOnna+tAv0amZL5Xx3eFkBhk0OaHPKE0ciuvu/LOShLg
J4l1AZvRMjrbDyGrGUAJagiHwbknOJs1PFWax0VRFNPLbdRMv6e/rCYh4x+OrFzQH1ofsVSKInOQ
5eGD800bjHuotNdfGD0xGpjcqFyZjb0KFI9cvId7O1fwPy4TLZOrUGUALmfeWRVOyiY4hzFJtUyV
qH3vy5s828pm0ImrrItcfY1Ggg5mrsfODeJt7MZ2USPET6sWFzVabx9UOY35rmkWoT5qy3DpZRPl
jWZLBilyEOgiHwd6kZVW/ifkDHEj7vlTfWtSvPmfOG7s9l518tDRZ9HZdl4Pg1/2EHR6/OoYT3hc
A2v/Nz+UOIOwXhrtUvwuyx8vzaojm2HPJtD6lGb8qG9A8VkSwsgaa0ll8ZyIlQzeS9qokMNu5mcP
EdTWmgfNrLgZt5GjtHmoLhjrWfksRIPce+XnavqOVbJh+6XvJNkkakzGkv2G+MqazNC9dHNYI7GG
Hv6lb6Ox+teeBtTy6CapZMly6aMUyuxyitbbztBpYOjYj0YLS67n71TV36G25IiD8khHC/ud3rMf
4FYIWDYoymZEqZku0g4OsrzgiTUviDavwaZxl2UGOusJDJJnFXky0YYZYdVoafXwL4wdxBRxDdBS
CUiZ3DJ7bAHTl4pPBeZoKlYDf7opXiTIpDyHuv1OsBeQBmZ3q/u8UXMWg7mXFcsYsBBSyb0HjMhY
EbyBWpVv0qGxH/X6tKNtXXizOtxbq9OMAm2Jxg0d70rQmVeOBH/Ykp39LIiZKo+kyyZlYMtUVxiW
Kyiuc3YjR2O7zx1JK/XjriaUVxduDSFBcRUHHGjjz8D5KXIP+/fDdQV6aePaGSShcDyThMBqOwlm
ek6FpxO0e1rB8ddAt6llvneIowKq6Wj69PAv9dShbXnzxgJINsm0JfwmsdomVH7+R9yAGeADd5VP
IgEw5qNZfbW0B7kBh3/ZLTNdRFJLKR71ur4/dxSPi/waKscfN46FGa3o8lzTCRnaYS1CY8A/9gb0
Vw0zIkPN/Bpki5Vt1m7CmQUodw2iKmXchvevO2QYNj22LAOMgu4n4tnwW3zjn7ga7LJOb/7JQih1
C19Tbo8z5z/cBUEHKROUAHx3eQ6W7Q0PAxaEz7S1MkyyvJRN4f40Dgs/Vt1uF2hEx6/jbRwAfWb7
WC3bs+0fq/uvi3MYz8YJMp4OpLnfvqGvzt02pKXAEYP/ulFETojBJEuJ+tSRPvexBGbMuRCid3jw
rxHin/9eNv+aFA/QpBzMSMZfI+yxuNdOemuWQR88w5dY57Lwwl16Gw7XtmX0KKzw1rKyuP27y2qQ
nDW8V+NMZDVSZK6zX354NbZ5bnPJQc7lYIwNTf6IlyIlh9pPPNgsdaDIAZwKhbqwgNrum0WTu037
K0QyXEYHnfDai1StaDNmypE+J2+YP+LrIijUx3fanxth2TekCCny/z/ULqCDUEZJ3N58SdnQHYc0
8G2Ocxl3DjHa58MawjggsxL5x0VFrYvfcvZJo+sS4jgGMtF3LYwPQIeEZJJ6zBJhX5C7P+qyLvQM
GzxzfiqLVEYb5JZG2DGFTCz0YW6+4Y4/TbgNJji5Hdhr2E6RywRlqTwCmAQCtqBXcHXYK7ceWSAG
YdxEJDDDR/r+gxI7Uay64LZZKuoMaKlUakh+aVXJa09xlYxQHKQZtuoGBwcMM2Qj6Z2hx6Sybrbf
lH+6K/tb0qshEeXe1qXsTuSjRF2BenZKvpoRdPmcEv/sVA6oQOGfSv1MGGM+nCuFHiWgL6KBo4NF
w/zAIGBnrsFo+uToDQTrEmNOzLSUaAFHNGnQ0BLD44npo6QSw0pBbot3SCi11U1uYSfT7zWcL3hs
phB5ZUM8N6Size+fsP8PLW8iM+ddP+xs0CqHjL70QCnOO34PqFbvJ6Sob8xz/RLJ1JYzrL0wrHbg
hVZCrx1TVxyFhRUI31YTBYp2BRXAk5O1RHgVyhKLoaF8VWaG70QcSq6He0Wq6ifd4QvWrcoypYln
cfvjDvaBN0pLcWr/IpGDgiHSOwPAByxHu2+8cGmY9LVc8m/i5JrtNtfY4vo06cqjoCC0V5whSBKl
4WI99vAsnGW0yqurGvZQgfDJfz/88DgbU1I/6HpRcF92mDrYM0bhPnqxlsiXdtMVCLQz09vqa7Mu
SLPWGe/R5le/RVpfjzAKVG1mALIfZve0eOuvfT/9pRMvqwnFV1X2GNQjljmKsgyPlf7wGiETmKeU
ZMB5dZKYqgUEyaNCuZkgJGZwvtviIyLuSgahiyf6ifNX5QEcd1KXRAO+H3WBYazlwaEc7+h4+N5a
qGqs3bFfbnG9ibNrjX/J3SKHXrdTRaFdAPvVKQWTIBXBxmsszkHiYm1oyTnfBTRBDuIiRKXlvjGN
h/J0k6lbDNGFyf4JBxeDMmOSNSZ5OA5Y7GBwb6zKLZBCpSCy20J2wPxPhjSUE5XQbAEsmIyWAFwB
RzjU/0BtWc0OHgLAhHlzWBl2/Hz15wdYTBp07WyL1/LqFENw0IgIUqcKbkAQO1lUpBjcYrjjT11p
YLqsEAY30lqLlKxdAMYue1FyYYT+jsUGoVHyStjbK3Wkq96yjkWnwox+T7xmzp/FDtSKIsb71zEA
v56tphSpEvc5yY5K+m2lnNuwKFh0ZGVbYN6nrPXtRLlpj6+QtPdzBaJNDLQsy9nSnY8xkC1FhVIm
y0WEiocA/azaRhNP2c4mKm1sTeDYSmTf9JkTJqsq+7pEIi0Fc9MUEm69naoxva7Kc0KQPlDN7iAi
BmgPRLadX6eOtYA4OKh/AKkSGkBesC/oeg7eD2ljusDknjcPO1No2/YCu2rf8czox9aPHz5JIvi4
ZKYWc3oTlrsVQHNPK761WpfEHD9LoWlpSaw3JQ4EfNBHiNwrLQFa6yq9Fj7tUqa8mhWxujrEVR1F
zQhlt9nlyh2+ruKTlv/c5AUAtkjqum8fhnoDYm15a0uoLODBcTU06Wol13Q+qeBDyQ6GI24UAfnw
OT/77s8a8gOXyR7jS0nZPq6RoLkY3M6ZYVE3y29zYIjxFSYun8sYGXCL3xecxu5FO66bxzc/ggp/
o3Anpk/vyld7hIDBhfaemC7YlUzUY5IU4CeGg45HLtBv2OqKdz/86jZzgTITnNd1WFRw03baRRSX
BKUStU5j+DmNHT6PBvjluVzo42F54sSon+R4Cn/EJ52h3Ak+F3J9b/pYdPutMM4XXGqW6VTqH4u2
F/1/rpklcRRpf7cuaFvpCkMm/ggGkda5g/EH7DLiaARcfoqiv6VK2GaZFkKtaZzFgy5UwTxdzL5z
oUECVsaWmbkxBTzDSEyUA3HxIS3M/ULD/7htOfd91cgk0n04mN1731NQAfhPo5lm9Gf3PEX6d8xb
ml2uGvhgVBBRYsU5GO9cVIdUA1PEtKzBsHcn3tLLYQMI0IU6zcGZjNYAZ+LGQLnjSSUvZcuxnnDQ
xcyQDsEXxG/zCI0FSI2rEpnYxqPXQvxFYK4wh5W7wee+hNatTXvXJN2JXLl8HmAPHP2bYz5hlVAp
bMzxcbnaFTJLrz5jctIvtVzW4oGGh2Bsx17WDg6r5RvDbxfoOmAXCjOv/sVwoMMl5DxpRnZ9ICKt
QlztNki0LSYRflJzS5CZqIJ5Hybpg+n7XG1T5oL10FhQWrMAgitU5sjlA1edLSwgxSZw+t5dq9ED
rGMJ8MFN4bwiSlUEE4MzKv42u2utzS8+Pt0JUub9AlqRSTt1rtAAUskYeKndwRexP1Sj4SpG9a/I
ZSTNXOsFtNHHoT9xMiBxeJJXYVQDNjs146FCg/+DjrzHmK/Jr9TJfjkFb4IK5mk9mxlrNCuNl/Un
BOScLt/KMk4pEXV7SxulT1M91i3hetv7dtWCUAS10EAxpCGR1K6h+qa4q17xLF7tloLpSViScYzz
LMH9f3pZkdt3h3z+VFtlw+WcBAwxwsSGp4nJ86ltF4FF4DCqBYLhOem6L2cX8So1MUlg8gfDkpZw
c0F1M81U67IZfYf5ic6qSZ6StbsUPnRcKzFuRqcuTqCfZppZ5JmfoWkkIBx/ezGA9ubcQacOW0k7
0LbvDYJpCq+z2NekGcQHbpvo7vkN+NWaG9CuPBKT2mHDJKSZm5vcsG0WPznQn18OYOOTekACXvQb
Ggm1kDXvn0/c1nw7hXzYDsh0k1QcoPqaBERbnAwHKVM60xL7iXeHxMwABYAFChNJ0a7dDcF0/E3s
ol+2Nnl0sAFXiLARvuMI9xY8oyVWtgp2aNp6r3E0cpwnfCEa/sq7HmALpdXGhc3agyA6SvbFBc5Z
5DqHx44HL3OppNkkwSSfMqtJlYWkX58O3dpRSVdto3YdZdgmlxM1jrvHk0F1vvEI+fo5JlsABWLM
Luu3740gCveJi6FuFXxuNSzPJVYs7q04yO2juoKt9jAOyciWQzlZjnChsDeW3qMreT60Z4VFR7x/
kufB8+/N7f9mh15gmP3++z886oibjzrFny8tGndk2KjTIyl7DUIdZ3bqmYCBg6QHxuKv7D/yqJ0h
hOURcYG+8kI3loONlQppNv6JvaPLOTOClBdgczj9i9JM6GGBpVrKDGQVscvpG97H+v/k/eDHw8uA
T623FRd8R2gmFaKEFWg9T1CDAuwx+yynwXH7ywFhhWcxGlm9PgpHybZ5E5nm5mrjvHvG/ZVtAONR
ehlxh0n5cwg5MEBcKdufdXcUIql088BZaOTklNQYiQIzI0FkJTcJyeNaAplK0OfobcWQ3rEd3FiB
zERx0Ij1oViCz0JohHKwjZRQrS6u96GtW+zvlkIcTGCwb9mhFkeP5I8l7H9BXFL3jzbpDyzJYBWP
kWfrBxe/a3NkuBfsiboxxwKwGpEqQ+UdW5tLqESVJhbHw7DmS0pJIYry6p4/ZAuENIJTSVaiqifH
7U7P4anadK4hykHezEneUi/t7G5skYuCp1D/mvBeY8Y9fHPhSpXnA33ZdRyP9vi7VN6xJjE0Im4g
bPLoB35p/fOSKNBYhxEFWeri7OB8ma64dKIri/119sm1YT1Uk+mnG1fARoEgl8LLkg4EOJ65pwkF
d3IAFkR6I3GBEJhvbEm7CgnoMh6w2zp1xGljxj7sfD8/seHMuy1yiPv58qmTwaIiJRSdRdvTXMDx
xhRNeaeGLHxrU1aG/IBhDhr3U+Xydc99GhD6SJ24jeLTV9BT8ppG4ZqkutRdm6w7n7QgejaUIU68
FGi9wEiWsLIzmx/a+s2qKVZ4Ys3sdEgeqN/omJpfsWDHaTxuAXRQK6ODeeoF/xIIG+73V5akZ2x0
18tQr4jIlwaraarRUIG9IXdlhd6bnatAhts8yrifd1ssAbtvqQixCSC3ovoQ5eaCXPiYtFyVbufN
J2RnHtAknY1LmhwyWb8vrEJTB2cP67f5/1s4Iebb8CQ/fI0ZKnWQEFvlMlllHGIj4mE3WWIRRkZa
Z9SALaBDXFBc0vahdnDpxzvBXY+x8rykoRAbZAc7tqAHXWIceHraIOwlmPRvhRirln1G3P8IQZdb
Bsv4XRypV7gtEf8xdWPzMyb8w2ZvIA88n8gcYXQCwjHRUfZMzVpfyvhDsGHKnptAioSFZ0sRQdoe
I9p0jSG2vqp1B8OmSfqw36wUz8PyMX9qK0/t0kdQzQ6hOF94pBjDdneyH/G1rgli47DIlbtgjJic
NAdFsXiGqwNpzToyHMiMur7EecVJNBfhxz6tqOfqz1Oe1+RnNCIgT0HaRQZxT4wH0oieazMTgPiG
rc1lCdJD2GmwGIPORRfB2URaLiavjLlm7ZMH8K03Mo+yxrwb179BaGc040c300c4GcTm5He+vQ8M
y8zoMqcSn4n7McMEweySao1jeNfx4+yuOixd5iZ+V/wD1peHUMTcqOCrT7kCDySrtt+wXxK00kE4
QwYMzz0vAwIiNICEtexMCWSBBl3JYlz6HSnIFdpH5tgU+uvTQjOD3Jnq0FZuyxgqU9jGRbx3bnHo
1CTA4dKHM3vjztNQ6o8eZFYK4rz6ofh4wVlsKB62eT4p2LwYPzyBvQBYfovR/uUqCLNfdFoR+ug0
1Ubo0SXFzSEFv6dOQzfft1OSqmzUxM4GucjFiS50eWgHDwfuDHcKjMv+LI6JZtT5DGmhuU29AnNB
x/qlnsETvvVmLh8BhreM4BSzWqJEhqLxvMKvSR4UvIne8oGPeREKNkxwLU+jshVvzbe3z/Q4TmFj
8W7QCTP0IWgBifd+eZT9NcfVzszTUfi6T596C0h4k0X8I/E0wfZJvtsNPmpvxzEs9QYOF/bU86Eh
twxyKh6V/UEeZw9u3bXkAN4tUJU89WvbpD309bR7AcqhkK/0VpSM867oMCjdMBOsKbrkXkaOqmiu
WXmn4nMPIWOEeIeRORl3dKnipdwJB7c9KKOzrGhleyNaxboBIqizQzmfs7YXebFVZ+qyALExr7Mu
fWHu8GbIUJb5CqSwpEEn89dpe4SRlmQVV7fth94moG1bdhVq2WpR6NVf0HgLVSyfgl8lePQie/qE
p5/nVbrnmpJjMj3yINrRONONhPlLLlRxbg9azvqZLy/ElbIbty62CdUyFdmwkMkRBlwQI6RbU0hC
w/Fb0gAeYOcgWoJuDE4UetpV8httCZNI4d9tEu2MCWQ96+DZLt42SNzccc35d2JSIdnNgqpSWGTN
q/iZbs8yG/xeJT/AhT6yKeEB19MdaS9UzNY788+gC8aEu7RL63p3fv+7dIBFKaboWqgaPlURC4IV
lmdMbd0H+/ug1EYp+BQz0wZ0J8dPVq8+Jo3EKujgNzDe2WE/JvxxqMhKjfNEm3eO5npFb0kHmfNQ
slhonYoncrFzS5xONSqq4RK66FwtRhTFV0UYgU+Mk+W6XcpyLT1S6gXMAlQ9k7rFpPKWf2bcO6II
p+KIkmerPdX1CckDXX44QHb06iw2KwDGKMrB6OYQnoxabgJFzt15b60EVQehSOvkQzDVqWzVLeYb
CNoLaUXU5WZQZsDF9m5GsvHFAMotKToWw7N+nJavPeVJavBnFJRz9mmnmp+wkuFQEnRlC+9jFspU
OAHcP30H3UzRzp9kLtTCswQF9h/xmh8JlM2Olv7S4zueiPGUR0wjqMYQV/94fSRR7Ih3x7gJwTmv
2a+2tx8+s6I/s8iTvU/XmiH8kQTLY/RzUNJvvG/5d8Bw+Z63zzKm9ynfXRP8nVbK21Rubs7qi0m4
wXNvM0SOX5DE2tZLUK4rIZv2U7qTL0FjNz16N2P9StMnzsd7uim4yjEObq872GJroPZdat1pw7mS
K1H94Yuvdu7UqbGvVmDYvx/TnuywfF0vHkJXVG7cpxKae2kKBkX28dTxs9r3U0Nqx9GYQPI+5Oyy
6ue1BrEtl4XeImoK1zMjJD6K4YkiESOo8IlRnXwCjZwD1lLMUAtdGJrLrFALR698PD3tAMm3ZBJP
C9DqiJisGREcMIDVIuRhDvdETYhE8vA0x/D7a54kMZCdHvg6FIzdhfTx0c1ng9pi+QrOlUjvHwln
1TeYsRrOr3eiiqiVk5R07JqmsBK6VIbqG35/OhY+n/grJ1bEgRWV3LL7HXoKJVFlJwh8xBzM68Jl
yEwY4BHq0qllM3bILSR2Utdo9quqx4iwk10u0J+GgwosYQHBg1dmAF4NPpSe308ObyNNfNUfvQ+Z
tgn06H3mAgz2aySj+5g5Z0vdnrVrb4/q8E/y21GVAlFogBihh3inRK1zA9dtFFTrPRms9BoOHDrJ
DT6BexUSlyccEzsxwL2lHZPUuzEaCMANojTjvzs/Bqt2Oi3E6uncFpp4vlSjInSVvXqHhMDhnVV7
kdt83sDU5ATZuvu/inxLTqo4hr1bYcVmollQa8jYVBTtxb+LqFiE6OcMmoHf/szvWC42m/3Emry1
GTXylG0x5WOV+LiC2dz1e9tC8d/cxPPTku7yUIrSZvPEmlB+pb/n4MVhebATUF9xJq9kcyCh9gi0
C+rvfM8QLnG64O+2MbUwwgdQbAtK8+h5l/63mGHP7sDnM4T5mI7hWYXHmDLL3lqfXWXln5daBt/x
c72gTeDv98SIcoEjEigaLq0/4QFTb0QqenLjkxFp+uuNKxjIDyumzwI9clbYBZjhLf2POUo0DwHf
NrkPt0FwDm1Jw3nFzdPoIxmwexckk5kCaXKtU5NA/Em02YL47a3DWIVBT1aCX3FMzo+UOFtM9EJq
CeqXX8HbsL14cMvsfhVZaFinQojAXaXiZeFqY2RAfgSORA2DkJ/ek+1eeFl4LCAMIqQZfPv/RXDb
+V3pvb8ZcPpqAjBsKXTMsjuiHsOXLRq+89YJG3JGc7F8sQA0foYbslC4YhKwkGoPTz94Ch/rQLsh
h8cmw47z5ky0KeR6DHV2fd3wuuRrPjPBI5+P80dcHruX1f9ytvvkAB9ReQQZ9Mt6Af3rOGaURUnQ
VUaErwuTP6KzE6z3lhab7CeaFEnDKAdqVSmG7odOT3267OryhlrgoaZ2yOG5KwEymT1VyixROSGt
djaBH05NWJGwWtTAlpX6rUdmFRwgYIlMYjgIz/o6jBCUQktsvyJFy1ZrVa/zVXavGXJBDwk9Phte
c4zUW0Mx9DBNJ3e2hHv0jO+9/qPrN4ESXEcWP3Uf541i1bvkqLJdq27hI35dku+KzLIXS90buZtv
aF6IVXgBVV+lNalvO8LHJvqHGwVCIGaIhMVBTwiLqm4P+LqaurKn2LZPEFWFMsStMNqtJTrLe9o+
aWRqMYC3nNMLSv6AHmtnbBPez/pSBCAvPdYvKHmvV5y+HrZOVgh2kxWamqjJslK87BifdBqF+XxB
Vx2HPcwPKEgu6B7omSW7Zd2/ejsiuL77Lc1NCzoS1P2PSa7EPOieB3Tu/8VeHadIWa9/ClSHm87W
aQvfkgD/A/Rm3ngRqRn+VX/W5tFdKojTUqaSNLkfcIs0Q+Z/Yj/iFqotllMNG5xaS4jnfK9KwDku
TOPhP0o+Ya47LEHMfKXef1D6m1uyalLINCh5W0johtg0wZgzqeNpxHmDMXHRXmhrFX2FGf4vHHb4
64O5wQzbYxxkrMN9YKoq2iBsHbW3q9yIjQduJOVP7k4tsnzPH2L/BG+Bi5T1Ha4jLCHrR8Zi7CwK
sseN9HWVkDl9H4RWPHBLnN+Q+eH+e5pu05r7M3boRJ1ZleloAuPwM7TYwKWRPoqxlhuZha84KEck
KwrixHnocFcQ3MPBf4q3m1BPHXXFbXrLnnGQVvetUQw6ulwdXX3mYDqK/IZEV6lRx7tgptf7F8Mq
Jq0nxpoFfNUp+rkO+QHeDafz64KHZAr42f4WelZOfj2clk6TMPji9/G4XuQqBsO7jYhtmtH3q3H0
cm8Xwll4cAohp1jIW5huBs3YPAMYAT1RYzX35Quea61BmnUE6zj7/UQ0gxj/Cnu/BPgU9CA+Kabt
7VnlD6/3fkt3+9G7+ChnkGgyJepgp7M3FkFuwXVnWq2BWs8ibFCzVqRew48Q15c/9OwpGNVkGGb1
yd+aA2XbjLc/D9wyLEf8ZX7T4G9wc1lc0uIxz6CLpFqfvUgFQ79r2KIO0hTgFVYJWaAPfx4CnCIr
KWYsoP5Pd1mb7gS5FZWu/K6US99e/gJM0FZrS4RuxuLYDx5Z2nthKvTAs9ksOIsZa5f8CRKkVkLI
TKDoEs5XwkSdIXJq0MpjynsHFOufhPLyP5NMjl01cRuCsh1sRRPx1qnbzevPkQp4Iu7FSxERlaiE
zRk555ETwekXvYFyEOW2OpEU07UW0i4qdcj/nfXRBX3lteJwZ/P507pM38ozZj7/b7qNvlIuFuiZ
3HunAC8WvItn9lxAR5fDPTcXROQqXNGKRpLgchXVqUDvrDfgoL+bwkW4L9W/o89InWCex5ku7zfa
6M0Ze8QDtWMQNSPJTMVMRwrNz2qaBCZIGvB5iE4UBggsT/1MqeMltIImW1d8eGm1vmPVSb4QyVbK
Oj9EtDo/zZFNl5r4Ml+z/6PECWEsYKKfxnGh29nkWCfD96vFOd2YVz7WmE2xwcnMC8MSOVayU8nS
qnXTDHvsSGsJUZCCgWMWofPIdKiIwsWX8XKKfIH8setol+0NzIVcNRxHsN2aScWmgeAvyLepMQQu
XG/RBoNCjRz6/yZEDHVpRPPl1Skt6CXzTA0ZT2LBoaqxmjxu4E4sVPrqr7piYoQI5t1M0JD9L9tm
U+iL2kyLJNQYv3JAk8K1EUeauNHKOwSMZQfmwTXfZcRR62ozAsWKg1bJNisnNqY7ZsE4Z96lC32/
EKBSm/LSZrqw7wqLMV2KMMMmneT3AuHrK41P0rw5f4HFLryM0wjTOIpT+0duFn/2gertiNCyVJej
14DMF+Fn1vzbE2/sCNeMkwdgfWKrdXM3IFUXfB4GYnfJWoybUmS/DrWQwnwEmSvv5djFYoO2xQOt
+DwgOB0RQan7q+uDfcFzbbHgRo8aQSdEO0soJTRS6OqsaP/TqerWFOzGGaFe5+hIEvbtQnlFPm86
V2JvTgGHLfzL1U+b8jEohGzjc9mTdZiECXIMyzxXZAUrw+iBJfjHHE1423AKoHFDnfT6j20YzP9n
rpRA0r2iVW5+T1izKioNTQT2bnmrL6L8ZZi2yNvMLmdIP530QRoTimpPn0VxuDm68k++N0qH2MUP
MSAvt92n7sdhmODI9uXKrr9o1nvviTf5m5wXdR5EFX9Vxtc2ko4qJn1Hy/GKdQBFfBJue/MUsjoB
ztPLKCBIol1B4WX/O1YBep/RUS2+vgq9BGDcf5hnahhoOJCUIMIAdN6OO+yjdZHOy8y2aKnkyX2Z
SazEAmtdGiD/7g47MKNoBVmQxUz4eM21u9Y72oUHV7FzcearPprxFtqMPUP6ZQxlNwpCh9RxpOd5
iBivBpBOksY7UKmvUwROJ9lAzmooz7dUODqXp8TNHxAlr3ZaoY2SNyp2mvBljL3mbuj38NMSbKNW
lQez84+5jPZHvsuGNUc/pfeelj1gv7oQavRxq221oRVx14y0y2oOlRHjfjuSXrijsinNSfkC9gHo
ZJQvlMsrzz2R3Z0UfGtl7pw2NXWJG94ZIRNrb/RorHwyg96K3vWIsNcAurEVa1nRBH+yUwqBNUQE
3Po+wla55igCYsEa6Zkk3pk+64VzBUwP3PggcraHCwJOBjfui4VxZ4iylNLXzkTsl/yTkJoWs+xY
Gf7cLN+fDyAm2pMKTTXjN/YfrJn4hJyEBhgZTAlw5ufSEEAOmfb4SnOteBHKmf1uQoV/KYhD0jv9
TMbiPcDnqfLtJ5E426sdA9BEOvuQVA1dtJcFMVMVP5Mwgf3VjADIBGPpvLlXsUuW7hxbLV+3zx+J
a/H7t0bTjoOYJHJdbk6KdKq8wG//jXsBzIxXuapkDIAJu9tKE/uTAmCrpOKZV/BW0SK1SNPCTR4G
+Tfoyqc6kJ6lohq1h8H4n/SpQGDMtZs7G/aR+Iq0huYtbq+VfDcBQDZlhnUo1oILqmgNYt0EbG/Y
wF8UjhtsH9+0ZTyPTayU0zoXLTsBp9cWyGQb1fNz9zRvMyFn5QagROiBEE4umzULe6KsWfkzqvx6
V2UdTG0LiVr/Ud84XVABfwMOxJgOoB1oSwYSwl0ldZbvpApnVAfGkumywUtk33l4EMqkZ0DwBlka
la7GzfPdofYFaucUnw4Ilq5DhnabZGDwZXLdioxptI75KU0no/nH071NzLWZx3FT0vDUA8LxWYfC
nLLNss7ySd0Q5RvgFOne6ZYxaQn49Nz8EjdV9XwrSGz5ZWLO331staVRVrNA+HppcwyebvMOOVcD
eNkuhNVRQz6aThTcT8Bd4UvY9o7EUea+n8dZodhHFLeiP3z9gq9ml53HwKqiwzruJagWbXEa9oQX
bDQiu4E9FLHIXefBskw07a5lSzv9GLME96i003Wc5Viww8NWFRz5BdTt9ftJ/nrsK8j+0qLGigm1
aPa/TGfLbGG5yQGpMIXdFvvxtHGNL5SyZCjdUQEJNGomUxM/pJrcSXUP4FXo9O5F/N0BAi1Oh8Y0
w2zab+eJbHybhKagjwLPwQAFnauzaO5azxEBnLjy4xHHV829c6c4JKxI0tc9H0929dB7X2kv7nXf
ypArGr1/tlvGBROctMnwxJKKV+FkxRb2q6HQtbkUt6prIogpOXJ5lkznyiIiyoaZUqdayTO9Ec9s
VwA/q/QpbnZeK1arwzt8d9Vto1mk6UP905NCYcN6rQ3kfBctHSU7oChJOHRh1vLUYJwoG5nEJWEy
kzCQ+rI7il3DTEgJcFhV7C0uqD5fC7KWN3t5PrMB580pWAp0FiA2Min88CuwXdyHRc7xEKqzGllW
FpTOSy9XSES8/4z7EQzg9RiDAwLOF5wfpc4CmsORho8NdyAuj2TYIqubC7+Pbc4KbRgdYa5pxfzp
vo9MULBRtPrjw4ur2WMBSz2WyTc8jZgiI3xjv2B5CitrBuU9RXkp5W4YOEgMSqUfl82VISe/+5PZ
PqcXYxf4mtzRw+XexS4+PIrNUgv9H22rwbTdvThL6nCkTt8OzW5F/SjSS/6MxdPnzCtDrP27J653
oxWprf7ytx+toVN1QOOOyJIYP5DrOGQ8OIVAF3mCvC6T3leUihyESV0KxnDY4W9rC0T995l9rwqG
w2z4Nsb4LlWRzl2Wn840u+MsnXdXJC7/6FDNsacWToNT5QJN5Ck4vMiWJEetgOjsu9nBfRHrRJ4m
0jcbUrsC7xtlP59lEodTjV3d9+vs7nG4ebEd6osRGwh8bj2y7ShnMj644FgobDnFkHqcPeH4QXF7
JMS3nCHrJekuytyl5Y4EU+dNT+p6m7X+rEbJzescwvpRESn4bV0uh2WPsYZF+phqMvqU9L3AqbzI
FMhuXUo0oyeAhXhn5VlVUy0EuhBzSgGGiGgcxHAqY0Ol4v9ZDSMTTrJW7Cxtebgfi5hU1jJ+nVwj
Lxq4ND8s37O9wZQ+KgZea0+UjL1jhIo1poferQSxp0nN17QIGpC4fj8noBEIV+h48XUM1skZuvjR
qeFI1SgP9cKjMVio7eYRntq9j+YUXvgvEHDRyE1xSqo6xku9zm+SUq/6ni4cR3NurLKaUm4RtXFu
XIPapi2cWlfY8LAiX8kAW9xWQzIat3n8db2CIVlglVKO/BTCbllwiObCXAcXnfFBEfXmTXfPg4XX
q+tT4/LYCMghXf0CoYJY41hMuaRjAgXKV2hz9x8QC1xUGqK8jqt5EykloxLvm+CREWh8gNqdbgzS
NEg43mAG1nmmBlK4BqpsuKOUb5zgQEpVFk3xGpjArBkms9Hl0dk7h+lKiPADh9bZGobUA96bg1jB
dO8vxA9mwTcdur2JLKSysRdeFWIaiYBbjZpkiqA3HfEdE7y3Hxq/Q2ydYrkgzh2bGmx8xI99C2hR
i5Hamy2vuUkvViMzRHYdclTZFI6H5XpTwAFVHjnpnMh7ESceBDeLzqfC6Plr/kfEuX9EoSTJAxDE
LX1c9Jy40gvwfYLwmSxtBLRa/BoH9Dg1n9EX6t5RkOCShwFInKrb40dm4200wDuwu3z/MybpmfLG
EIk7vpZ+rMdi1LlURILmy0YXTvAJE3Ui0HiMj+FxbbmUubSKmzr1wxjdiD3QU28sLlYC+/y20P58
FZxSZPUOX7O/Ls7x6qSCaR3GgQxIVX0kgW4Uta4xjWErIR5y/W7iqzf+ziviPcBjoAqJyuFKLV7k
DvKi0I7iUDuQXhxfy08vQljZ4PDxJNhjSWZ1bgmR2DpIVThHvhDVjZnk8KtHx6CWrXE4zkmpuGoE
0Q40Yra6idqJhQPx2f2Ol9hWH5tHMO2pK+/MdXvMSsx10sl0X+NvJ7s0qHJWOcA1sw9mD7WbTmpx
YgOW4kRT3EwhefWWFrtTp8H/HPcg/bwnYld6eOrK/rzaMmQ+ss871X83C6lCdGAu6a5ohi70HR5a
jrFwdn+fuBG1PSRWGODThIKFv95WlWuK+5DDTvRTzrBF16v29+7yjvXXn0HNW4luB/QIqYKZrCYb
1ecCeLMrK8R6C3x8ZYZ2/fF7U62MeLCICI9YfV/h9Wk4cF5GuQ/lL89v1DLqGxU5BIKDAi5aPaFS
NaPb7KRfKTUIs40jEuaeBtbXk20fm8cFmulNBmh2U7mH03mhuH4zEquUSSKE6N6jULN07noEq/Rm
g1d99MI8GfIHcqAUzmjkdKUgXo5HvqDA5wiI8BZThGq1RjApvGhqyNxeHHuEJwWJNev2byS70IaC
yWaq5MWymVNmuafxknk7Q9fe5I4mOYwTJ+L8u/o1R5mkDp7IKtcO2W+z0coNHL8arA+KN1f3uk6x
UORxf4am2XURfnxqwkRZ7xtL0MXeDYmsffFp7snMgYzr8OsQCSOM78xzTAEh7d0pKzsSZ3UT8a30
5qqNvGAI/N/jaN8k6e1rppJXQdx8kv9q6qv2Jqfl+HVobeLYMLA8SD1cbiOYOPmXr5Fun/LtgE7W
TIUNkXlWnW810iA0adxtluhJchSA1lpEM+iaf7Zi62duCE9N0AcfLtHlox4UqynEYnCMTPFokPZg
MFR+zz6aKKOdARQu47UCXE5bkGZ1zA8DDnqIhxFLDmw2d3pFBcvny+mF4zG5wplR+p3x+PJuaA2Y
RbvrWt2gTfm24sOj6HuSlobVYGlRddvWwhhxqqazVEsr0It6i7Qi0AURr38kOzhiQr+nwaU9AWa3
Z1S8e/2KdRp6hS6reuy/3oUG8K5KKhzto2nvdOkajd7W6AKsRM57SG2C7SPpMoQjAuNGzhrvJvST
yEw8ADRhPIWYdjn4yt9FWCPpQy9LbBNHHquSdGp0A9J+1dnex3vuZbiM8KWPDR3uVi6+VXoUItxs
MOkSNsShQodR73jXb5E18jG+uwZVHWiRVjx1eSjyO0RLA349FnCIuMp8UG1ArAllRAUfekw3OxhP
RKxWf79agTi2yt5wYcrQ9jivsVdADEE0ZRt9SY2EgDwWvwIdAc4ZYtQGj0rnG7hI5oJpKHhgbbG4
7UULZsE7ScrufovSDWeseXvQkFEEEYRwoAjMp0JvBpOIoDVFRnTs912MMdPPGu9jsNAfjM8lB9cf
HNpB4lo02MBtj6PARUJzZ6Wa7jd8cz8aoC+iAq/uFrd5h1o0WEL3QqmHz3R+4SN/DUtHbwnn0+f0
zfSYlI3oqkm/NC2Dn3zE88aQq68Txf0bIU4uV2dVLDuV37pvMMU5W4N2YhTsgVvvVGSlNRcQks8y
MlhLm4eL4T8byLiOQQFY6YxHk5BOPKxxHYyUfDhfaGRRnJ1Rlxit1SO/st31isauqvoszEDeQ/eG
EbX9hVBOjHxY+vrJaEu77KsY/9q9ZgldyssYJvFfUxiDiSjRJdF+RlqBNwQOY2ctBXbf6akaOPcD
mYn+p+B9WRXWNVvmBBqpvE697PrO3YvTqUAROFCvCcOHhRcCebZi9+8JIvBr/ryoE2V/ha/mMknr
SjYxp72GW10m7ukytcDdETONZL+lVcA5wD2drIprTPewEMJiqF4Njd21frWRlqX522UdXCIdx4Ur
KtgceehD05xgsDY95yR2JTrz8JGlgBLuyDmRUY9vxUfbUVTPAiP48kZ8jb2cC1XZOjUJaPkq0wTx
lBGlzID4QavL+x15OTUfM1tylrI7YJ27LPAbV3RPvGTkFDKQXi/22Gcy7tWtKqtH33QmUwGkGKHE
IMdHVHL0K/OOGogOXUDWOgXES9DQoek9QI7mzuzBY3D22PgPJS0DdR57owD2AlIbS9jinMoLnMl6
HOGu6DgbIff79VSgx8x4oMIGgT5xtIYKUFJPUEG8/qqSveRUnuvbYB/zNjkZN5fTdHPvr0JJ6yiN
k2AsyQNr0tzLXFPdEWd+MH9ZkZ+wi6ecd1v2l2vBnkQnoy1xnMJyA1q7zerRY1D/4zVSpzY0+Gvv
5rt45w5AaEf5WoyLEk1Q+U45O7W3Qnd4eYnVRzxEYlZksqbYHi5VBTI1JmkjlBrcoP2qHez3eQHk
Cqk3nnL45Tv58f2PNcnVw19MLa5FGN4sDA7F0IUxJaG0xNP5ThntYS5Bq3/cLDVuPIPFXdKyVw1j
DMs1yKS6nht0totmd/hGqcYlXHkgN509nT1E7nhuWeb8GlESL6as/H4/J1C79/BDn53TUWvtqj/K
BKgL12hRSjpme3jTdsIbVzZEWQLepVW63LluZpkm6wxlUtjfOwAChz6VbtyV7QLYzYVWmabCofur
B60s/os+0H7QqyTbJ8RQsTvMe8dKV6hi3VS6HWn7TinOggigxvo8MLWk6fwowsrvHf98BIHciXG/
8oR/UyUSbV01PTRLPnpwUf2NGJFfdoHBZte0bpk7UoMu0M9O1X5jhlorJf2kgGe1GtSZCcjkSckg
ZxYuNwssH9DQSnKAQCM3TyQxAWZ3HtnUHJuanHehXmIUoG7i92IxDGEonNCLnXYRIwnlnMha3c1n
r1QAYlgfwUGut1HLJaSrOT45d38Ptiu2qQ7bigJpiMxBlqAi3ukY75w2M0lQTLemzq2/Y4PNzpgI
CF7U6MY7goGwRcSCkcIXDqvO0R/xvdhLKROJ7ki/kRVN9YS1wvGPjaZ0nQlttbplbHv90MSw+YHI
MmdLKSM9oG8DzmVAk+HFx+oMfE3Dhw5TQrR9p2wEC46BWWZ6NNK+iIeQe3p/MwVleyKT7ynqNeOB
ONlT5GaG0cKExZm97FF7WOHp299h+8m2dgukaOOGfIUt/JbYlJl6tuqzKV47+3p1q+dEtn176htL
ESiI/hNBDHFnxrqT8ODLzNC7bosMFsP9iXM/YYHif1+PACPSeiZHUG9+m6NGFYp0UOM7qkENlYZ9
1Cvvgz/d2bURf3WA2CLjestW9R431mP1GVVK9u9yd2ebe5+d6EQ2wZsXXpjAQMK8dshqvqXTpy6m
GeS+iSRG4WZLbJ6wZ2jh/UHL+815Cv/C5SvXN8JGl3prrj3RJsehoEoJYPT2no5U84nQ5XYX3Y3G
NO53jrpEVCxY7ljpypwFq3DbgtRAhHmfzlHJjjY4CbkAdkD/IOBF2YnTKmNgKnrssGpG2q49mLPU
C3bfjyIP3oXLgld3jJZ3CqJuHc0bsTepL+XmEcBUoq1EOweLGDy6nxokS96WmIygDJET6tDKM8/t
0s8jODAqdQ47klSoZ7jZm9jyqBTb+pOxGHUYqwNvWpTQm/2/eq6VMMieKtR3MKjazkIWYoIozP7F
DEhY7r4cAe/RJz0uhug3GNaXdgn6C6u0ephav+Npm56z8cOQcIzanPNDRJ8qt8vRKxQwaUwCsjIw
qDx0xS+VlaQzHt8gq/8Nqujy5NZGGt/Ak0wG/OlGetTLcNHj4GhQVMr/ybia3LsQwc8tsi7EJDsx
+VKNB3zhtWBORsg5wd4TSGGxY3Xtkb4JS0dzEGtHWSizq/LNZ6ehrJAKu/EvZ3osYM1IfpN2fsCT
y9Xv39LHFnbVDjT25klvcoFy9N5lYZq0Yii53d4R4XwxM+nyYAqPM2MINYyTOuhsL7qNZVB21Wdi
04QI0o+xi69lZReMsylBMeSQh/0LibfbgEHUn79kyW5J0WTMhnCGKqKBZlTCgpkATezx/MqxbXs+
nkPbG2wpFOG2J2AmrQly75y85M8gFXNNSccbmkDCOPIVxRZP3v3QpBrXz21ubmoV2wO9BA6W87ck
XRW33ot4q6VW2JZN2ZOPVQ+6fmlNKJzS6lOFoYUgdI8SpYmXOoekbwpu0/wYsahSP9zpxcIYvQhz
IzzRqVRvvxuWA5b424wNySDA0tjSS4Gcip1yqSMqxyeULjws04IZ3Ra2mOCXpfZzgQKDqkoqN+fU
N6myYKpxrJpgjbK47X3Sq7CsGb4GTX5TmcNNBVLwg/d6QUSvgoJuxzLfLiLPvj5ror1Ikvm54gCm
F4Zgycpv1xftTFC22JW4aUq3/qn/wynlXR8eZiklENcSJC7TliZhdnFOEiOpX3Edy/KiE24LZEgF
4nv8zCxb7U6F2NXCvwv1+nm3c+OqDJh3R1vUTMn5WlTAAb6CYmmAHupq5WY03kQbhMmctH6gVcpt
6dehLQAYBMv1aKVVWWpbOw+D6qmXQKLUtpFPkUHq7jidmisVWvFU6q0re4h3SxuoH0aB+hKOSCD9
hfUzVWXCRnAOs9ZCluWGpwqXnjjFR0wflkZJ57x/cBTByWT48PZ5PDLTzD9PBsoG1H7fCjcoTUoI
+HGkOPhXYD5RBkBPm2Lk1jPW5GtWv9JxGmq3v6VAdKeudsLlrnKBpIWXGqSx5W7zOmdTSZHFoR3K
L3FUU3l4yN6c2Ez/o4an/qfjKg/oSKS5l7AC5kNFMcvfMM9heaxs3ytHqOF1HM+vUmtGjp4oQnR3
BeLxMVsuLCLscNUIMtLG91sK2x42pM2YetwGQ2y5JeWXzLKjs4G3KuZePWvI/IuPuvwPrXc8Fpao
VvRKH9oVPAvF2JI1Q80zI1RCaU7Twr8NZkzsst8SjydxxO3hVDiQLuKAHgPwF4/asspXFh/zULVS
dgOSKO2iU+uUpnffz89y5U3JC9bMWZvBb95XWJRJv/jcrf8mu1Kv9pxWhbmtt1PAeMBpfgNQI55X
Jxgxb9QO2EriXuAKWZ1NRNya5sARTDxx96/MFDt8rVOGKX+dYnNseazjtvOA+tgVapBaA9QrkuP7
2tYK+FRNoGrvpkw328yB2cFEoN3/VL3/fZ8f7s9S8j7umKI/uHY4MOKj4jIMeuVevimxZlwWy/bZ
BIxoVZHg/6q0wtl2OSvykwnQY52mPoiBq74gc0j/zW/GahP16fBA7UoVjhaat5Ow4cgQiZ6ypHbN
S5aHANWyv63C6MoG9mk7F+MloZhZwWNTazkRagOb1O5MZVkdHUgzu1PRfFbLqNMTKEeEzQHuDY59
6GWoAiHuHNMRiG3Lc/+MSTj5b/spmskHH2qYV6gPJDNZbFk8tMsh54Q6WERbxaTDM3+EPODkkEfF
vTrIP/EWObbV2fXGK5N8PaL9WyZWmkNl1zZHlD9t9OnchUDOWk/dR8E8JnF/Ww13ncONmLl716Jw
Y641dkxfTmXHsjUEyD3gN7aQ+Gn/qiQXg+mMoTzhhJm9Zy4Bbx+KthiOduX7STds9NfizaBpadyt
Km06a0Y5xF19Uye4n2STlB8ml2DKEglLiTLEYFlWB6OAhfsZ/n6vkhar9XUnNWuPAgRleUUcooK4
NMXu5Dgnphfp57/UMPLCsWickVwK7nomLw1FqBIoDNHNXc0+FHk8fQE0M9z6j6JF0YtLG7vlRnXD
Ko1ivESeFn9rqB21/IjghWDJzniILP9Pa2/7jaitM2rADAC7Mig8MLTXJzCbwdKACkMZtdIUMYyM
OpnsooSumQmsBHbzaRao75YrVHNbik/W4/8Perct3uLA/iEAf1T8ngiwPtYBhYES27X4IRmkYaTN
jnyerTNLrJZBk2C00kOV4LoboTkmi23L4CdJ5Lajg2iJ4PNNWQscvQn6esmv9uQzzvIXulcEF78K
GCIoZ//Ve2MhHiJwYfbXgYb4mU2R+iGRc/JddJ97Bfg5DpxzJlqux3Bsk9aICZ8nEVroa47ihW0G
3FniyJM0GWZvOPoxerGHFeW84VpsIt2WiUPtxKiXjhekUjr48tYHz7cXpzgnUq+lTrQm9aVH/FKB
5Uc/fEfaia6RJ2xzTHWnrEXuWGKdZlWtgpbkW+h44jXEwryIMBSwy0eRfpRcJeZoipK0kJXcI9wW
GTp2vg//bUINztk74OTZiYkG60Le1PX64tuSpKbtAv5jkOMF/1z/r6JGnba8CN9bZmjS+qXaDv41
FnMEI3Sd9G0QeeTT9wVgQMgVFABOTjdHrGqIjNmAl7x0gu9ohQiiqBbS8xezB54kpZRDBj5eV9/5
6ylgpWHjnPwjMNyNyon08YkdgjFxKIxu3YU+5bdllPSEXm79nC0KgRTpXeJcBuISILWLjb9E8Xlc
s2ll+2u9b53NWDbMZcPAMQIqDR10yQJLl22DfER3g0pOkBiHoTz3NE5Y7/h2gEo/MZamCkkuc3OJ
v0tem3VVNnXRt8iQk7UT6LOQMSe9nG0KewHGQzUejGXLHSkwpoOh2BRqbrQaEIzPjc1c+tyaHerQ
0AOrR+VqcbIoSoE9SkobWpy4wYRJNdojphtkrhINdYo4veZ2xQuAklQe1HCMLcE6teKYg6ajL5R3
6hdUriOaS+yg24vOD7EmT7xRwhoT2aMhsTjNlcvImZsE3abHZnA0Rep2xSHJ4nk34GyIgfduCYZ8
SqHhcQy30MKlGx0IAToWAQPV60wxvjFsK5CU5/NqO1wvx9MHVrRuoTVxieJEnjPPOIIVRl8x+DuR
WS8DYFnx2mtGcjJCCEvxmveacvkUPNMWUM1LEAOiJgU05ubZsgVfOjaLzeZ9bI8L9HvFXxQBy12z
whX/g27eM+65m4eFbxurRdMSofokjhZ3COLkAV6MenIm6oIOR1QLtmEACaWLkylW4Iit/1m+sCHh
HUNdFO8zgK+2UH2k0Vsy5RH7Ty+t7e1WAsoOyHgiR+z8i9a+Askd3sU6jUKdYKnMLiuzq9Ib/Ql+
udbkOFqMqz2P7d9vAKsasBtXTwiYsPh57GZLldH7KsCKNUfHFqTMPqkQYIkSjiI8+whd1mnSZPnU
mFow6RIyBc+f8xactTR9fcIgc8hfrUse7NEQ9BAhVeXRdZdOOmxcThYSp9BI4RSsIX4Z2GrJWhsy
T5CTnKvbMv4RkaYVgCyVUQ71moLHY5GVJADQ3OPs+nANhAbjZP0Ew2NFlUZsAMRfJNq8spcOC3SE
o+h1pToAH3EqToJTf++Db0bPJojt9S8FT7Fui1Xbachka0i7eIPnP8qRheirsLxnaFOHnFhaQwAV
yw/J1X2gWAjTDhjnH7tfyhmL/CY6FJDgHkBA+K0R3SX84+QOWK8z4JUxihflMug6EtEQ5i0rWIRd
rVBh3LylDHOaUSjip1YOsoQoZOk+AKebqxx017FQjAQIpdD2n1EqEe6KXF3MMfSflSdOBoZ7YiEQ
ih5SgnutRkBkloUHP90Nqsvf+D+AymCGd4/sv+7TusKWrPwzfDbEQEy0jVPLj8gqpQZHA+hTZY+f
waliWDwurB5/5gzWIdOwlHHt4Ewg3zmH+uaQdPImgalJQ4x6vH/4LQK4IO9AE6lsSo7nt06AqMB+
eKVO5eEUsMNOdbei18dn0S6yDducqYSyOqCv/Q8gtaAOM1al7iPa68v0I7xrM3OUxRLYfnjJGjXg
HzER03e3JqECvEuDKys1B06JNEkuQ1aslE5SJ92Bg9bHzuioBHvzLNzHCzhiyNX4EpRbqrXBi+Kf
F/BAgsGEwiCCciUKiIbqZJfbacZtsLur/9EFRDB4uWQAni669UbIIzlCuM7vHVa9Q1zNtQid+sLl
FOCK+xat1HrhmtSKS9G83zE0Qhicx/3WnZ5SOs8zwWiY/1YlRGRhmGYq7n/TCdTcOgpAlTngko2J
FEjChAhQ1Vzc5rV7SxCbaYpwJHjm1+29NK1oAQzGB/JNoRELU+bm1rb6qmRiPHPl/DATcCYDSvr6
qxsGr80N+xN1txDpdoaKRO11sc+v1ZLymxA5D56rzYcZ3WBai6pJE3WMvmuLpm3G0h98KJDZlHn9
IxP5M//4dRbxAQKt+gh20jmelbleWtakSuRYWvFu5Bjq57jWv4vpOWogJFxUmcJpOmE0bPMIbh0w
QaARdiCLjRckIBsItSmaOovAfN5gPFVdtQIgNNoGGzEl7skrBshz1+QYwtWS9WmStp/+gcRh+pml
9pfOHeATQA6xKXoxOaSFbPFD826hIgSV55hEu1IqQSc78IFAD0Mltsxk0m0LSvwFEUsCQ3pB9E51
GpQoOOffPhXCvlUB/8W0qi7kiQk1ejHfboiDNOAeZZPr1JMpjWGVXN1lHmD6RRFv1/kZStvqh+kf
sl6y4OZ7uQPth7KRTNHJoyFQUm5VruXsdL060qvvEEer8/0cbMZo/bDzcytS8v800Svt4VjnOL21
Gd9jJxZ9BxB00pF/itBFzSPqLk6ZE1HNJJY+O+wrrH86uKVmieTrYiewh1+Hc2+Ml6dyYfX0SDH3
CN9Ho2sLKjTLwC/pvbDQjIOH0IBHbrtQuzrHE2pDvf0QDIqAlVGgwRGPJyoIBMGgfVk38qiGsrmw
2VIR0Vy4XkovD8+ExS6G8KSnuruHXLT5/LCMHEsxZbS3VelxCmzZ5ueRfGXO3ocSdcHdv3cLhdLq
X+nC8lXPhixCoVhFEw7Xcw62HqT1It81+n+PXf4hEubBxkHIhYiey5MfZX04DDe6F8UeVfLDUfOk
81LZITzYs/vikYETsXy9+9vVTY/fdpbFy6PkH9WJFETYECbrrVzRVUbboBzGfhRcOgHYgh5/NI2V
RU0hAs6WkOM6MDy4THslj0UMmdE7bYgoeSQPYdg4ERBbZ+CSwgpxlcRAuHAUBO5gYvUysz7RTu4y
5vuDM/ePFqF7umsfyXrNM3VmKRE241mBCz6fr+GLLIcCOixuLdhRmDD5peWndr1zw7NumGbjoLUr
1nsk+zAL4xDNPLbVtnjczY+uGJS3VnodurcQBNe73qpTykDhPpdJAiFWuSNLI8fIVd+vv4npsOTw
CdDScTo1EzXmcpUHsX+4WxePuhl1MnhQ1CHthUXemQdKb6gdIxGtQeGcS/9zgxQYF1sQ/0MkOHAv
FFq9fxPZMyzrLUztUMXqHg/RBukStZ92rRlBNKXrd5xr8GSpEoBniXfb56vHNs/bzFP/QqLYIAq/
A9+7XeydQPgik7anfB6/MdWFTjTksiE3fTDRNUjr7b3Oa+I18pe0F7+AeyaDTV75xt0WHjJS3Uy9
VMzCvqIImhh+16dlBIIGdPQNOLgEXGdDufiR52erylll4EMxZ9wWV1BxEQwswzWL/dm9ZniDuWy+
9GI+kjmXfoUtiTP6QlmYPU60cvHSwQ1VqS0hrNL4wq+unNmqwbvp59s8Ef8fEy+27+l6TZXDAIkP
r0Bt4uAcyehPjLIbBeM13yiFh0+WUp17b8SDg3EPZ7JfDKMtELOJRBnSAe32vFUq0cNSUHvr8obd
Br0jScftS+6fsbP6OWeBOKjryNgW4d/w2WQ8eqBWtl8tnAEPD6BtteH6TuqkMcEMmTQ3PWAQX9q6
jR3t5Pz5m8532uc1ygu9dbQSbBtzRxC1x9YZgeYjYeuaoh7dS85KyAMrHm6XOZHhP0vQvQ+CsTIR
mVoXkG9I08EReOxMDvh1wctr7OEFTBpH2V926lFHcBNz3kWZ51wTUojeMrRcH2c/TBoadPeJC88C
fdvTdaQAvYsTAGNc7ZtKaJGHYKHvwrlPTqqd8QDlVox/oJQJGETLI4Ii+g/v8aCBql6l0mdvMtH9
WsFDCbRIVz8TjCPg0aKD1Mw8XkMmHdFi/wPXze7+h+ljlN1oJ5EvIGGIb6sa2Zy4qYZt1V2MNNRb
Ax0R3M7xRwV+3NNBljJ2O9xrOflLAvTa4aVWsiPKq+pXlnnYR90afgCi0FOEScmE4h9azrlWRJJM
46aoyu0vBk53SiAGw0bWW48fMGWH2IiWlH8A6mY8XEufkwD+UXVT+f1Fq42gZ4lGFEQU3+z5W6TN
WTZyED8fRXZ5+CkW5ySv8aBHqEu1uduHOXsoqrWdP1S9U82JG6QuuKphWgN71uAUcpSbsB3sARi8
Zl2yPxbO/Y/kpuaWj2VkzYDAfFI+mWDMx4dOivSK/i4zilz+55FpSdpQQTXxbOkOXARRN/z6gh6K
8fbmql8+qyy5XsbjnRAfNcckIh2xAkvbtOdwpPW4DU2w0n0KQqbbl9X46TNA9vng
`protect end_protected
