`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Bj/yHUFjAzUF8cEUTKe1/pZAeWfjdXSN/aTCe7XGAXYSniHyCm2v1DhSBJpv/i6mzTaRfGHd6aaZ
3tHO68MF9g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kofYye4rsh+U7MjByPV1y3bveFCiWxBGISmUmrbYp2FNTogf2y0ontp2OTeVoooBcGe22M88v348
SbeUEMJdduAc27rmj1SeHKe9TvRD9+8tB+d1hHOpd9h31xzKqQFD3UZ1V6qP236ZdfhMCtTl+MAX
4aE3FcFPEe5HAim6Zmo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aCfpxvpQDv+zaFXt0AL1Rs3PuYGSlAkXu3QS0xwmus8hQcFfOH6C84x2MMsbVjbBFVs9Gq5FnLwH
vxlY8Mc1HOmU4jov66r/oCY8wreW/5gPL5xmxxLRaXyUyWBagmUfUxEIFHiih7RN/I0AU+3/X6NR
0rsB4PAs2HlvLuZucOW87cAmNzsMO7lBqA7putu3Je1gX/hBa/7XUwINCuRD7Xc5Mt1nFYkm9vtM
EIUDyYI8VeEa32m2CDbDKJSllpYENi6cbg2bAUhtnC2JJJFPsAjZxRMwex8YS2PeSA9XamQ2lwlJ
dhTMA5cbWIYARZK5AgaEezDmSVoaLPrrZLP2HA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xI6YrNVW2xjsrENcPSR0T6a32c2BWy0DPDGXSC4fR27ogoaKpCNNsBSstqyozrdS2njn7ulV9StV
udROkHL/vcew6+bZo9Mi7w21Alz80ZF82NLJ56kBWybXvAaLBDLmI8jzcThgxnJHjAGEBPVa8Kq3
5zK8YY2/svs0+JUSIvc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qdUBPQkXcscSZ4PVJn0qjDfWKMl7N+Uw4ZYsaY6KD7VEiku3K+nZXA6TcmDk2W008Nitklzvh5+K
k/9Cc1ipQlXo73ZVRGPpjk/Jwm81nZFbA6pQnIYb7UE3YKH/DQTEHDziafJffdUG3eYhiH+Iy+cI
bKimXi9FptjU2RCMPI2ZDeRXBr/IUIUk+xSBPV/cwF8XIZjwqFZsxT0w2Jc0WqVoSrc2jIy/hN6T
clwUajTvWyTSShSX6qz0eUIysZlQN2VbO6lM+Quh+sXYktVhw4IYk53aXo+KSp5S8MA+FHDchrtC
raTk1I08NsmmoFN2pxzhALh0hd2k7LBeEa8i3g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 58800)
`protect data_block
tjjHg2+ebvMKqx3rytXk8C8FVV5wnXDSoSwcCJlo+dIxYbzEDby51sl6nA1iTs8VEPPmFTiVsPf1
tc8AAtLFym005HdA9tDu9/tI4FL8RXo6cCOKfyK9Kumk9bU9zFY7W3CWNDD5GtFZCAKP++sY70Ri
BHAoGfy8BUczMI52m+R417G5Vm+g7FB3RW4ABWl4bFyV/Pd4sDd/j7aZuGwBE7G86lnLkIkvKEc5
W9n5T+1KNGIzP6d/xLJ8T/ScEZfVl4LuGHZooxJ+uA+bM2R/GLoAXEQEZDsNqKDUH0fUten2SCm2
lYFJQl5Dr/yNIdNpVuCR8Ca2vw2lbwdU5WksKqMGzcAz/TlrWCbjAB+zx10QSbJFM7mQQUGM5QKH
zdxSZaxr0IvHfLS9q0mfIxsshhA9t3lcbL8XNkxttERPUA+66LCVegu8jITlqQxeg+az/92CTQY3
rsTq5gtdzT2DLmd3xQzjL1nP+yelMdMzC3PQ+aItHMHBVjRE4IEeQ+4e9/uF0+LX9Zf5UDBdeciE
p6PHT4nSzGVR2lfKGfCCfI5Ev4sO8LpLIe+Hyli3aKEMoT1bX9vPJyP+l9NAnAmg205bKP8184IE
pFFDZxPXxvpm9Z/JmtAdl0xtPQiFvktUI0Hy6xpYR1d6X9RZg9lrfrN1FrJjkjnzjKeZ3w9X1FxQ
jDCfDBYIOAaZuYEBLklun6rPPV0KgPT+jKpFxryEa0UzceLL8b2FOLdOhCovWCqlmccUK85E/Sbg
CHASNGWCbCF7ifmXqAK1Lq9ZVLk/MkyKgTvRnKRhtazpTe/XOMFUmrbvNXDVF176VSyLAHscpHrq
MCcADtK3dSP75HAwEaxKVOFeDsEayo1C3iQERbTdHz7wlnOLt56b+Ix2wdfmirQp9VjEUu0OyWQk
3H9e5YWmtoSkopCsFfoM7CPZK5jlHWogJnCwif1djGUGIRi+chrVpvYJGYwUgyWFA8RThfeFwc7d
eBkeWy5ly0UAtkxUqxyr1QuPUCfKaEUMO1KgXoU2YU6gQkIxxinjd9bOtdhP09JcorfHGaODmPtC
C7G4e6dcZrA+B/JUhRdzDNj+PUyEikGJSib2aX0pTcoSIWJ1FUAvuRdS4dxxBQ/9bKwhm5NipbQp
3g9Io5uKY31FGYccCVP1U5mtcDmFajalCllx24TGk4067zQhr8hKT3ik0s7gCJYRp8KnfdlrycTr
gRIbj69GNVKnECTVOPNNTOQx7A9uXqQ+pSScKxgjF5AqmVBuQxJsuH0nt13dNbhglr0YkNhlw3HP
V6luSqZk4QkBPmIELrgPCpMuZYuEQClV60q8V/9H9EHYuPENQhHmsH1tULZqzhj7+ehuHy04PNhA
oFxZTFgAP7wCC5UpR+fpjCPUGrKJMejmblN0IOTTPbOYaf4tlrW4EFZfQ/n626Oj2IzUDqAAWOkw
wGb/PJ/o6bKqYZ6G0tgNnvm1hVTh79f8FOysgVr6XR6uyCqpdVVgKgY2lMj6WmX6aOClwCnOFaYv
hb+ntgYE3GdI8FCCjtJ9I2xVGuxk38skdrBkwhllXXCTFKtk/YbsRWKHXJfoefcy7BzPsTVfpMis
vS+n2TFOPSVKaVt7fJ4bl/Xdk0F2Nth0c6aFJQr2HgAYsggGiem4oZLVZlBoiwjIEBy2XLKq2T/e
Fp9OTebCBzINBfRGJyKCwCJxKW+N+KEGmst9M1SNl4WH2lsGLb/zW/c06dYQu+vZjwLalEvlWgSC
Ih2TLM4FsUSF9GvINGPU1ndl/CQx6M9nAHNKuUDr5dyymdHgL3voSusLt8x0dDJWOGwqF0UXCSGN
8PdoeBRwYxl6B5+FP0OqIxd2/iUwrx0QWcdJtAhJg7hQDjRstsPCK8qzmmNVUDCefmpLf3g9fMDX
qlXYJcElHK6iP4qE84fEBlm5rn6SIdYF5wsFL/uWc3fGe8WruoX1dBGOGA3FDL4kfFoN2Oath3az
kPqsDeFl5zWH0wTTXrv+1Xo2zKL64pTsfW9VeIkt0OKCCjL4ylz+YQFXml1U3kCWoyTYEHw8aMiF
/Jg4i4Zeg0sS4uVm4Fuc49w3JojCbF3+Xq8uH7Wm3m8K0piB5kmcKuvm6RynYdTFZRwurR4ROPOi
tuN3rRSZ11JxcESl63tqzu/kc7rOLVBQkYyzB/zCkvRNzug9GnZveKw9lNbhwjNjzKIA/VtZtZN5
qsjQsqOqXWH0dRC+2wVVExT6NM7ua1s5p99vHClj7fLNExe9bMUi6927+rEf/+GdC5HHVVnCujaR
FV8ZU5KR3yRPV13tqy1kcGj9E/0oMRHV09vf+ShmxbnyR+PoQZv7GqU7IDCzZnOt9ri+nbvQ5UL0
fg0QwPlGtgGcBtE8NuPAHB4BII+iJMmxlLBrhLlEIm0MhOwoeqi+ZVqcFodmHiuj9GLcMPgioceb
nBz2azAX/NVltHhKf+rccF9mp/AQsxVjmeqK2z4spRJxU/wA6CC6QOtZ1ExE90LfMPBNRXm8tbts
uQDvXfTN8Yhcu5/eIw+T+wN5vtaCOj+0+CkF60A24SRNkAs8nVYu9tL7Rc9L9rAYAekRXjv4deRg
fycdwCRb+n/aISvyH8/F8dmcxHbn6f/Vnq7tkmMNv7PFIPSu1hGK5gEjP/IKXhZdyOJVEdjMMvDs
0RrdQ5BqtKt71/g8y20sHHflL0C2+OWpQnISqajTAubM59STWBgfcSvIfmFZD4hzc7VLh9EOpjzI
Ws3RgHwAOAWPO4N05fZl6f4gyejMLv9t5QPpzvSVPf3zTEBMPYkBjlvzumBdlxaSVsHUXWlwkf2s
UTnzFVkzMVopHMBReT4XUcMxzymem8grZop9kZbCiIJqpUW2al1xmIMsdxBMt/bSpxCUxDdelJvX
S6OXoplgupSeE5Q0d/7R9cHM4d70Rap+2NoSsFp4LDcIfTAh/gHxaMGeW6EeUHlPHuRkDuWeoAEl
v1kJKczHtzcu/Jk/+rFQWCD5k09e4C7Jd3s1rkV6NzGLyZnIIBJHMG4YnGQAUwNfrmFjRjPholxI
L6/Xe/AInB4M358g4t5XLV699xQakt8Ya8Q2zLY57nvjvXCsEsv5AP85t4L6b4j0zGfwDEzsiaVu
rwm6obVRZOyfwCZgyxM6iVuXRNNGqhPCaamUta4hT9vbhi7eBhXaBF6Q5mUTRCJe1l2mSWlhLMjo
lkk5wXYMjOkS+SLHgPSFClf5SSswZvaUz2+eU8JgQXaM6V6qAyMcA0rmuWQRMrZreBUtCUSrI6LW
Yx2j7bnukOVLfe8Y52VQTP1HPwwA3IfySX/6P+7XPjhFJvmcJMsQfNh+mU1CBdKqf3R4sQeBPmIK
DkbbrjbN8owJ8TJZ/vlbURApxsax3r+7GYSWSALB4DGDad6NPerOrhkQN8i5ecJzCyRa+ou+k+fj
tORvJJ21j5whvAQ7i7ZmslQ8hM5bS1Q3VhEVziyqCg16NjQPy3u6X0WaI1sAf3i5Nm9th0Urto/X
komG2hh1dpmtDGmz08Sb2idx8abOFxPQIt42JXuOPOuaHaRpcO2K9vaHHWTkRiwuyVwjN7E0B3xf
Uoqt6LMaHSRU9auNhhizh2UPL8PJp113tTJz2K79jvZ8tPngPXosHOVvjDR6TKcoVqjsiB4Y0T7e
jcxnyJ+jXgk6bIzq2jhYQme2gskQcI3eWhgdg7cLnv20DtfPlL81T/X1kj6GmDqEnEY3v5qTEDGH
+0hyf/1SQBIxZurYE8n41ZzxAUqSCE19obvQ/ZLG/inQraTCvn3N39mnFrJBd7YTiVHh9a6FMkV+
xHtsVgh2jYo1HuWqEKf5zTEvoUOQxozJrxPJrgO+/wwzeyeUe9W5AeWkj3EsL8n7OPVkJlAq58/U
9M36ENgF7CCqRB4qr74YDhJAJPjqnY63F9QGTA6HmE+fZvlAYjNM5Ysac0nJd5/FfAWnpjyMBGL2
Ay6+6vAFiZ/P1gdiDj+zjBjbqsLAG08JKuBWOAFVCRDZZGplE8Rc1/CP7269mwolD0EC/4MDBpXH
Ima8zi2UgNfr6H4TOrwOpixzZjVqw7JeXYQhTWgYKyhKpQBNaQlNy3zN+gAX4FVTXE06knPowloj
lriD6Mr2w0PPTYOeNkjfLYEhQILTHcqOppftkTUjJ2FPFmAu5EzSQxXVQ76rqKzq7VEO3tMAzoO8
Xe8vzCq2SmpoWTELpGhl9Mg9ijOsXyVJUlFVi3bOaAvDktl9AHMvMziHHyWPLj7XhtWscL+iVKxK
BTWt9vDntF4rMZD33k8vPrx9dNzrLw4MBesbMt8G7xYu3JN0J6LRExSvphG8F9raf7x9c2X3ExSS
rYVzAy7KzYpiqyLyRwLRnDshi93GqlKRTo47xtQNxe9PcuUz+Morp5TmIdsoW8EWHboGKNun9g+e
T1xeGaBBSrbJEtLjmr4yaSOTj6p4n2hU+gX6LbOFvODvlbYaIdfbkVZBpTdjeEPMQEMIbVAuTbeW
CBQw/odKMhSpS6OV9RFYxbbyjm5HGDYYQHTLfuisyhDPStSAWWYnJ8jK6S7cLkpwTGAr0Z/lj8zC
uf87mmnAUDkR5jDto18Mp9y3szxR3ihSluFxNcz47vQVuNSnDzcTU6EJBCDyLixEf4q8ewT98FiN
ZkCm3emlGsn8xNt4qAZxwxuEgKCNnkkUr5QS9tsYsFNMu+Vwaw4jpKnEmCYf7/UAUxYaaoCWb9Ao
O8UZNYCzb1OUCldFbk+REVQ9IPFKWAs9PjhqAYJ+AE2wB16LgBUytbFZJZHgFf92Ay5IN0dQtq1k
p3n96GP54y4TClS+oxfuYg+DXLYHUS7kWX939iFkNPxenlRj7uB/gkzeV30xMA+p9sxTCxJyUN/D
ToevSC6n4jbn1fcBYY7riy44AgGZrwc64X5BfHfe+E7phgo6tPpOYMqT+qrMkxGb0d+lgkOqL6Nm
MFaXmRAIk5wKMZObRCwr9x79FgMndHCmRU74I++B5olO0F9HkLkkN/gc6QzziFWB2VJXbzaWSTGJ
OsbvZ9zIjr1C1Mc4j6PJIpRbo9j6obhdCurL6k4rlzhIf5vpIKupNRQ67tlWgc0T+KvZD2IKxoc5
cnLHjrs2tIb/QttR0CoG2nYbzL5JJ3hbhGYiqnBqSzAqqDGPZ/VgVWI5e6NW0QHHNt+6CcVej/cF
TYEeaqAWIWX9UvZYaPsyXCE/udHP1rKXzXkVB2Xx1HYRtVJWnq6DhSeRcPKTKIxS+N1gnHcovYM2
6uP3KThUk6NAiO5qnMVQ7ExZr9zT477fbcuwtfrAvl8/XXXMYHvXVMGrJj95tMVUT+nKTMq+DDEQ
RJ7cISDAlS437a7vP+7oypMljsduGjJWnvouqIZu02FCLaAVgTMWpxZkrX1P3bWxdlDmlDis0Ubb
pLWLvB2DSiuChQ+IkxA21k9EhMOFG7MgHmU/XCXh1s1FQvs2EvxIw65w+tMkdbSc+6VkC2E2dwlT
rVVHcyBdLXnOX/EdOjMXRE7XBTV3pbcbyA3w5S91uwDOk1pzfhfz7s8324yDbfhCB6Jh0xDfkqRt
99Z7ifahw/P5Gz9bolmbiJY5DONoZaxTVOhlygDV0tpWc8c/7luo6fOqzfDvfcYBNyd73WKjCHtP
4ZqVzRmL2fJdsEENHDxWmShWjiIkDC4nUbV8FMjcfaEjekM4Y24zID2HJZP8DW1Q4f0Cb7te0uUJ
fu38BEA26y0+bvnG3D1dDHEw+EAuUxDpDz2WCSz3fiYr+5xhplVX3NkwkcLl1h3m7AH3Nkp/oBMm
o6IsnZp/t3A010k0jtBKi9bU0h08BWatxep1i5BZuKbNOV5Um3wd244s5+/lWGNIeO8QRjxIb6RJ
poL0s4Kt4JJy/B6T30sWSqDomVcyKYVSaNhGQwMycVpizyv/m1ALfpqRnaEJChZA+/+zkFfAxeAG
YCMWMbb+c5XrWWpHjIxjaAxF5I7epmrW2v4zxFq9NAMwKNv0hzib4wUG+9KEmZEkFzmV62GyGKRr
oNmQ65+UxQt4pVs92Xt0yMTbdQk8AM3aLR2codwIoBBhygYYsPrtwMw5CBkT188yGW/6dt90osM9
DfZ4OnvMTCBMwnH+Xjo1MxDx009YwcbiNe0VraLW2GAfKFbzV5Wqwt3SHu1z+iG+qxqdF7d8Maoi
OX95EUlThop4ZOcsSnXAP5lnYAxum9jvdlBQe6i5Rqf3BzpRqCqilQJkxwFyguqmJmWmB+/xKBba
oM3lwbd/gz+NfpGmqHcTbgSyk+z+Xl/f7gddyz2vQAxJ3TEn8D7PcSJMh9Ii2Rj991bzchTU94lB
ygfo/Abl9wsyudBvz3Qu+QKD5PLnbo7HWJJnKNgqNW4lTjaWQ+V7UKfn58LeH9ZnoHhwXBQ5GMvm
7Aw7aKN+5vp5vOG1DV7CFT2h2QbqvtQngrHlgv9dwlbtNrMgQ69HLTAx6uoAJF8dDAgFO158xhAn
lJW8uQjMpKZyNk/H+bGrXwh2FUF7ih/Wd1J2VKsQAHIHdONLLvK1M1cAeqDgHt+pNE23+mQtDdGL
rO5WwDzLqU8yZ17Osu3RMp4ib/9NH64e07hzkcvrBQ8bg7mzHSF6YaLHfaBCymzFyC9yEw0RIWo0
HZyXbI3rKajCOB8dWA0KAv1OJi07Hk1u6f65Rwbqi2HyZoEvycewbukovLn2M22qtneNA0uYZdLF
kfZ4gR0Z11Pe5rrbqXNqHG5ns8DNIUhrPnK0K37F1VwPEq3BxDZsGlvo38YOQgqVqjX2gvM+/bmF
7hC0BXkNW1q76UCFIUHfrV5vtaT/olOpIvO/lvSZCaHT/F1TBD7lfxMtVuUmd3ks+nhceVvRP4d8
WCBIIVKoA2Ll1uXeDLQmiek18T4V9KqqqZas5+72bfv5V7JhSJZ/szggQR51DDMHZuBqg1Lb76pm
DHwbFxyYdlXjH+flS7pHBoo+E53/rUfOHotsBN5+Hap5ohG0hsQjg+ovEZ6xeUlXIWzNBeh7JO27
CVZfBePColGXohb+5P2L0qj5aANF9NeL9EjrtqV+8qk6J7S7mqvecbljecB8KlHYASr9oO2cSVUf
9uD2ZfMvPLtguoodKrI99TNgUzYdvNlxSBopzSv304uavPEyC2D+6Eas7lnoobJFnDaaD6j4C/uv
TSAHtqw9pP/AVMlHhCkgc8trTb0NLnFDfkwc6bNUmWpJ83MBmGB+T3G1k1QbMJrlTHKBj1u2naNc
fPXiXlLMVXiRpzXb7loSdH+KdwAHms68AI3oid3+uF5WbmF7vPPn9KiFHydTYoG5NcFefDPzltVe
qE7Gm/5r9Gjc0Fk5/vYqsxoDmHxuYJImkEf18JsdVE77TGPap7qoUm7KNVc0HNYaK78wbPj5Pxvp
UScyW7QnOck0FLOuhGNW+W2TKfkRZbZ2Ahz0j2xW7ylEPkm+vfuD8Pg6XWs1zZZ4lAsoG91Ej726
65eTRGTajLLUp7Aqg64BCgjXV4zw7zZkynCa/P/Bnbp9sNpIhAd3fCYerEXZXVE4DH89a6TbeLv/
x4uMCMwgycOKb1PXZUKYz5hNnEYrCWMRvsZuUK4sxuC1gEFEy0JgcHVShC9rfJKqYGlCjPO5i1X7
JU521kgNnPtgv8d195l8az6StGomMX7n4kO2YSiyNyhDlqksyBZMUgjTNJni7o352ccL/vDsxhQR
0NKjJzeH4gK2y8AT+3HJPeLw30PEHvubvQTzdRn2ui9TI1XwJWe6Jw65Wo8M6bGe4gb/hXGBYxZB
WMojZ4XpAVbbmvNwKJJKIplC2dBE5ITTANpq0sbCMsNP9UiHNNHIz3gvCAn7V8cZRaH8QhRH4QEh
UneHuBFvrrh7xYlky5j9SeKg67OdMZts4YJThISKFgx1VzPtjWUQaOisZ2x49WtvjxEIggVwhtez
GJENRef3VmHABfE/rtiy1/Fjl+2lyCQ4D3NnnrED/DLGxKkuXVbZazxyZtNul4P1Ktag8b4KHdSO
wAjo9Dr50ycWKCF2sctYdzPscFuUE1LT9sAHtJnspMkUGGbHSTtL2SZIlFQCW4dPh7NKimA2t+3h
PkWODBYHp6hsXrnAxhqZPWZm5mG3Pp+COHCMEebqQSdxGVl/gFT6BcCXo1ZpfsBe9Si8AwviVzC9
ZqnXekC87J0jdq2KckHaNe7wvdL7zwAaHqfQtRARE6hSEy9ct/nnft4DEFQAKPZSne2ZPWlYZn/K
8bxKnhy4VLf6JFoSm84IdBmaO/akyjAzOKqos4Yzh1yMteVvjpTJ1iYQYbOJZOLbSUYiXaKTNfri
yb2p437YZwjrVN+Oanc1kNSLqkknf0q+moIxV8t4BBM6weXEw+Y5DyvnML6dla9LuLsWZ96Sssiy
uC3q8oi/lrTVFyQDB8HfnclBEotKMvUUBZF0j2G94gJB/aCyM0bBxiR/0/nRWqyuEpknYRtLeIDo
rUsB44neTgSGSyx8OXoIrzlPxmTPE8iGgovc0Vz3yFwMPU7+C9uR3j+lnsA4hnmwL/r5OLkjkq8S
QH7UV2/IXkKbdIff/PzipIrXuRIhyT4FbpkcPSDlDQowco4Xsie/IrDvaOC15ifXuq68JABENsL3
AgmYXWLATO27DLKjje82d15IMqJRj3SFggykLbDe4WQVOo6vl1uhBs6G5c4gdjJDi+dGvpM8YJtp
kaah2YMaLYcrKArEkj3SCDDSv9rU9XFvV219EbVogC9E0UX44+EsGmuqKT01MKBOuPRtXN1w6Amv
n9u1CUsWWy9Rx1Um6VEvK22ZuXkymYg457NgzfAGRMuVfVzBlpxOMDn4XiLCeTs5ocgF02Ki2ctU
sorP016ELhDQwEMyc20gftzNusc9KnmFVSWqE5ik9ZDmxcrAet3Kv8bfaofAUW/QTDcDk2yiQ20Y
bID0JCR++24FQ7eaDEQXLYEfDLXL2mBKjqq8KmXstnhkEsn0YIJs0+/idRPmHWmgOtwhuVJvqQj2
RK5M2x1WL76JMWuZk5j/mAkPN7AocsXAZd9MO/o8eFqNp8Fz2VxqMxbBqYaa0d0QfdFtplXMa89k
6jXBMc1PoUTWC32UTyluN1qxYKCQD5zVb2rVdOYcpPaQCOMP69Q8t4xCEwhpcd8RfYlQ9ek8mBj3
9y+BKpHDPtgIaAW3VIAZ5ZctEGt46BWQ7EG+q3XWzjMLlP1N6JhHrdL0zn4zpEy68pWiTX0rWcUR
G+JF98BsKllRq7ujHF8wo4P4MPTZxpg810BzBgACPfMiFzRlvdCiCMQkUMP32inP4D1nGtrbau4i
XJ2M3KZLF5PYAgqAdaFDAifoonlIh5kE4PF7knljkYio329xaaOpZPUkJE0hgFj/ds6rivwVviYJ
unHEcNGx4stI0aqv+OBi6Lr3uHC+M10mOolUTccjqN88tLSvI4VaF5ojMmqneKz1tw12Q4McE2W1
2Gsnos/dDyYIh4/p+aQB3A2YwGS4v2k3FxAEZC4/AVadg8nxjZSfaqfR79cp+XOHWiHU0TV7MjGS
0uKOND/1nryQzb9BfmyCaw6QAzXOah9/yYigJbqMpTK8G//Bw+v2I7CRYfayxCe3fssS4XpMRdf4
5Fbf2ApOk3frEMxE5h+FbitfrQxyUnwA+kAMru3rIxmVp6vF5y+Kcnm/Gmwjs5T/B6u1dewLkhlL
74AZ3eXeLR5zlRULu/6r+Nw1KniE4NAzBlYTtpjpBVzR8RaKVdVGCkROhjDCWJNSw4sLCfpQBC0U
hOFUdDAuG2eLwUKabx/X4d2OFsriGE2vrw6gDis6/qRGSG662LTdDSPyoJ13V6IXf/HwpSC07DKC
LMrTDPjdEOAdp5zk8TlCDFhM76UCM/ZA3xwCyW/4yxF80HjnN0zm93VB+54F+/TOakWfpw21w09E
32Ct2P4+juI81DO1gm7l0r/Tj0dVBTBy/NZkGNGmjSS4wVEllIepnzmpexnu64UcU9DlB9Cz4BRu
fmokaOAo6ZDkw9vbxxOYIqbjW+jazOecFTFLot1EYAFnF9djXNSCmjtwAEWHYN6pPslfnhA5dt11
ZAtVqCRcDHtDp+Pu3MvvcDtlc85v39eKlCruWakeVmJekFvJC9tByfMT4v0gK6xnQFkJroSeD9W6
wjh9S280knsmksutKAeUUushuern1FhlpdP1XtJO/jbrLaQpBlcbqhDCFmrMT8LwTrK7BSGGgxdJ
z+aP9i5AB0RdtkDOuMQ121BFg3TSdJ8Q2A5FrHY6RESloB1GqXULtYrhx543MIOX4Baa8SI63U+O
OiDolQnhMag5vazFNv15KTlsDABXQ6opoz0FoYLhJ1NUamlsfBxRPuSofH8abqRPetUYbMuW/04T
mM4sKag9Onu5UVlwJo/MxbLQ3t9AN+4qHSWGxJuGyjK6FK5EZyhI7DF5c9ij/Hap4Y8uUJcf6aOQ
T4IDCsB6YCsoGBM90s4JWKGd6mrKH9/C1XsXUy7+WF3bniZP/oUTZ9Xprdjcyt5EQJwKdOnPwLni
KOYCaNGYMgTX+b7HxGlQQLmF5xSf8o/Ti9GCON1mYlwGbCtWmIoM9mtlD96m/N/NfBBMQxaLVz4p
ulD/fZY49jswSpWPu9+JXrYh6FQNU978Yj6my3paIEvQJZzY4XL1d1E+p6KWkDhQrl6CF8DICuYn
hW4vdnxpuwpHIhYs+yUXQDe8DkJQdEdXOCLA1iFze/+tEpVMgkzu3VdwgHgd28sGo236zqH6PVMP
HwMGGe28hqSCTnLN+/GY482STSgOKnDWW+ZpSH/Y1VuB52ZzHO+XL3ZTOSyxLOBozyhw/jJJtRWY
x6UeT6+ZUqdyY/AOp+u5Pc/DlAepO4385Q19zI8jziWojB1gE3n6qZWW6VDvICrozaXD7DyOSoun
69El8KKRI4KG8rtrQj3S0ccHbU3CUw0DFvVsZi0TNhxK3lARWDetL6Myf45T2HUNLA5kaX2gHncd
VSgP4KW6yJj8pTF1VohUjHBuE/3Gv1h72Ffl90mdCH7K479QmD7gf40X6gL03+wZtTutGkKde87p
ePQDNIuI62Ri7e7xvZG9MaFgd31BJ4+yRyReYJzDh4luL5eif+L17HMiyHAuBIDsMlwE6GwBo3kA
iZub7VEJJWJjnwf8oVe7GequKMgATyaEGHe9bjowp9imf0uXjrESR6hPV2qKPnTwkBobyOc4XMxw
yf3a4o4TF027OhC5U7HS2C7gXEQJk8rlnvyfMQLw/OBd9K3FD+8C+BWZD3ys4C+IWqCweCL8ULWy
RdCqMO+cIOMdN4BfNnrQVr93fXF3Y6zNk8dqa1cUytGq5YhSn59ZdSu5OcgFMtxzVGV3BZYYwnWX
lRP8Tn5UHRBl+ZSXskjlUSy7k1mvOC3mDWEWRpZglPfuC+9NTIP1MyPxIxD1oUEEoLPEqPTdVe9D
HZuzS5p+6kMWcghLeJPropqQJf8AyZTQgZrwwPjbGQeL139+1DWFg5pFZCWHXNcILgWvp1TveUeg
HYinimhiIb9cZiPQPkKIUzDGzPQdilFnVMDRmDzAE12mp/8kaMrRBUMfFPPb842Krb+2EXkVsVsI
YIFaYjeioZTRHuNL7SNOqs9HkNdrfOUjGex0JlOVNkH1uOywxQGyG9DJg2/FChe6Vc8yqsRPfVgx
fec5mNtbiMUAoIMgrvrSEBQmvjbPS+KdfdGXFimCMXPUmReXUqqJXFbtLlXcG2s/RrQhPFx7t6s9
5cNJdxQ/G0fmR5OzMDwCo5fsFbSpT7+/BLRZQT5IALlt4Cs1uOoyQpc9OBXe1Y7DiVzb6Zy5YGd9
L+Zel7Ton4iIu23tsrTZrPIVMfydFjXFsrshqygruw5ApLcXArnvdjxVNAw2hxHpTgxtS6fjoOfn
IFANXBdHYoA4U+wRU4LiZyXotOVlcIugaQoWlP37yBah4nqlyFiZKuUDy1Qmsf60eWG3qKwa0NeG
iihjKzMwwyYdPuuMhIbB0BGEjKD5fN/58Mx1g6ZtGZFhQJTgJFAs0Iw7EA6BrEszY+mqWuglwoCE
xu6INhyevdkr3mb4dw8QsaKdIPGn7lI05hJhwlXg1XJjGiIaTXDcpux4t7r61JxAyFUphC8D/XEe
DhV9YulqvAFet3bvzoAmdKba93TJT/neRmI2hygcXasR173+H4xcqmT3XG327MSqdYU3pUmKppyI
jyjPZjAqgvT6CPEv+NUOs6KC641ZLM6rCWwp0gSkWdie74VOWtqmfmaKzLL+jpm9/JbW67Z9tqDn
f4L+V4WOWVcwpZ5gT5PdX96AtXNps9CtVP7E4yZytjeR4c7rY7sJBZtQk1wfIOg7CFEdHP4OGQnI
W42immSY3RG1RrxHRmo/r+bRj3H5dVDMsp1q07wmXKHOO3Xw34fCLkhfEzWCrgBbsQL+13Y8hZPk
SlzYIHMD/zoyKjSoXL+/bmkOXZHXv5y8Pva48YVHKyCnyNAINjBqsc5//mgyE/7bSDxrDNLhm0mQ
0H1KL+iiWwYnP0xsnjycjieHTgSwGzWfzEWVPQbK4zAWW+6wQEJWTgKSaWWTT10Dj2LEP4iE7J2b
HKvvaKRROFl5jU6ifX/Y06y22xuPJ/uiGNzOOsyulFYYqFLvuaAPRDUINchTj1JjjTa5O3r2ivxx
V0FWjC42SiYobQNMRH1FimzrG+ByweYBY0JYWdxmaM4EY0YfEv9bFnXE7Ui0llEoyXqxbP8N6MZi
Ng1PwA6J94bdbSi2s8YnXlo96YAuHR9LfqTPf9PK4KRhXTAqqUyva2MSe9EgS5RCexwZKBz4MJwU
Fq7Po93SrCG5Ciq4Ct1NHTyZyh7IdWuvv5rvhQeOu0ltxJhIjegT8rrJ3Ja7EY5Zv4+XHzZBjzgq
pZVE1WxPrwnK4h4eLoPxjj83l48hf0SF0ZNmiXL7QR8ipoJwwsChjg3+ciDtVnFQDrcaxteOChzF
aDkOlYyRMAQT7gQTjhXG+APzRQHXh6jKs0XwPZl/y8OWjjL/vfffUpKnfPgDPFj1IWL74u2O1iTp
jt0Nj7XOcsh3DohJ2qpRr07BOVa5BIS3uqKM9xSL8jvdh4HjABsTWctpDx1S1RUWnJ0+8P9Bw9i9
NKgqIvlfYCzb+D62nO4f42PJefwd1jIbXRA3wUPrmcCo9IwdeFeA1BA/zjxbe+BPF18x7svy0mUg
+lWmaChXexJ2K77ElaFicLkGwOGJLtoEhS1BUGb+BPsCPzeQ7jIydJSqdahQMQAPSPTtzwYmIniT
4q6PR2rHbsWSYrbUEUJ5MIkDPdUDeWR6tCGmgqTKveMw+T2D9ppAw1F0FLpFpAU1X1So3noxQrXa
yMOvdud2ce5NGDwrtjdtmr+JACqHMhnufhfnxOHxhIAeo33fWI4B69jbX8ATYO07hoPo7g8cu6yZ
aluvv1N60NKpQDp/99n3G1bccANrcRqYtDgliaPY8YN+/OknB4gtxxRd/oWyeX1r9VoDmkMvmx0B
oEKEWCjkn4HC3h6M/H2mKzzxQMLDcjyxD4TweWQs5fB6hHsAlEgJPHNT/BMNdZN7NT3AR3r91WwV
pBqr9Q3fXeI4+ja5YcUE+gfqXDkoXrKKf0T7jcWBJ1GV2RcfaqUcxsO+FWBqbdlwhAiorK6OOQL6
jZKP1jjD4+ygv+VNlokVJw52GSg38U/wVZSs5gsjKR8x5XwjNoo/488TNjKrl/ueppZ7rRaryduv
ZLbw6izz7swUbn+VDiM25eaCJCBFTzf2Z0QsusBhCgycQjhldD2Tz2e6Nv/ElHv/tMsPbBNgPeDI
E1OrIKCzy2LMONDjFnCShvp3EJ49LbYeMnqLAIJwrYTV3lPckkaQ5uGMiFQM3dwybvbvxwr5iAB5
TEkBCp3KRkIj9zQbbEnZ6thGkDfKIUCj7T6qC8ZKq6E9nLAM9PVZdP7wlRp5WA5RrDf0pTZEpjMY
KBEfBLD8YuEPXB96if93Tdf2zKsqvTf7aeA+LmMKGQsspxGAyT6sJ/2Ad9WqBYXiLK9gjQjDU5mG
NN2v6hCn+vo0XMhWzqL1uc35wDhj94vtFDOhUOheLNcAwFWQ+PHAPBjzUf14oGh/t0cPCGMmZ+Ou
NvnfPmPwBJKZaOtWpqVSTeMxlURwbylK/tt3tGQbfsvnEBPSaIdbmR2IqAN/LqLR+Ba8hqGydgxx
jbmjnlwLeyORnCk1xZoto1AInYm3D1wcS4ligo2wAjQOLm1k8Jwft2W1R9t8piVJo5h6nNVan8ZF
LhBesBjL2MrjWSBrIfVPWPMK5k10WPxzNeUzt3ZWnDbeRnOUkxv9hZd5kGLQFP0o0www2PCifiJh
C3GjMWXq5Ti97DS1qhwbwipmMT8qVd6eYUOG4+4N3Fs1qa1gL62fpO6VfASZ+Cwyh+DOn9zRZif/
JRWfQXBxes4XySpEmeycat4/pu8j4AiWTw50HYNx08YaaUqTOQaDM1MlMyQ3jBx9kp7WpQT+3fsM
Nkeo3EaFH5rfnHdS3L923cxwBBkOkAZiF9SbG0SqGXWtMZpBjZhS1f/qy8ApwkYpYnlo7X9GySZb
LyDaiwOyWRmJ7tKiWh4zf9Ki5RZ22tIO2h1kkdN1Ch1o+ygMkuBySGLIJI8Ed+30jWDXrVmFXmZj
E4F33EHOSN6IclprI49jcvFnmXsaXX/OxF/f+LRx+OZaelkF35BbhlslmnDCyav3wkG62G0mTTPd
e0md1YLVvmrbSeCd19G3UUakiurhBz/dTAorjn7waSKixPDELNJWzSoV91MBoBHBHIvGEJM7PpnL
X2wzWE9ROMz8LSyytVOIeacbPfvYW3r40jXAV46l7JF/wcGTsKxQFSPV41lYjeV3XJirtid94HnP
dJLp8sIxB/+ijwdm1dVaKPznPhAscv/dr3Ug7b7oI3ykjc4JsKqwNCqEboc1rZagdhY1bZh3bnG5
qtQfCxauJ9/HmWxmTkLQRCT3ojwgS7fZhmRCKVa2blKNHOWyUjP3txHsCmYkekHM+vOeZ8XELqOB
zhVtlXqWbw8o0aIjboEMqYKa6xuNhD4uFRJIT9CPy63VHFmWwr0hmn2WZ8ed2xjoUrwyJtTmyG3Q
vBGWhgc6BqTRt8XqL8Qig/o1yx0yzPslwSJxb3ETfSXjFVV77Mm4hwL5+ulqqPm79D+T59G0/AxD
y0ZHtcxI/8VES4ff55ByAo8JE/22jAdl3ZfpW90kQAFAICJi2vEOMdAiXa7bQGMeFQtVwAAi13df
SNrmLDt8KR5DA2mR0HmqkEdWtLVbnHV498jiaacDSLeXI5k9h3V9KvlmVJ16zQMZEg9pk/o9wuNl
E+wBnFH6U/0ZoPWR0Z4HS+sRnxW58rPOfRGOFQ1XZjvooTVzA7klYDWDLLn4jVYgdN8zWYKHvs4j
lFqy8sRyFePMjBHae2yzux4u7Aywuec140dRIM5PkXfWnCqiu9/k5cYuUL9cKhhy/dDqgslvaYvo
sFZOZ31bHmojFfRsQYJZjEPtGr8lH8+9iKs16B4hREb1Q2XzYXClI8NJGmlqIAmPDE3RJo/FtvuC
or0eC/I9BVgTbzQHtocSbpO9SDxhk5IEHPTraXm+HJ37Q8dpxTRZWI7Hm/BuyiHRp925q6djsfJt
+/tdanM3bTyi+oz8CqZh9VuCT3nppSx7SCcexCSggPAkpi64EZ/CCJXTr8g1ui94vuIwseAvYJws
8lsJqBhjWPQm724322y4D6KBrLo0EVsdWILzOC1QUxs2nbz3eD3TpbFizOOaMnjV9PXrBlQkgBIZ
Btu32B2/J9KohCWo3kdm5r9XafKKwWePXW7EPcIb3Cn/RQj5xSqzvdbX3X3OaDvAKvfH9wYj6Jou
cQ13h0J20Zn7b5XiMmFj7E0OFAQH66HV2oEKmbPflW3UCXR9xUOkdm0knVDacDpQNnAl+uXrADZN
JevOoTwFFlz47B34z5s/sJUJ1cq22aMlbgUwbtYz7LHqCBXyP2cTA66cdkeGNdmni882FIx8FwkL
ybX2xOpRB2eFTe2t7gfmyoobT1WglxpuDiYpuYxIXu/OWvgu9IkAGtpriPHJF2a1g8JheMAjmYTH
n7jvmHqh12nrbqj44Ckz+BFmvSqijFF9yfErsK+vZ5RsiFam8Frg31oYW6sjfsRavS0dLdvOLBDU
jcV1u9bHq40HjIeNw+eBdsEMGSUOWyDg3o+2gZrhh/vWJWhrtF0nWjJBpKk0saqgFIH6PaaMIxxb
cZ8RxicaoQapGf9lyTgERKpmBU2TQoI3ft6BJTbR6OxYsPgj50z0mQhBs0mQVmyrTzLc4xJLHVfC
aHx1KjGtSwVI0L97vL0RD2RYOSDcxZxQkRG2y77enPATNXRu3WWGTH29SLyr1lUSEFbP3O6nFvKT
a2olvPhXwa1iZSCuCoRebPs4/30peJdr4MKPievZwGP9x5tz7GYrheI+EBsSxNmRJHRLvzlQ9tHM
kE1izeB+hSezQoyTGSDzQYoabt2cSLEpEFf1f1PvNCi+OGhJV82Vw1Djd7G/zD83i4YvdTe6zACI
Uo8QaTdPPJZPvYzChxtaToCMMLdYs4/pHN8HOnZL+/j6dVPKtczd/L6JlTPDJDotCx5mYMQZmv96
hr2GyZntBcR/xUvE0xvpd5pQ9xL7fp96mpl9UBYe6A/n/zI2iRgYUFqiioQCsEHfDHqTCU6hwGYv
oyMsp3u6WHDV5GEO1bBEyOEPlTbbexh/HdqqyECHCDx3doIMSs6D56+14E6joykduiGDM4bJXbWb
iISNR1XlnKj9gKua+zBTDMT09v0et9fX9EvA+Fl6gR3C47I9Cwsd8O3iOQAGxfyD8srYOh0ku6NW
EOxCf6CgvZRXJdHUz7HTxVG8RZjpBTopdM1ELIXQ6mjcQBEd1y2YJASOMFSCon3UT/xpgmSc+poo
/T/APbd0ftKSggXA6x8v7numLeNuuL2Jm3fg5kzOHtZHKqn5hTyELF7MsvCHoI6ID4S8XG1eKgEX
ajsgVVs8JvLfKU2bXIow7YaD5wQ99hC2nkaWkeKpnhD/W6+W2ta0bG1cwhojqQ9xGjZYQPtSn5nw
8jLbDDeQGMZI+xPChmp8paTGira5/8QSHnNnGnHzNguk6Rf26RRi8AUPgjytfSPPS6J/CGYRVuc8
qfYed/kC6o2bUA5yon/MB1KctIb2ZH029wkgQaxyrP/sVQXMT43mrqFh67grd4+/AanwxL3iDEPJ
ZRc9oxq3q27TuqTlUSjFgLuJlSnWxDBdXXZ1EXhxHGEdScYnfvv1kwP3UsHEtt2s20s1/JoeaeKm
STPDNJ7bTOjehS7Da6hHLq1/7Tibv+jAci4HE7m1V2ZkPxuYzNz85JCNi2LWuOBTs7I+gHxurk84
ofZOZgYXbpiVYv6TZJH7UexMIUfii4BkW1bPRQo5q094nvwBOq2jww9uKbCpm9WbtqZgEjcX3eTE
gtu7JKqxxkQsJRrcWhZmLRKptb3cz7nxSOMJTlGSQ8ETMxFNVrvoy0sJGg+nYBjRnCFJG0qd9iKM
lFCHwBVhhgJ+0yEeBfEzzN8179ZgZaanHMTV4zrYL9L73ZJhwt7hK9T4WOj2Vp9eEJgcEVvimu5E
r7ZD2fhKY0cfPxRJjCArOQKMru8LY2GSegHqNkdvSxBqMk6M9cP7E0WLIQaq5VCIexry5K5HqTAg
0Bsrd0p7YAeOy+SkM+QIsxysmHknf0Ze6G7B21ztmLKhoxsodzLUcEPxNRlgG0/JGDG/lenbJUjx
Sb6R3KkZTZsUNVUGnNXecr9fGnZ4BkOXlp5UX8AhTotEUrZUIz1Use0DbqIWxX5ieJEytQurzuFb
7s2Jw3Qshpgv6o7NsW0HP6yCCt8qcmLd6q5mCQRoY1iC6RovFys0QFKFIVSoPKkb+EQ4NLYBOMSO
1mOiF+la5P1YEcMWXDgS3XZINln8HJ69Vqyg8z5IyMRNvTrTxjY2Zj9psXKQtkVovf1MRDFlS2c7
TZ36pCwJtS/r/48sM/UrKBSsdW8SITXEyZqstqEddy/BgDyC4PSp7ilwVMCCZ0S5J8xoUwb1ifb5
6pT7teLD9H4Eypam61I2eOSBxn+/k2cGu4JZC6e/KdnURh2YN3/omEiw0BZggEMHciE7PKq2YS5r
w2gTBEIh79f1pxqhE3RR7KDO949S93P8ED4AJCNW/5AJ36PPafRmw1+sYElTKju+JkTH8ort3PwV
mDVCl4Dp8VgRaXj7YyQfc1rN3WA+JisAXmW0gjmFdXxijdBe7ILz2cVPrCIKjpxsKdLihnA9thsW
LuTKsp8IEc5U0ECuxEnIa6z238d7QrDbhixk0KxF2PrZ7BLHpUpir/eVxRI7WFV30Ue0k6aqgwz5
ykKB0qY6cZ9Un8QKx+CmjL0WgINJIbzJ5BuJzxtNDUlVSdPWSc2bY/OK/GsSAOcILLEX1IcgQJk7
4TJe5HReC/oaAYOkhmSNqd+Tw4fCOIMYvsnb28q8/r4FoFSr2djUarhzLes6L9+L0NSaOvVefQLN
pRoIaWaFYJgLrhiYwz2aLo4wcyQc+G+80G3ZbJx1uukDkyZqMyz67EkcFY3zcwEyHoS1o+X9P0oG
GHnedUu784+/2B/xCk8/alvnwJjPmRNWE2yu0pyn1x0HehsDtT+lSVgUrzNVtzVmZg15FtiyN0B8
9aBLSMtKPlPAM1uQbm+A3NakYHiJy/9ECBodvB/nT/DIqjK8Y5av4RtLq5X2OJlFLtIVWicDNuW6
SDW7VrfW4xYu4Ooo/tp0tqTqC7lneJVzP26MieI9o3eEihnJQ2XijuV+ThMnkc3bEJgaKyb8T9XM
QivmYmcD9hMPrU9CdFRAM8//0CA11cDSc5WUOVpZtLrPjLdCzj+CbFNG38xFNDasImMm8K5vMNjt
F/+BzY9CJBX6HA5CgWbcwVMv82jYRX4cueMUSnk2BWX198VCuhX8F1mU3rMALTaszTR5r31E0fyN
aIk+t1ZnsjAlvTyMdmzcmDOGnx0Z6ynU7lAKH06ssIpwvBLaNu8GcvPCXf5PdNFjS+o/ceaciRtn
bo8lOW9Z7IQ8C5j2InHaJ/Mj7QJ8IOzAP8VGNgdABtxIxG4kwfCOPnTsIsjs9//ZRhrS7H0uu7Cp
tnQrGPiB/ovfxx2j+W9uDjah4g3H7V+VdnCGgkZnv7251Jqco+TNchOlV/clpNXxIUvRXZAjY8Dj
00JAJB3iD9OCBn2NsABovbwCsRgOgP3G4KTV/8s9UjzOUMlxEb8DkQq50Hb6QgHbd21FDVirQXLm
/ii48t8OQ4fnH6gnbAtkOzoUgPI8A72fZbDRPOLIyzOGTxbDu9lXUdzwVnslF6CUskkbvzVUOSUm
U9Lg2oG9RPDYxx/fHhV+2qhf0EWPmtZXmb0gyu42l1OVdVlJxnDGKHBnJE/SbUyRN8FO3ASWq/ud
X0onh1qFZsiAfvuP7MaoHsC167Ycz6Qu/xVtZbjUTIxjve3sE2Vl2udgevPk8IGg4ihKIz22YzNE
hKbiD9ZlFyYQAxjuNN8zoAjc8Vpy0EtrvLdJ1Na8r9fa8A71QGqegCTQoTMnQCRUuBrk/0vLO5x0
3Qrrm5Tlhyy3NiuapyLOYgWfeghLMAXRldc1ySBzX1PuUxJFBQ0E0DYHDd5RGzS542cguy25mqIQ
3Xyz5izeXFGB7NmW8mm8laa/YWKR9R8PeeWh3qBqEUli4TjacvRNAldtp9mekxL2ZiloTE8sAoYp
ZuzJuyguzCuVuTgNg6CVHzf2M/Eh8lOhKA4cGaJsdm4TBaVpx0k8qM2EqyIQFuwq55OrkxW5/HJd
7+YsFv6EBqIeweaOehuuFZcHihBimZIBu03KsVaKix9TQastBD1BHnBTOBsA6dpgGNoNvNiKxiAj
+/t0+q4xuOqJJoaSwLmAo738rPRkGu8u7Rs29s20EJHYOOljXmItoZ9HU3HbpUxxF6JK1Vb7rgzG
3NtMuiFGGjimT6z1u000v4ZfKdiKlYFf4wH9kp1l5Ly3DoR045/skHMOllvRs/7VtYV0JBqXE12K
mAIgugbdkNNkaKRrHjd4/b5q0aZSGGNX2Dy1iXS69lAukvJU8wbzzDVGB4a1EUHnovXh0EFAFSCE
AsoCcFiZ3HY1JJn/CsvgAI6PTeiEbcnJCj3m3QLNtVC68h6RUrY/Od6Y+Wv/rjwY1aumNly4LpSD
eIsJHTdB2WNOB/hLNxYbhAPP1oV1dhv+Ea7OaknVZnQBNiuorUESt+8FzgRNbVwGJsQB2z8c28WU
VXH7r3/EqjhWD0iDgrn/V94+NDA+9TuLcNE1e6JUBcrzEa4HvEaSvK1tOA8FGGJxadhGRgsYZu3T
Y0Ele+VHarkN1IMydVvsuPgGHMMbGfWHpxB6eO0DwAt7IX9WZW7/x8Mk0op66hTXJ4aHoVmA/Q15
i5nVw/yvLnl1K7Jwx6lPCyRWfKzKkTbf/GnWzhMwnmpJiFaHZDumhYLGCa5WswZso+58dNV8ZU0R
nrm7UlhKMGnY4qHpNOOhiLCIbV2+Gw+kcz3euucK3ckBc3IHz3Tazg1YW/r+fjY8kP0FFKObaNgb
bhKfXkBW1ZUQiIM20/aWO3dQTrITFlJOXiHAJH40Uw59q0vo8YTHHtM6FNVPKLuiLow6HS5NELlt
U6lPwDSUTtIErEEC4CVnX04dIHNn2hbWMIhqvX6fopvRpNaLmcsroqmJnVliCn1RPGlPixqTJmlK
Wh4+Axk3CEA4IARhO+sx2jX79xPEI8f1W6N8AOfsSmMhzKFjJ38oHfroBVFs6ompD4EMZjEuem+u
22EI+AkZup9hrjY87+2zFQLXd5oLVm0Y82njSW/xfwkwMisPqgx0cjYIFFnz6Z6hdOli+jsv6B3N
+JLV3GFWFy+/jhzOc0nGG+gi3ixGyFvnt5jFQyjoumu4vZDJ5kixYourZH02aPV3GiY0kwnv0ghY
/bE/kVgp1OhI5qIhnX3+VV2KR+//tH//ZQgplpvAfGZ9U4+SvdjjWD+VsquXsoFST8BXDXBQDCkW
g5eJSCxmzR6AsUZJ8f45L8bZwrkTWTC5RIci69AML0610PRbKLJMujXubKjzR+CevHukkQKq8tgz
YZzLu0eeT8V3ebyIFc3FwedQXSdmja0rYvDI1oYfbQDpAxUjczmCpqHyoACcm3JO+JGnMrt8N6ta
xGKDQ/+GABrPliwA1k7SHQywhSUbBuQY78JeCeRTrDcdHx4wi5Yk1KL/DII9kPxJvcGNueP2ekgO
d8S1Yu/pEPQRQfOznBPpzxKtXe6jvcb9Ug7ya8CklEaYvOPctrLg3dE66Eh4x/yns/eI5Yw4CQaK
59rFs/YeEbc2Z9dM4m9OHfk94ZsfQ/3resVKBYwxvN7KdEZqWym+p2IYIETz+vgqojVU3/FkjwMA
O3w851gRZ1/Jp3NCuBLQHO5Aofl1NxXJeOEYf0I/ALyZBYKG+IsWVCqtz25hNT7T61hjxhA5e/sm
p9Wr0V1cHsM/FAJR3vIizUMqWUfNlE+TkBmGeoEK/CziHnKW7qOEKWrX15Wj1VNJo3YuVw+bmPzB
7VIK8G9aD8D8zDMJU1LfJ0kfzmj7C4QHKnrmTFNpRWcNrlFMAmU8zvAOcai8NKFACZm3rXn85E/C
IOiSRjiMoCwvEMMnytWXdEp4qaxTYpKEp98wmdGkoFiACiGEGGtMmy4I/BJa+8xfLTEjsslHNhvA
09LJksszK0BVnj6afz4/TkjLM9MsasmE0IdGEd7uq7azRsjjSrOmk7z6JwOl9Bfd4sfQQtqd58ZO
8wIwQRtStilHRzImBEPDHdw3Uuw0OfTovIeQXoSPNy52DZn5d0xY7hg9FdEolp6KPtMtFcaOONAR
Vcy0/O5D4ajiTAQcjLBm7FE/1T0NjxWY6/oPhWuVoumK5OZfXNhiaoAADjkbJ+82TRT7vRnJhAp2
ZJ0WtmMxyuxW6bTQlS7IYa9e3qNqe4wE/G4owNMSr6fTjfpRYygHVNy8OGkSqySCx4OhgsKvjZrS
XUmfTxsPkODRNMZbCgY1qHsgPxBHwafOmeg4prvhdTvs5xzK5R8dvWOw+a+0FJaRIOaOQ6y2vqyK
o6ykEO6eqhcADNI8Z64Vmi6rbZfth/e1RCyCClJ6TK40UacPdltAqcghU0OHEVOZmoMF7JmqVgFm
fT+LlMN7Soe+V65AgO+97iE9nvmu8PEWdwrzZh8tWIVsmgVJEmPvAoJszDt6CUdyZpGBVaLDu852
D9u6FOBNlu1GENXutOz1AcwxN4S5StB2TUzf/jiS6DwjPJEHQIi5LetFSUkXTgMMO+elzj1Ks0tR
ObwhNDjWS2Pe+QZq8HZ2WHfCviPo59lCdCaJ1J4mT0bSyTvLTOIWeOCyahFK0wiiVHyp8L95VqRj
0w5MjNXEC3mwXNP7YepnmfBWsy7wEaOo4WFQ7vNb8CEHq9RIWLIBNh7rXQnfXgmw50odRcrQm44x
ATNJhfLtiPdiJrXCy9WoG0Gh7jVFBKmG8GM8muRk//BMzEO9KfPQMyUpR4cGwb6YkDAJiPB1qpgH
EE9Iu05ojWPWc5aVKdhwa1VCdFt7Azf6EW7DWdsuTLdcg+Ns3RdmFqEzCdBQwXZrW3VQ79v/lajU
UpLyKT9gGxGgf7KMWcf2lECvHm+7Lp5B8641MPPZ3iSp4Upi2jS1g3L8jNpbJc31hi4hUaSUR8UZ
HmREsRtr01vxTto92omChwzyDx/sh+NmSqU991gGeZG0uvzF8RtZf4gM5oeyYJERdUAw3Kb7aQUk
XSg4lJ49xUAhr9nOuqyR+SHDpQwnIlf3jZAo5cVWWMrh2hBWpZ+mqCLcc9wsCyG03vD4UZpDe0V1
BFKkTXJAOzTBpy/DDozkwximsjHgto2caU4c7pdCRahiRZtdfSlFk8Rcf49QJwpBGA7wjdz2AKVA
UbWl1ocVUHFcKfEV1NQwrVMEWHAMB0jerOS7E4t1NIEkuiuXt8mcQrSRMJvwSW/ZzbnPkj+7HwYx
mOJ/lT+fjeZHBdSakoJFs05XQU6fD9xZwd3jDnzWaF8gQDpY7w77DSlUvKAczB7oIwTLtjpwV4rF
X2IRIlbHK5BQWSovXHCVSYtsMJIwwCnw3Xmy4hezaBu11XALTkEdWVmtUBYC9RCkwEB4KYFrvLyK
X3QstazsOY20/VbWxKX8aCBHCt3DSJu5DOj7fskbALiIKk06umwQuSah7kG+n2NDQt1K+cn7On+K
0rmS3ylL378QY4x6SAuNdrzwHXenPQmyJg6PF/0kCdpqMiJDZXibaRhO5NUn07kzZyBZ7T9bzsw0
u4v5d7kQhXlwsw5V8KJ6Q27dPPCU94zw6eVLvIx8477+mjAgrhofUUWhcLWlMCPWlBL9SVp8Dnad
iWh23OzElRAojO9WXZRc44vqBSeOgNkuMoX5h3bZWVuVdk3X7Y4z4gdDKOzfQH/3B7Vf8MdziW9T
3s9+gdt4z2yrIvIshdgx0tUwX0aHq6z214D0BzU2GfeRailrF5EfdCEwZOL3jUf1JJ7F6J8FzRM4
nanC0JSF5PwJh6GRikI2folzBDnpV8rdcn0xx+b6kNI9cQAsh2C0vFCOUamUOyf7673LEs66wtOe
Vxkd2FvlK8CCQHtzQ14OTOz5j37klDV2poC7uBB7q+jvxp2fta67iNq2uno7P6T3p+UA+n6+ez4h
47jM1x+l78gMpCQQuTwIwPEvrtrXnBK3Vc0NOJrpiAxB7ErslCls19H7teIrk1Q++d64YpQzaleA
5fNr9S7ZAfjaC5qa1TSJZIwSxSE5vVqREWTo5asK6uH+LSwidH4VsN+D3Iw1lmy8d05GviMjc3q9
Al1MB3KVaGB0+iqqyj3E9uavjGDX9kXmCPcB2gXNr6TXLwsk7mhA1I3qg6nEhpxD9tdx6mXegDtJ
GJGHGY4DA1MuVCrigMtdUru5ITVcF3WLmGDZBY4jmh0FRhrOIDlSJN6jJugnTLMgZp+bfMhazrZB
TWxJ1og1hz6F0uWR1R4UlssN6Gf09gHD/3Dr3xBP6c/jsh283/X7gSnHDUGhy4rkdk2CrxmpUj2R
mnjQeghnJDBycSGaZYE6dvtxWao+ls0feGfzcQiKSHFHtxlVEyY71SHO11UcXh0+/J6dWN9QLazd
3UOf3NeSB+nAGQ0tcJ2ap5I+69rD/w8VWrTSUs478lg9wvaMtMB8dQl7KBbUBMj3Ct3uxIRGY3+7
5qcUi7M6ukhMe0KaIMj5PMkGH5N+6C74zcZC2fAG3ZbmZ2u47WAYfvgIIXtqFSpnJpRZeuNlseCw
bsd/CQoAe9qdk/HjJjY8SYXs+WJ9ZxWfLWY0eR1asfz85L5Dl3oGrxQ3fMmtJ+F17bw6MARPqSSN
r6KU9uPfh2OKWrzozdVmn2+gojJZILa0hAPyOs3DAsoqIW3a8ctogJOdcU2XgYoaFO52M4sz02aY
NRncNQNORLWyAX7w8p0XBfGbCzLJKmtFTRB7kc2waX/8+FB70qv4VLjCtv5TUr4YjOxscf+sw47q
bEo95/HK+FYKzTBjXuIEM2OKP7+KAADwlbSimNDWi+aViCTTA5FJ+1jWKBF6xHRpqQDgcxrGH20b
fkMh29BkhH0eLLEeL5GAfK4HtyPSxF199HsG3jNsG1RuKJtIsMIE4REWjksH9LZHltRzooNhdeCH
F3K5N7hnzHUUUXoJRDcvqTuZpsm09Gc/C4HXUA7lV16DVH8kqKUO0o/yF9p91KxpMDhsKfSRbvgV
HCd9G+JjHhMbq6YVmgdYst4b1K1FZlb4pNbcoHmhGA0C00sHQfgVHQH7FZflWCNwU4/BBNIklMHy
DjMZ3GNkDDAoS5yxqGGFVpIuKs9HOkj+iLQ3Rg6PlZbYF0AlNpo8NJnsBx87nkAbqD3sm0aKGz4I
B11DrOc8VEIxAwfXrOXmJlNNRL2wCdUwUK1V+9c1AaNhQRxCHCfNkF74qWVGV250VLtBEyBpMJk+
LPRB2/eqmNYSZ9+6F8fMw/UxXV/7PE8YxTbeG8YXSYnotbFi4S8N3bDskhICHYGZoDaT7LYbLPim
CXt1xF3nQgwFqbdgP8EmBC10lBo5flMBIM4jL0EZ4Fkmxf+xYeA2cPXXid/Awa4CdF9yHo1fknNT
suvkx1nxit/tU3UeVKS+Mlf234T9DbIF1A5pOnv7R7LAwgzNjyfG1pIkwkKdU1oP3HhLJ4e5c3AL
uhCUZIHXCjySttwAhYmQbjsulzRZryzs/0asXdulhg/60s226JHeCgP2rtgS9drEADRIKzcPbJcR
WAD5EgIegZPfpksGbFC00sKBTP04mgl1s9sERhCj6r/It1ITQ8lME5tJJNb7JvRz6gTHb1wVHZ/e
KtQHXHA61Bc05r1uZCZl10P9r9UQV6e5zabgjNK1qPrB3nNOp0weSN65CSToMvD0QF6KRLff6rqH
2XmR05EuI8sZztvo15rf70xobePl4r35dlS0zM+5HN+fG2JrizpezG5uSs9i8MlLNFeduQRLA7/M
R5GwuR56ZB6KCeZB75iAgNU07Qu6hNUctLWH576rxOtK2zfPMMSBg/oXwlV525fFo6EuUfqMNhg2
HA2KnsQNZfkBfaQ6AT6SYcUpVQn5ET+le4PrRH2oswTyNimgzGn0LKSFj4p3UbzyuEsDH/eVTYTz
iSUAwhAiMvmcAViSg20syIyfykkor7nVjAxIT+5/A8irgX6k7+T+Zqqx6SIFnTcMDenAi12Dz+9w
YGSOuqAUR3IIM9tj8wEoB6iL7jbXKZR4A+i4c8ERT9JRyp7cFkumA+BmQDR2y2/jPK0shKg/v2g1
PbnWINAkM0ZiD9YqUcnaesZ4bK1J26+FuRIaHrXPz6pfa3oG2lLkZk1egHuU0TgmxCudXLey3B9c
CjVuPnt7zrhB2fQ0N4EEdxdv7Xrzy8VCj0kNIq+L1Jju+Zx3+W6nBaAqokG5CCMwattPMl4xSmfG
tPPPFommGHDdLkfgUmXH5xvdH78S6F8voaCv4iHLF4BMnP8RqD690CIB1TXcQXMSztH0GY2S027J
8t+5oSk0vYo2qFfOTyrwQKDjuaFsYsfUmw9BMx6wmJsVLTJjFVdUZ7U/WqUS1zuymX0z5akpMsge
SPA6Wd51iVw44cGH2sKIjnk0BD9cWxjBTR/4YPCt5Q6Oj/lNjtzGbnUw9kJMyWy0p0PQGtzwvTzF
PaMfS9LzQWiOeLM9qwT+LS8CWjCTtHYqTHYULyHTMyEEJXlDvBR4FL2DHM8toHOcCbSveTwhfNS1
xq1JytUJrYomIEmZcukbgWp14DeIUtpUlXqE4uT/UiDOQo+c4nr+2EP+F2wTeA3LqWD0J2ujeIMW
6dKu5fLTEFVdNsiF1/AWwJWK7t65v1H0OLh2ZkMhPeJvEMXMxLFHxfYVTI15AdMDy835fa8v79mj
K6LD6oZDkkBhPcEYGYklwBI5eqBypRQ7r/RlhtOI1qzADMOJxswZlqz6bvcpBkUu27gWlgMCW4os
fYWmSop+MwoH/tii9Xz1sP+wB2gOsNt3l4I2ttqi6wNShywy3keq5d2dynC3f5rkArf7ovr6swCP
j9f4qwRIkxFBE7NGhcoL44J0DEzhza1kvYZhVsk+h9uDLSGvaxKx1VutlWz6AE9xaeq7/gDMyYpt
oMbh5c7AvBpYIntoRiuDelN+utXlE3U83NZhuHrn1UrWKh4eBq77FmyT5oPRnGiqfmF4btLNiH0F
YYNqkYfM8iVDoDPKG1CkXiw5w5V9afWk/8lMsImcrrTyUKfcUEFAdyT3bHsl1uqkkycFFLnKtjQi
d+MRVjiZyv+UsKNXLuNH5XvVM3hfJUv5lCYKKDwEWxw7KzgqRHEimSKMwEFSVCA8IpxYrYQuJxNs
N/BrvaucZnc/dI9UlQhzbvNvzHfqLNLWX7uLwSkL41YrJH5ljov3M/SR5PUA3O683H6cpkCZpIFv
5KaWjpnYcKxcfq+tqWeJwlTZ98fPVyJKc5EJaA29Ph13sv+FHb8YUQH8L1rO3qdEJsgKNuR8wGwo
oiQOcw/NOJT6fjXxpF831lZRn4sGXmG8BKlbFhg8b4fh8KBd42cQkiDF3r/80hcYtpb/UJjBG+iJ
mMar+d1cB39nqW51knaEqM0ob4mxhpaxQkW5wrgRep/8W3RHE6EO4MtORS1XaJ33GSW4DMmsOE0k
uqhvJabqVBozycIOZKuue5rXWNbaY9IGoKIn2iH2y7rjM22OcnyhH+GmPnpVuGnMIpn6SW0qXzbs
JbE8tcejDUvQifuTtMDQnJ51ejS3juWkrMEDryvpXqYe0zsKDkpKeB+6w9qOvObqY48mEFSPoyE6
N78jpdvUP+ZNFJFC2egLNKlX6J0ufUPZDnEKBMC01L/bh9arrVdanhpSOIeejN4OXYRsdbzEJNop
oPKkt7It9SSd2vNkUe2mmTkpBicdSIvQAordD/O+zvX3vS6249LoVDPR0W4TB/J0cBYnv41E74Iu
QG73o6rnI5PtW1xKEcQmmLPGxLrsxebrhyvnd7zuA7nAXfoEbxUqzM7oAfasx5DTrGLbOvm74WJa
lFPub2MPQVjhgmS/JQSw6B65SJF3T3/pyt4Gmo0OlTkjkjEmEJ/jIjj8A/Z1uiiO8YiT4eUC0W6T
3HScbyCVDsObFdAcsvdXAX8noY8I7gcTZcjhAO+GR08tZf2RDRrWolJ+3oLh112yqaRwT+CRrYHd
2p0vdVSaCGrXXyLDZvEXK0qGQROEyJFNBqNdW5X9amkrcuI2DRLrm8Yqkt7W9tLoQDejdOk6Ngt7
OWh//BFeGfZ9m70r6ySG2lVlx1HW2OHfnIO2y3v3DPMHKeFzcc283QaZWDNGKnE1hhI8aCyH6vP8
TSlVOtBr6XVqbzRoR7Kwmt+Ixjg6NTHRfJxE3Ur7tvDZuBL+haDwOPBe/x8gG1XRDfqNZBFGtCY3
kcx0goxustg7HrJzMIFgN+yYemYB87Q+AYyCiyUM690ulbP5LAVf8AgS7KhmLU8NvsGO2gfc5Rv+
/p/HpNoXAV48MKE+T7NApBrR1HGWqjQDtb6vTqnCJ5zDFSZ0e8XnOHV/duLfoA6nqvNOLyvBzJ94
d3BgVolGZfXfvq53FLU7epqrWsWSmHIdnn7TXX49xF5VuZ98PnabPNUU7HSc5NA5pkqOrhx6OrmM
eCcRAfWicLl8NmbcUHGC7/vvNtya2oCQCDUgl/grANO5s79QU4JmfpphGXDjYavN60Qk/FaIhP1c
5jzsoOnVjBmn6orcPn8PnBL713DjtTAkLfXNevFxn4Znu1TJXf1KAzLUlvzqqt705GYVTxaOqB+M
3ZRHVSuip84eJDayqn+jHmUAh1FtIIrQCo71ADQpha6jtWn8aE4V1I5XMXKr0VRYkqBJj1J86UJi
ztR11i0s+bZWfCvhX3VbG3mOfj0PXSRXJxTQQkobPPL1w6AvipOc99MdTqpsQLjhPjCTL6lmqoK4
UXkIGxVr5nvsiflUwmY2kww0UUHTtR/GFG8rPni6YZDcryaDh7Va688aNKgbrLLyBL/6TfdrNCm6
JS1EwBnPtQrHhFOC4oBYAyzfY3cWXY4SnFwg/SSgXCWKKH15cDJfaZzXLBtIF733W0zks1w4hvnP
2bSFWlaM9TZwr6QXjXuf8lx8Ela3UvAeaumirLdd2BS8AZPX1QDyJvQjObK06cALbhRnzft9uGlS
VyiP0ERVsZagKpzFpnkAjLVeHoPAuStggUjB5USZZDIcoBdVFd5gUmypvGGnIhoxHfftCbADg/bW
fC1TeWxcNRfgD54jNPf35j/t9xxX0wUdyOLwMD86tLvHqrWg7icrtazMST1wZHZPt1PaKFByuWTS
tLsua/uQyMdjjgEmHc2KP1b6mqZ5AdbdiP9sYy6EyEnK3xhv2FH+Cjx913/k6ivXoR8sS9ftxNhS
W43nj053xUUXG+BHqz8SmF5T4d1HnyVTn3wZrV0Nq/KJcGVBRtM/UtKOfEkfvuwsGm/oXvHRTeFN
5tE+d3rRkeIFeu01rL6zwARgqiZ1YM6VGXRUAApKsuqlWXhkJ620JD0dR/aSWE7YYLTBAYiKEVx7
BxyjS+Va/Qd0Q/V/DtEEJDVotiGWVA/dmZ1AOa5s2x+NqqugQU/dZ+MBjTcgOwFpJKDx1NkeIH7C
G9PqfdRto6Mg5U674S0YgGRaBDBgcrbz8agamfsnVXowq2LCcxeX19bHO8dgKkqpBfMYNZtQNx1Q
Jv01ZpBqwB3Qv+TWUPMJ4d4Wssi5r9IdkE/p1bFS5Ghs+NdXgkrqmjoRMUJbz1IbB7hfm9nQYmne
lmI6hij2HVlMZ6iN7qFI/AAd2BwwlvQ3qtb79i1ULFnBH6yfKKQlu/MkeXEFIRuMDy9U8zzfzTuY
AMJtoei51fMA9voHYEX4vDaE3o6LaLGfS6ukyk83gQekDSRkD71JvjsBZXG1xW83Rk0gJl7nk9io
TJFXewGFHRvSIrToMJ+iHi18N0obe9CR277Mhzt9Rr0qiTmVo9pmU72OZYhYJ2SoRd8SZzZPvvkb
QwgjG9r1iaNpxo092s5pyv9qmy+qJ1nDkqGGcDLPT9480hUQHVOQVxsSQOeMLBPnGPGloi9PsRxP
MD+xSGiW/6yWvaFUzhR9JYItfWG8ae3N/Au5duJMgczfxV4gYuk/S8sH7eexmFlxXWMPsJlpjmCc
U/8aW1Nu3H0UcIluVi5/uEqUZbLq6jQZe0fugwUF5w+smH6q2L2H7gjQlQ7eevkgoNmqFzr26TkY
coa4q3BE0EdPpm5rysAOPkzzagSd1UjCZFX7M3GhCaQfjBy91VWT+Pg6tdJ2ZbGTXHjW7VcBmcUT
wyCW40MQA/krlIZKYOh5QZtxNyY5+AZNZm3b++asldW0P6DnrYI7rXfDeVO6fnojVcx2+mFNXRNp
EG61eETtCoD4Xx3+jjyUy4Xp5Q+4bUYvtfsswNSfI6X91RPTKWf0//uyUQMmdrFW9HDoOBE4Pss3
IwKpfM+ss8UN0lWlBtGHx/IG40cGg+3uE3ILfTg+YJC3M0ge3VMqz1LPq5jYJidkngo2ZcnfNZj/
r2C6GUoBYwCCT7ICdwCCIZ4AQY55tOpDXdkD7zDKaYxckn96Nfd/mFdf55GCVKCPl6NScAkPbVqh
dpX9KGG/FV8F4wdRvfrUc48CVJCpfuFsH/l0MZefb+hgijuU+UMSOftdNula00O7RhAzIS5lC+A0
wSPTR4OuZ62GaX1hDyjFiUZihrZqMWQZxOo6TaRkp+cRY58tiPp07Z95QnnGAPEbSVSkg/bmgr1F
y5LRq+4887re4cC7Ot5y0Q+ULwilmHPq052V/JmK43cQV+73ZAlpGCH4ESluvw/nr3JUyq0vvX1E
qQvh/a6hvuVUZfL9F2Bm4LRj4W2GKNtqsxVriZ52y0LXNRbobsM6twpxerMLatg8GFQjXK2vSa2S
uPXWDkgRftIy9obi/QHMSf43veO0BzhQEZguVcC+PBsramNFrNhnIm4EIH/VTOmQB80SMEYeLLKG
1ksdJrTTdDz2bA27+Qxq7IbDRGMXtdGh+KTpc3AGhK3GSUc5H2ArECjEdTzji8kAwJ+nLLzt1GgX
t4HlUAxr5SS3RY1PulfAMb/WQR4ZNPJIihEbFxrC95xeSZve+xkI3TzalZk0GWfGO+2Ei4sdNAh3
3yaJQ0Z9n3D7gj3dlScsM+9WsrStT1XRhJbAwf7w0efrxKfgMwhiPQYPgkRgXtUv7pWSVq+hgkVt
MQwQdK7OH89r1R9CW307/c+W5Go9WuYsBEiYMPApUzU2ReSTrvFgPzPEtj5jkDIko/xnNrguoaxG
Ea1x+DwBiZHOweXcmIbTvIYlBznNAcvsbADGM2J6VMZxRN7OON7Vom4DESAcb2QJuxHvqFJONZOO
hLwJDgGdgMfAAW9W8zoou1Adk53pFqzbx1uy64qY2pCUkoKItr3Dvs41WXMEMR8atwt/iX8P90mH
YkR+1DpJ/IlXJlv8M+FpKZzZZovpEUkFFyhSeMo59Nn+IpSbnyTxtbKJGxF8w+MnZLvBd5fnHChx
Cw5d04GKLgktAWsT7sLUV0oUzFKigCdwuXncTkqZt2UbJ1gKYPjq3bIxHe05KJlLOOGdvfTf0e0Q
Susb7yuRacWdn67CBFtfkedEZZ+3xKQEVQK5734HbyuguMzH3M7vP4CHZ6xChsjaYTzf3mwpiFLU
yaZOaLaBzkeagKOYKCLCyLheRLNY7GeMfHaEGcU8wQGrmmypuCQ5LoBQQOA7VnNqXVIe5CoffTzB
OiP2O7X9CSVc3WQ73v7Rphjdhb2eqLL3qQMgsY1cA2rUnc1vwCRoNmDDRWw3HgKI6KKRCy7yMmyP
7pZSI8h0rYvUEz9OcbsenRDLtW/PpI6ZyZi1kNXoivmefzuE0g4n6YEWzedaTM96cTrrUqSg8iVq
u2j+Tu4mVYVhVQ0bU38eGyl7KYvF9Qc2F/dMWqch4dBwWVP5TfIs3GUuVdMV+ePftn0iFBJanjWH
Jx+Nx5VNJY3mpetYsas/B1bKCvvSI0UDPpTCZeZi8YzM5FWfOeSIY6fCYSJ6VHq6D75NZPP5TOOw
ZUr1AgOSRL5/Y1fdepYxNHERPIn2a+/ZnQ+quMWOS6zUMqdch7wu2fY1UEUaFAlXtv+b9+gf8mAO
19m8LEup1eMyE9k3ox2ko3awBCOkOKop8PGcvvzDNbRqylRvE61ViT5Y/QjAalhXOJkj3W424sSF
+/oS6/p2pUuy0e7y1SwW0qD53GVNI1IHTRlWe/DPjiIyHrJ74/ySdAyWGF6HHFcP6NATD4ETQriA
N2uwt/Y7svCxYjidrmqy9t+7IxHkdUnuWjcs4xFoV0nf00VrPlI2/q0XBUjOG+QxGbkHV5+lmwC3
KB3i0rUWSDmsM1b8avjXRHyKQV3HJCQn/3FL1o8yXtrwhSz3fXAkntSg/KzBqg1MxRB5VWFb1q97
BD8hgRmHoGsdvHX1XfJWj33hzl5ED/mS7u6JQBb0Sz96XPLURIBFHy1IemK5GZ1lBKKOUHCCq1rT
hkuJWkTuJ4Pu0jeY8UHlkK6FxscQz/haFvS3DhUOSXuEtbyf/B13XE3H1yIbYLxsKm8fFa9JcR5v
bygZoH8ElowFI9LWaajAdgrzqtJUHm2id0wcNoX/YJWV8lWfVkuCKT1V3o2Vev91oJlN5g0P+q/j
m8pgLDsP3Fjssfado4pML/Y7KLVOT05jg7tp1F+B2pdxPxvu4oIGXbVLcwCuAnYXO1bA7PD9wkQJ
cFIjZpaUk2M56ZGP15/DGaoU62YiU1YlXon2qJ8ysfjQYG9aMyyG7tdhGNd4U6t+LuOjsBuGfsg9
q7zVoCk1yzAavVLgHqhiIUna+iK3+V6+GtV0gWGnvz4PVolqdBjY4HDQQPf3dfqIbQ72Wtna/9XD
CNWN8S/JtJ4JlGj3rvtzhXPilac6omXNVL8quyEKlf6ld0XQF8Pao7vkMgyUA/Hnds++PX8uXv1b
8dyJu6/DH55mCXCZdzrHBb+AYmHxqbOtmE8U1ekKXEZTUYv12iShg+725rHATLpo9uAXurFhhU4f
pCQbMWrLlUQxN0/PRU0kGQ1qi+ArhMQOUTMvFmwobmZkMbTuKAY7i12NB0vA7JCvKRJq/HL3RYJn
yWGfI5nP2Sh0ResxV3DFd+5IQ120FikelJHW1Q69qWevHlOLKor6VD0UF0jGICE+NaxmcVij75Oi
kCUyZlW+QsSXuZrxexf7Er3Yl0E9lZE0RKZCtwlPntPyzc6r8iEwt6NkVCj9eHemkjLyfe2/558W
2ycfvVH5kfH179WhmFmqQOIoDutmYbq7qX+Efm22rH7BEODr6cuXsEIYZvjb8+QMVEDN6wKpKmoK
vIBvjEqLLQRf2aLIenwn1wPB6VrUOX3cNf4owY4opPYV1ww6S+cKsZCply0uhhWqS066j2qxn32o
nODiwMoaFFnoP7ZNs6I5ZE3sMc/FEm5ybc44oOKAS/4ZAYhlta7jsYEEo2bUAZ47yUSNHRL9sfXp
LvnpciRawRdD4JMLUARXj0HORb/1543YRlHZUwJX8HbdFx/LHsZ4VDk4BEkXSJ2zisYVIAtY7WjR
AC41tesEU22fJiiVAH6sNcePRmxxPc5i7hKNtA4VX5EnJ39ROZUML4izI9ZdLatycSGdZUMACTON
22NYWUDUrWW8iTFOuZb5/9nbGgglpx/ZY4hIqx9DvcToU3jG7MXfkYHAjXkrDK62mHxJta2+1cSU
00mbXDwav9i6HsXnIchY6StnNg1OGtzxZR4gKrhYZavqJNIZYSbdqvB3n4CJa9YzJMtsVCLgks81
eSvUkLn7BUH5uvs6aCCdUcjaitknX1XyjD6XdLjo0vZKyR0wrci3ZDfLtj9dgXIRsZWIMH3ij5wA
cLXtCScu8O5LRnz/c1uFO6M4RXU5F6S6Kztgid3V8GwL+Sk08iHYayZxGc5/p2Lp1EbL7GvLeKk7
zEhIAcLauc0ouhUTFZyY285a7lmZa08QrCdutbAI/5ORTHqRYQEefK/dWY1Y0GS+iumhP8d8Gs7L
PBYseceargF7nOG7SJJymal+Xnfm3CsaH4i3zvF+KyUbQB5ppzZJr1VWz7a1aTMk5mkJKWrXDO+j
g/QhtCsnDT1JpBJCVfE9gJmZJvka6dIplTeqxph5RDSqNl4VL/wXmoDo80XGC8kF8vpYCBTobtCa
aqW53LYdc1HUjhqIt9yWQyQPt+tdUX0EJ9Emclozn9E9m26b61nOClD1lFNhcb4hZvC86ej7gdiP
LLBgP4qnpWUnsE5WCC0XsFwdWqNfa15JTHEPZ8Hw4iZ0XbMkLSfxu9VebV5/SX/LrXnFPW6FYhII
PlVMACxy0XJa5fCyPQ3HqZsHU0gyEqrFZwY1ms6gOY2z53HxXpWbNilvXlesW+m9InNa3PJxNeS0
0nDcPABhsPtpaU1R9ib3bpbbS4t/rs+CuQOtY5I9ajuZFf3YXuwIFXx9bZ8u93tDl4rSskgJA7Ao
ll9dP4saCTKFmJkpw0vG7eKgPB28WOidCSCykRfHffRTK3+XYs9JyVo4C5CfL2dSKVaGPtDZ3w66
xc/KmXqxPjRO5PT1OQ9aFVpADzCTVdwRGanxElgLtolFjFcIIsxJL4TQsUfLb0msdEUxMiNlM5FK
F2VZ2fEKBHKWItmXgQ6qQ20VR3kc9GEu3rlfAo+GOqBErgQYZJCtA32dd0FbICAgxEUUnHogQ3lZ
k5mKdoPCzlK01JNKjTOP+qRDwj9la/bR4GHo93vfIEBxLHQbUKchFbMRGET0vphHfZMNOXLBA2l/
vgolSstnJB4wp2iq2T/gwwxhijfcnfaqK3D03C8zDI4rc7z9h92F3kkU2Hc5QOynDn7EsJmk5JM+
f3sRite+GVBEUbRKe2Te3WZH2nFbK+Ft1DdVZ51Y8Rgab9lqcVecJrHARx0csmtd2TlpSI/sZPzQ
wc8+Al89EryTiuxJdxDseLvZGjqHvDDnjU2gu5+RhU8zhkvUYYw5594ymqyxLUm6fsS4db/7L/r9
OKVdG94h3f3roz1ymB8PhhDD66vqa7MhPSowp3LRmtnJNFZy2rgFoZwyZjpYtL7URUH73lqgv9Ap
BZXFnuo5QoJN0Vnw9yFAotoGgx5nzTbjYezyBXek1euHRuc8AhNPFzCgTgfr9rQjCLJsVLswaBeO
mJFtg0ihxH9R1LRALTQusR5EyTiqI/RwHfcQlfLd2wahc+u42kWVQNIUPsU4yUK8Z/qY9pkCFE9B
EkoKUyT3Ha2Fz0hlIOU3+qHFdupeni4OapsshLkX/xgjS4Dd7Ck4S2futc9R0UBnrUUxLkmbz4rg
HSxg4ZrTQ179GKki5N4T8RlplXMC6n0JcRSvUx2x83rb+9pG81+vsHy5e5gAO+QWs6DHv2+/FJlh
iZWf3/82GYGiiUR18Tj2D6WTpxYW8JFK3kZC41e8NegcK0T8OKbjMSJRQMwcfTjacsDCySqCkrq2
Kng3v+MKYY4AcCsNyRqc24vntnWLAmgdMx1Y65Eza+A44NfGXi04jOj4ntItlxQ0oUZiEO0yAwhs
D3x0LFhebKG1wJdGsjZM9f29bIedXNUA/izZXwgArQTbaBHymfpFEpSNGxowmTKQ+h/v/M8BcY9Y
3df6fzYM8OBl2UBI2XMsswuaa3xXpZOWDTKAHUnBbqqahLclSE2L4kydCcua3YCcB2Pwf25SsThx
LMuUZWa7cBuSlt0YAkrbMttqY+QNxozZR0VQ/eH6HtPwy+wKp2NzZ1PC/S3POM75LgvDmxF0J0R8
oFxkZCYPrVW3NNMY5dBQ2KKRgTRPYrrOaeODl+rJ/Vdrq7hjNzKLoGQnIJsCIf/JIFMYAjpLP4lw
KK90HZ/zWyLPc2IRNCFtoYeALevPk6aFcTFCu54mig8XxolxgkRmXeKuE32UTN3kEfRE9Y4bvdbg
foEyImz7JaPPlGODKHhM8Ww0ymrHIBtXRwbOe/G6ViSe7nQlih4jcMmFyF1hPFX6ySxEeKYAJJj4
J5f3huHprK9z00srkNCfP9n4oo8B8qRViCO1Ymj5c7fUIehf9emzdcpnx3D8R1dymbj9gZ9Dz511
Aa6wwqRthKd69RiOL9WabqpvCDripMpK760+H8LJsCHSmUJHD8pdDt29LrA0lok3AQw2ike5GU33
4vgSu4s5ae2KiCCvupUjxq1CKSPoBOHpaqqUxVVGS7B+KRhPsg8qimwIlIiypxSKC0a2K7xUjZfx
+ZJhoXrEh/xEZqO0xkI0ECgRPczDVVY7E1R+mTJJcbbRwqM7I3LH3nT3EFjmLX4FKYS6Xix5RZq7
OK7rhVyBn4COrTvj7GIClqq9pKrYZMyhokTxI/NA6OP88Q/7j2uZq3iSDnzI2M+LImWhMO0K0Xpy
Ih6TqYRLBvc1s7Im858Kga6Y3YYUJacA2iEbZyLEs1V6S48m9HmS6aujjpQpBBEuEu8HBcxjZpm9
oxYBsqgXXmPq2IHwub7AudX+Plo2czZ7Dhki5XS2EYgSRG1UoGymnQKfkuK0k4KFG9ZlpzvKIoeX
7Ir/a+jBIWyYiLg+mU0UMkG20sF0U3boQIzf86hl3UJDOWePU4bJCeKpQ9Qjb1BwV372eLtnjrX4
QbyZ3Pb8VjOdT7LzWdnEBrK2f9/CWW0M3aobhJ363LVaRFSzjNwzPYCAALVvnJhpoktl6giB39PX
rOj4/Rcc5lukyDyNnXZNpBzdDfuAleeElPoCcMlJGjfct+q86GvEsQdpKVHv1xGnfUN3q2U8N5lE
GTrT7p+BGwkZhBNTfYGW74tLUFCCP6/LZBC8ggMy450gMj4KgD7kqG/BZAn+1JmlCw9Qct/gB52c
vdciPnUHDDW2D7QI09PDajEmlK2e7NFIbs1nxYKiNqywOYA6XAExYOOkAStCiuzcuoucXuzQOU1l
/FPGIKpRs+9pTDDOtMwjG4pfAdZmBZTub3jjCc5KBbsAkVDSgqBgiWLQJ6RcB9d1paIq7VrQZxko
NYHKOR9NEJN2hI5ctmLTv/mIuoad6ShJfgKXNuzPXlAl7Q0FRvpHsZC0mgYlQVlPK2PeLpgJMUx8
i+0HOLRFk+65z8sNt7xRtaOrVvPxsCgojJY0mFs6seOHp3RUPA/uRR3djfDbjDoIRsN6Tnvvrxlm
Hh7dpzRX/vdAFDve7WCLp+myvthtyVO+Nd5FuBM9cxOA3fcq3ni4V2uELswZc9X5MRtQhhNAybWo
DBhFdjD9qH1sLNNh9nqVUrjvPS4d4RpuANhN4if5btcslai0pr3ypWO6ZqYmraxA3pgmF7trOUXV
/9yhdORUZX1j1ldMXXRCmJOFMrxfQJP8AzBIemfuzDAESdKdDPDJtMpMtUing2KDenwb+fMlzYEW
k/K1SpBfKs4OdR3th+/K1V4Rsh+pUDaQetB/TOhTyz0vI85vTe9JuampgeA5zNpGC61m34iGri9Q
cUKPALEUeR4GzTkQry69pyRBcmK+vbHfOb5Dx2UopqYl7NkL0XjnViD/jcJcz1X5Cj+N7LJ7i0JS
YdANNstJbW0e3xNegxdiwEAEiK3ARyCHJZlWO9hp4Blg6yBoZzuEQz49bF6y5uxIOPGT+dSrCexk
F/iGSIn772JIPVEoWf/hTqwfrdaaJbotXL/Hpv8HIwwbclP6kBqLYQWVIJorBA33wvJlLVmeRwL4
G5VYJJoshKddbZMS+TyG720KpxgxphlJ03+suCfvDHJD38DDR/OLVn/SQj1euUUHz3/xQrG6kIFA
OIeYxrPISOAzmTMc1ylXI7ZXIJpRIWMQaJDubyKLCANzyE5fd6OtOdkywwvmUtP3DtbVzmXFD3UB
8+8bThq+jPJJnjCOkSf0uTeHkn0ihprkmYVQ3w2QstXwQEUFdqIUddC+sxpMVRr9nvGpNu0zsqmu
O+KwqZ3/Fb3XZ21og+EpFoYx9utlg1e8QL0By+2JDTOQlON576KKXvadjXpc/0WT4X198dyakslN
AcRhEeAyR9wTKJr56LZj5RudeYe8UJ9ke5R4Py58IttLBhVR6u+SW0K+DufasuZmZq3zTyXPDJUr
VUviYntZtZg/xHIdkmcE3QtmIZsxqyCKKuRSjFwpBVTrZXBAG/kBH51ENUCwWrilVyO+MeKXhheO
tJpASTBhGzYF0xR60m4ehAVxYcmYvJ2NFOMsrRV2E0qdUdM3evOgNuP8YQEG1lLqOBfe4o5/VjS4
IMUGj+Bbc5c/vG+ohjvyL3DKHEf1SoxApKoxjcr8y8qbKIQDOWW8QMRUftoDyAIejxn98CzZZv5q
K95RvRO3ftXug9oS5ZMAm48JA6EcefVLl2kZ91S6YATH8xEIChPcFuEmNJ1PA91DmjgCtO6hYB1l
FJboCrBj+vhHt2IfK069KQO1zwF0dcQalERIgB/vcLw+ybNDgFRQjQ9ibIaQDDK6GIs7uG84qpwh
pr7NPCLbmX73RQ2e+m5EuI1t7A/ICC6ROSZ7QjsiTvdl+82wQJ/sNVWATHCD+oxZNfsoBmk6+cST
I3YtdTjDZIZisokxdIQpzR3JD9z+JnIGlRqAAGc2rEIo4x4F7mtMesQTOd7beXoW5YpOqS2vJ+nx
hhl2qdJJHnz6Y2IigUx/KAFV6+b02grzsJFI5NfpTYRat9VK2xd86LEIuNbL4N2KoUdbmlxBBUzJ
8GhLFeUXPn1w9NSf95KLgihl0rGSsOgk3QPTaepz3Mr98hVJdoGZ9iEpAifiyfxbwG3UDczDETOM
vwS9EakwgB6ATW1YriKclOZcJuAUP6fm3UYWCMi7jRdr4Rg4iQvV0b0NaO9aiq2C8B2Xqs8imfsk
jwssIU4COI+mYPUWNP+3LWpeeiRkTbbPY0ZcOtUkFZBSvdnRNoUkOZsN4MCP5TpnWW7KjhADsqWs
Pa1ZFMWNjSSKv68J4bidRW+hUJ29yyIcXa0GJbZUR1K39K8FlmhL8MZ8s9mqoxg+K4lOANan3GlC
+EO6kIIHlDq3NkYIVhqlzHleeAQOHAmsV6jqvb5yeFvRz/qeTU3gphY5jO8B+H5rHUYGFQqaftAq
cdZwC/6kB6oq0uQtsGoMG1Sjgf6perzxi9GIl6FdHV7+J4nggb5Hi1j3pJidw8lVM+O8RYA4Z9Lk
y3RpUeyGDDKXHBnKDUPHWg7uLddpE/rkxkvaqjTrr6ajT2X1ccgvEH9nbNH0FDeWR9a5B2oh/2nD
yrwrdQJiCGiyMdc/8OnYL977bkRPJeIoqXrEvYnud5tUu0w4VLr9+LiRoiZKY0u7rpXHm7SU58Mo
0DVwxsLV3WKp06RX9NTIg5cvft9Prwh1j95vMMiWNrMxZlj5ozJyUgKX5EeQZSztWhxVoduVx1z6
Jm0Hsa60ODaz3n932ZYl5QZk4ulG/ap1/wd+MD7PCIuaIOt458aa+HXJheqWRqljTKD5M2yR3Gz2
2F2VLvyn3SCQcqew+8Ty/zWi4U2kDx6cMvlE5xvbQRyz7VpbAx53S85WhQGN5eLSwP1NpYVTiUoR
PGRPfaX+lyYFeZSEqvF7xxsZfmxFIXh+rr8lV8/Ty79dBf/WPBZ9z4DKcSQ4glnMzpXKTkFYamKJ
9KPFaOZQ5Av2P/9njIEkcrLIGCEZi4hadKmbkseNzJjSNfT8O/2SUIVe1R1OPeFVacK3IfN/EnH8
O1vK/yKYkLdvVMdQXobbqVeX8TIcjdwOpk811+La+uvONgDeJLX9QbeBgdX4TmN3QMWRsmAXF/Zr
WBdru+F2AjFW+RlhqKb+RHPSAu//txu10ktG9adf54OV1I3x9V8vPC1ps9Q3tGmw0b250m3C8yqF
oj4F3KHzPB83oCseUCNvyWI5RLYTekw3vSFtkilaxA/uacbHr14Q7nGbSGb1difo8VMCjMag+qpi
NOA7PlIAPGXU+B11wiarvLcpoVOQXZOjpnI/FpFovc29arUo7Myeg7JH1JuFgpK3+O2xkkOh7oTQ
6NvMHtG07oREHRteRXD6RjJrnPnZndop1kJ+6r1PI2zpUFYiecmuD4ZupdFX9B0LbXMaWPSM21d9
Gh+I93PUNcCtjKdw7jUk0UEypUbCoUCIR6EcKPVfVVUMDduv+pJ+4NHs2vfmTYMQhHgpAHvajce0
MsfHuwWxk41++e3GVQ2nc2f7+FPydrhi098GOLYWjruLyqSS5qypqEIzJhoMVb5nd58AwLN9fgUa
ElLQHpNw0ewK05vrjYfgAWGYa72eixcF2e9nQeCif4SfSmNp2A96dvwjk6hYD6cZHKFIPl713tvg
DNBQc2ROTkh56kqiGhVL9XeOiVDga4Qeam15nu3KZrKernHjurwCzcOooI9f+Tp9iD7VM8M4YCLg
rF7tDVnMGqSY01cTE/ZKrgrSPGxgZuzwyy68RM11tGjzWOxd89i2JkjGnsOdce1SvGGvDbZgFu7k
hEz7p7ZZw5+S2dCdCawx9EggB8F9KP76bEvIxp0HXqHMi88h+eYmvw7xhw3m3PM/KBov/ewIovQP
g1blAuGwHltfvz8tgN82DW4VVXcrpd6LBn7JXdoHTtkZNe7Ehw7KoB3JIIQQHRasaWf7C7g0Uxr1
ObSizR9VkyxnWjUVdIrLeIRWorAQUuuqk2tm+LreqWZotaBoYI/JhJ6P0VVNAX/kkYzqWUqCCffb
C0o8K8b9k/vFnL3LsfG6DBoQ33R8iK/0o9VlcRH/NKv2/+b4NzxUlBqxmqxfsepDmwBU8WMsI3hA
0sA+f5+/YQOO24bpuGYZh9zt+4l9qxnrZrsBDsm6lA6f//uAetzFJXn6lDmunJFdTY5H6Wj0zQY5
OLOp5qgI7DfDUlFWnOzdylGKiGCagmf40KWm6a9UM/ipk1P8QWhzm74lRZ9aCTcaev1WQwP415M1
bhjrymBeoj9gLTQZYJfxyc05PFWIoERk/zzAchUevLM93jtEikEMc8IS5FwA5Lc4ZXaVJ+QtYco+
dUrS82lOvXUf/whGvn8RKrW/Nf1x7PG7fYw8jGPaFSWqVl/A7MBRR4XFv5yBsToy9UWMEPE27I+k
RX4Pg7TyrrZkHDJ1V1bSHBWaigLp2dZZOj8nEhZRHz+GRMhvOaSYxShnceDp6/d67JiVEwSBfe6+
FjnYwT4yCowen4RnLaf+UpI52KZQ2Qv2tRd++KHp/VQTzEQsvFGJpnFSU9dkNYhZfiW5im+k0NHy
CEm9YxbuVJcRQtUC25jkf/YBEKG08nCz56f/CZMaHVNEXKzn27fGTcEmZwkkE2DV00xo6WA95es0
9WMMXCgB/WyCoKlBTucULO3PJ2weIyjti7kgFt4nVGM7XvrQvwxB0Tatu/3w5nAKx5ZVMwyWVnlD
rwdCg3DygGmXT9IdlCbATOHOHOba5Enky+yQGS6sjKyGTmlaZDdg34dLKl4+1SaBijEaDCjDf0jw
eDNAv2O8IQk6lSCZqyBgKl4693ITUSn0jRYHTegTdhkncc7IuAe3OABmnq2rxtERPwb8DQIDlq0x
aleShd30mZ/cKh+cQzwzBfYDazzn/UWO/LR3oYGQz7qeVrS1bwSDJNpJUFFkgd3vIZ/4Gy1NN4RR
glin2Q/IGe0iNU5cVTQfsrCXwcNGAR75fqiChHlEjvw0N+/+IbT/468I9vfwYqPELk+Eh9suJ8HR
B+W2jOpIfT9z3Z80MeBjg4hXqHy1RNd3Dm4g5EbaK2afGQI3+bGHlpPW0OAtunPFHf0Zp292FP8Z
vxsxpjn7HIMFhzErlDXGJEMym5j0uRj5FUmOiPdjUK7CSW67+psS6nnm3QImI5OETMMVXtSo3CF/
lzVpKMhplnkmpRO//W5o4Hil8q6QWINxiPrJKWYDDGQ/7sQy7PGlds1XjwdsBYXPcrzq2cllW3qq
+qizgDUNODyQXUU/ZmHlVgSv0l1wAunmbvxp+wL1xyuhXwMKrBt3RKsGEchdN0SXik888bgj5oo/
AgL0n1IBLBxh1NGrvLUwg+uwW7P268GDctfK1w+61Q+bNKTFg6V2NSBMIU8ihgDqr3meHw+2B7EX
R1YM2OYm/rkvpwp7fOkWKi7VFPV4CSOYkcKA+JF23PpGxp6CeS5/DzSuXpiM0eGb6NznwC+ShFP7
NKj9mJhuuH3/N3AjBVRmiyu98u5ux9+dLLLudckR7IxvAnoHnqKtXa3unU7dOThRywUgWJyrOBf1
3qTZE2Q4Jo6m3y3hOzNccOeX6XLULdNE6I0bVc25Y3605IMaPpuwtMVRKP7d7aiSdUDtOxZzNhCy
jPf3p6w2GDOzqf78reKj/350wg6toY8IaeeluoHqpkDcKyTf/ntXfvC73B9RNIX42m5wddoRTUMd
hud2oWO6ghvZqzeWSCXVA3Vs9UI1S3IQzddzr4UBAaPNsPMlNzkMAqgz4vt5qK/8367ReMV2dlu5
tKuCjRSUnC5It+J23iGeFFgAT0RN9WN2vaHXjcY6+IOOyxVbog/twkwcyHdGvHyQA0QUfYOiVa4R
rz+NA/agEuy0KaOGz0RcxEO64aCPE7b7TGml7DTYgCx8Z9rmsfcriQIO93u51OzUFTDK1QTa2cF4
jwppyM/peZc0ifiSV51NnbWVvo6uzMjovPYNr5jNbgLnyWw/tfblY61yOqXy2F+zWkHTvtkrBnuf
M3Xlc9YDDsUtpsqb2jfUyAzH0elirZboIkhhzgUZF+DmGh1fkLEe0L3LJTHY2PskYPqxPfvaDJbM
3Ud8+pFRgXG5/HQe2YuE1ayz2saosGFZBXVRbeVRaOE6gAnRb1pCnWI/hcWLXKGVmwtgH7WxNXau
d04dFpTTXlU3gJRfAqhocSdBZXQediXMNmCSOulhJa/OiZ/Vl8avJBV0G1LN6OUco9EdvFfnYnPd
fmPG2phDbHlmro6ZcI3NwRK0M2otHDlSz1gcS3L0vV9oUi5GLIy/8WsZSR0wJH3lfZ5hLgowJXo3
bEHCc8ws9qmLjyvPO/TAyDpdVfJWOjm8BaPnIG4spZk6E5sQqGv49bNrruUK3kODUTPAmja04whn
NPgBBsJx1+NAMZBV0OJ6XE/znpWFx9nxHQPvQLuTiyZvBkkHuo1gB3w+0Dl9CmZtQcf9Qohy/zPw
L2Kj5Hn4tFKRHadz0pnqXmLt1x4ra0tVwJA1J3o/JCA+waoPR91Xy2fuN8GWPsS7mbq/7F6udeHB
ZjrQsh5C4o99VFZOn9qgE59NAhkSiFJng7UCD4RnqXlxMqvmKLJDHuWuD6TdZSdKUr/8y18ROVuS
fswcqgMw10/VRxGgVHfehMsyOSq2t6TAOG2ttOFlPG1mek+SxR+Ouaj8k6On6DEB7K64xroqBvEF
tkCdjiileotHpng4c5e/YP8w7wEw0QzabfQ9sGqaz1YQRsgmzuRwbwrZGIkc/a7iOqXwfGAbvpCq
NttBecLbw/TxWoACyDPfmFrW+HFJ2Vlktd21p3WpcVSOk9KGfKe3OWqTbEbHIRLpoGObGgyKk0cR
ucA3mpmDe/QpOkHSuN1OQ1Q/43lD6wBgUZTKjWZG9ZlsfVR/P4cQwgt8NzW7jqohDkW3Ityu51lu
REBOrelEK8bZHj+tTTrUR2luAEwvSZD983SjjHsy9+J/wE2aknHLzR8bWUNCUnboOtJp8Ni1wQNo
KdrsTxmq1HoWyv9ZmvEtUBxu1mWywVkYN63Su1hXkoA4wkn3/Sgm5my6btskQhmodwfAEToS2YrJ
sjpeF09W81qG94TGkSzm4Ca3eTBoSIc4ZYWv6YpShYek6NNFYN8VKIOOjK9+2iYSxY8wyTZvjA4n
G/fpLlRjSw7yvUDWKmo4A/SlFAy7FMyGDUbVFu4MPW88sPVEW509C/LXcPwDJa/Stj0C4aOM2PWN
HEtZsKacpe5eba2hxN/DeO4evv5/Bwg5OITS2ty5WmPeQHaPvB8WeOuOxlkG+6gGNEPhROPk1eBU
zQjBszRQu+pb/qHYj2/7X098vrbM9z6rdK8xx8amtJXIDppBEnPuzpZftqoI8dc9tKYnRGdNfp3G
S2281phcANxp3Of7qRX3JtwFiUb8bv1v8x6w68+l96n6GHZ37X42sRKPi5ppoh0ZiraN2w+QmQrl
CAqOzWlPCS+MXuejebQTbzfdn/u6gZ7M7xmbLWzGduFBPqqEgL0GF0Hb3nPdExfqDrV069y87oDF
fJ7W0z6fpJX4RyT/3uRz+3SCGvAMYvAKeFWrtgN3EsOkf/KDXaP82qUwQk5xp96eIMooyc5SAXAz
2OkygXrAI0qv3KvrHMz2GPtRxA4gk7SHk2YVD6zCkTK4L3RHi2ORB87Xx24ocmOnDWZgSF/06Jdv
1qMXyLVgod3q8wacaPPrltcr2qs0oWhUF+zwEt6iUNL5ghZWl3HsfRsgnnzXTmkzrChrcz/YTYqL
udPodq5+KXoarF4GSoPikaLXjMB/wEC/ASrmfZD6MKONcVJ0o+t0YVKrb8Eyy08FoEc9KDZFxOpE
jWIRR4A+PlRLeYIKvsKChUYLU+1k+7f4ZcOwu5ez/Zk7xF6DnlGcOzmo1RJAm9z6ncP/FR1+BGkS
ZmSqWjFQ/Y8rmYNPrvjmz5V/bY4qnwM8/IDzuaXWmKNQxOFI0YgPT/cIPtt+NycAhvhKIqn6wrf4
EaLnJ1p+6RP77xB6jYXrlSFtPLQI30IlfjlAqy1t633oUvCVzBbqPj8Qxp0gUKD+3jKsfLCsk2vu
qBeQ2BDXxAn29dLZcw+2Fpnt7FHtwjEh8Oi/H33kAt+Z+7bKzfnvF6K/G9qD4fq8BaySGHFIAVG1
Y94TmM85gyAkkFeDh+0OmLCa9WLmCGXn4N91c34huRnR0WUOQcUbubYa7n4hvekzHrvcuEQmdvWv
LFYbfxrXbXY8OoQVL8S9t4Hu9BprVwTnH0sM8x2+EBX6eGh9cPxvKbrceywxdZkcNLqx1dWPtllu
KcFttcjkpSF+zv9Z3Jz8JvsOYWny8ku/OeFmC4meAbvAfFqu3kFJIyq6tWt+nLztDbg0lbFwDKAq
wFSMr4Bj5fFOt3u6nd82svc4WEgfyK1WCHajD0PR57xqObjntWSEEed91EsH4a1Q2macBVHISmKC
BO25K1eSMlFK4aBXM8U3t7gVza5G3i1CcQCZu4tIKAAa/7SpmChD7rOVMCHF41tpn8strTSF2Zfm
MyMtqX/708xTn5dM6qTGa1RP5AzOIDXk0MSujGYcG0VneQvqJ2vD2+iOeaV5YdeD/lKz2botB2AI
ZKovhCNDiJkrmFPMku6TzKdC/RlB4G/0tTTudKPcuRaMf8O9KW5sW5HoMl6ZMV+hn1+lD418n2I7
9GTUBqtZTyLiP130lmCKpI+iaGfl+tDzHo0PoLU1L5V5hkjaMPftYvYXyqQlUWJK2LfRY8Hr5PfB
+B1PTIXN7g1p4hbMd9VBHtDi8mkmZTGjTDnalvtBRliLKOsli9+Yp4fAb1gJlbbBmLKD8/MTOnlJ
47igrUNk///0oGnZ4myLWRLTkowSm4Ftiyj2feM/N2UI8s7w3vPZ+naX1KUO6K/zbZqSlEhm/GQY
aP8DWa5azDu5sZZYNETcZlIDvF/8LUz3G0kCfK4Z4mldW5Bi/jLInZIy65tqr5fzbrfPuUoFV2pf
8j1cS/yTH7YMmoH7NMmsWuf4voAZxgb/yUAVBuz/DB6/eYDBuYS2qyz6lCZJm8N/upx5y5b8HDiH
1AtCFZjrC9cQ2Zo1BYhlxTO0JjigHjnqM6vBYgpmMrUbO3lK9bo2p0Z8SwTxBYyNLKsg3aYNwxn4
MeqonQfoI2AfaTCMnG4Oc0L0SEpN497uINQmjYmHEByG84o78yLQM8AkXJU1QS/X0XxKM6P2WDgw
USlYd54lGjQYF6lwTYnbpuLwY74D50eZ172vzooISdrnzGC5VwNz78IVkXkTbeRJM0n2sARGbVmx
rrR9t3ldgvsAmrUpFq45kGasHm/gkDuxmyHj7kBMndFT7MPfdzcT71CMrk0Y/1Lo9sKDGaqMBFYW
6WEk4zppRYogBnxgQcz1DX+r/V8x6jVAGwoZBb8WJV4Gr2aD1Ta1b15UL7Ubk/xv488RtIOBPGL7
tiFfDJgdph70y0+rq53ouqjC/r95Fzmazsf4SxIpUSSHfxriZ8BkRqzGJPs1hUsmcDII9DLgUA0j
aSH77+5n7+berVw9dYyHJptGQbF24OLQL0OG/pzvSLO8Z/9fQfV8qatH8RruMILuGNBMFKK6B3L7
aw4xvT/USv/A2536xlxUv81HQohXN/ej4tf9gznKtgDDF46c/0fUskM+1JOrqTzNH5euRKbNnjgd
8zO60wzRcdbBIaP+M5dikS2loUCXvgIlK364QIFtVxcr4AzRI0qCteA/GKZe39FcZnS1TaKDW7gh
rnXI8CcoAiSNoemHyIwdWOBLvYzz/VMjt94JK7rzlOpun9X2S8f4zKMh064c+6M1bmBEIPOFyFAY
bLK3eo+Mo/ZaZKqjAaZXqhSqRbSKrM0mUMHSJk7T7NzPZOu0BBY87NwzJ1e4neRbd4wQ/oMN1yQi
RQlnKyj6mpzttNQlZabppIrcsab+9y+ZFK0FBpX3qgHRdvJqzT3Kp319Zdh4g2Hb6hZSm1ha8K6i
sThv5fegry/BsciOw4GWP5/Z5kI//czkjPqpXkLxYEh2hfNfkVR1fz/8lgmU08u2yEHgzYSJbgRp
3MbEJNC+7RT6CcGLRgbhwgGZARbHGj8Ulwa5ivpiOI2mf81D8P85afw89DfwWmCb6tE5wtjwuqNT
IC+SlbV06+7jmeWzxNcLmFp2VrEV5DAJ0HVmd7mCHKzih4j+cWF/hEMQujYDR+1qNs7dHmuZ4Yfx
AZuB+tDiQx0M2yNxO40Kw7Rb95aw1mpLtQWswlbeqoaY0beB9S/mKAQrjq90xiuk+p0wCI6Emucj
iBwa3+tkG+fzjIDRUNsVvK8nKdJuxPzd74qPKlwUWTLj8D11luOhsgWARBg/ShPjMmNMy/Aug3Oq
2UGKCM6KPyNbscGKIjeME7kWgnUkWv7i+hLh8RLCbCrkDoD9z560MKz+3wnySAR6gy2mzCbmsjE7
rqwOpWzMF88Dvuzeq2KBW2nRY2JZ8Jyz05ZH8fJOXEZ2DyF3HdeCX873BGtsqj1xfWxRVXQjIyCA
xP+2RMvNErzJr//nSfuogRibBtAF6rCQ+c9cKs2rc3O1ZGHOaoy4Ba8v9DgC5yluUEor4CG9ZsvT
Lk84bOP7r43lFXgTy/Ll9TvsOxOMOuggDska+xSlh1QzO7iaLr/FAWjmZ1Mup8iwyftufze8eO5d
3u6lwHs0O7Lv0nkVjfVnjaNnbxy5oxr+ScLD5008NWtfEuSihsqb0R12F72upRXyh5Ivjd3Du4GR
BGDTniX1Nv1BlLQDlgW5kjUmaWn+uXt9wrJ57HlwYCIcXs1XEd0QqG+NPgCXPYFVtucIZmr4P164
FrOxA/suyEbWS/pu7A3puohlN1DnSGO/zh9zDTxqqXFAitkau5gK5OcE6838gBicaBFbChb5L6AS
ytFqtPzFYTkQi0lfVWdBbFd1zxs+hdlZ+/fgWp062mB43yyiG6RYHzdNzb7c2+eydMelnRaYahjh
pzDc4+bSGcZJcHlz6fg3uBfw6181vJ2KciJ7gGrcRsi4z80XPDXxJksU5GkXZnQ3ONtapi0nt9AY
gAcQJDpotknBZXCEiTFt6D58JWsk0ZiOZ0bxUxjQ1IDrtZmfdUe22hnmDfyPg/TNCekuksb7NL2k
W6iBHrN7gnjOvivplw6k6rREHfqooz0JO8l+4i42dSHHsXYudFN5exY5pqKRFfiv53EGpUireHBP
04lWJhwRvXOW1jBCGSWtLGuFXgsH0NYVYawKDVjpYn/RPWvUJlidb5CjubeOa25oY20aVcnqXMOL
bjIRqTULKes4J7NtcJmYo7bnC+0VfGq9fbpCWnvn9l9L+7IIF8Lun5IFLtBYr/LSEV2aLvkloMOo
QG98c/0L8OqJSMWvCAa5SP5+FdqKcdtJDYWGhkPjkNe5Dn7KXrWe89/NNSP1GlI134C9XK51gaTp
8e+fwJCgElWN+j08/N2Uf10LCKWjLHdQgFGEchSPg7j24s2mKY4yjRx8rTIKYHLL0Sk2mw2If2AW
495fzqTb7Tsk173BJ1Y3VAYFF48m/r09R1JUKbP7Xsbvx+34T37hufEZswa/XS6hC/5fvigGXzqg
oQDPW22LhIV+e+N+X4nllQxkhMvzBV6S9RJt/wKkkYoYjU+vM5hmgvotVsehke9+RfdLZRI9VImB
26fTNhlcky82tOhgQGXGrOQBSBWjC2K9lodxi9l8Q8o+dOErTRVPa5bA+cQ/WYCb4u9akYRCJNKe
Z+1daE6iMTmke9xFmtANW+t9nCvn4unNyz9qvwAMxqMtV6p7T4baHNlebT2L7lMAA7qYbhp66h9u
QB9iSRbh7LrNuNcYexmN9QfdBN4WEmlN5KvKw50kcwRvNr8mEYrABUh81PawuD3guKVOnNcSyXxE
7n8p6dbk24FNw6fTaMBR69U7yQVOAVfK54bEckFjMS0DGnf5sz2rFId8OwTMkrQ+PQrW9KfSGLIv
zZJ+Z5PXiq6YBJAGe+3f0X8cdu1j/SHPGGFWpmNZyPt+3SdKlac5bevkF6fnL1reV08E3jE2veD5
b+DYa/Q7tR60CQN144/hfbCintTLkwODd2VheBwZ6zBHSygPGBVn7qqBHalWLCQqlGB7xwefzzrw
fNsR6jooiJRNxY0A10OPcSY1NWJSay6S7J1Esb3xB4AHzoMymhY4NHUMz71oQYelVgVH1J9lr9mF
J1yo0Jp1ksaJwN1EzpF0IE6UfEgeHeISnLlYDD8G2W9ggCTNjPYkwl7c9iUzI+WwZZEGf0xzfX6E
c7rttzXG7VsrVz4GMqgq7kr4Kj2GPNXhr0toghvYTnoYr5iNY7LuEY5WkRgKvAbQi7x8RQaIdT5n
gjz6nk4Fa91wqnljcFnrOmQ+i1JL/J+X2+EMCK1F1SvHejb9P6v9AuWf2VRBiz/uGMsuZnn6Yrb6
KsVb7IsRtlDVznSdLGEyHlQ7vvw+3vna4uaClxrXEoGOQ2zQHVt3QkdBZDw+gbMK1oOobPCVs1gF
OhRRUIZp63fCoYN8ySO3GGg8f2SqWGHsp77NR153tK9tAWszWERUgzOGVTNEGlM8pebS4zDKx06N
C30ieAN8QD4xyXudcBmfqtb99Xmgi/N1R1iMW8NEkqBeuJ5Q+K/WADSEWBSGcER+80Qcu/Si3qyI
qEFWaD/SIO9GjMqofCxLBusYWxAa8VgD9vtcqxE8n5MdDZswJxTYH8dA33EF8TVsHiSMYM78b5ew
Bq3EPAGzJGelkqEjTTLsPBvDl9SrmvoqYHFZRbGW9ag8U+XpBwuIXrar8NQT/FOlUXIOen3ii+i8
JlqgnXsPGJ06T+VYL479TmIk5STOS6MJDO0ZTm8HJJpeQkf1lLYBChqhCbioCLjqW3VoIUuJZU/F
cifRFPpo2v31llwy8b+dxAW2hXkh76PiT7Ums+KuAHGUHyaPJMoHVUgMtO78Pkmlmr44bUeynHGH
mV3qVQfLgWrRxZESARO25EDYs86XDRoT29PNyl/OcXQGNWTTw4blzijYjinbqkGu4d3uR952dK1I
rS++cpVAj089kAcoF0O6eplWT3cbbilOSONaDk9KJrQS2Yp/KxQg2u/iB6vdeV1mbzrc95yIubSJ
SCaO371hELbuhRYTfwvTBUzlADonz6jfjfioiCTSXWJvwmwa/xo0yktDjPGv7ytdEk2yJgZmL4BM
g5MUmJAWYLglvBo7OjHP6Ak7xs2jVeMjbYgihteQlIIdvV2ZuX35Wb6hsve5QchUaKHPxEmd2Tjq
id0jZNtHhL2OxRIOvpOfH2Kitsq+zzQnwePrl3n559Q3ZM5gTmSlk33jKX3aRNLivA9lyN1M6SxN
TTZNgs+RP7nB19sShn0BuXR3eUeJRkKP6p1vfUqbv+ryWLjOkz3KjxBauir94Uo58bd2VeLRARam
GZIZ69L+UkssehhbYVOxWET+EVRy6IoZ+GBdssLAcQxGHU0WGkBszv5PWID5Ytzonlc2euQdX1D3
ipN66FrluGi1XHFOhl8HVM3YjtQJCZyJ3hWcWbNThcwNuW3l96FE0FB55Efjx6WB/qFx+680os3k
ak9xDzJ6W+kIJaiLvNdAdae7FqSER8KLGA4Cr8vQfKaYXWE4o8IB+FrAlIg2AYfw5QpnOl4tKLIw
tv7xSKvaiomOBvYb+/cuZFtjzveYb6gUyvXG2dei//LHdwEMaTKiyo7h4GPiqtVtgDXWTH/ydBCm
Ga13gOnyjxd0i2NAhntA04grZ+qpymFu3nCUMGrGA11wkDCHpWQTUrck96U6fvemKAQ5wUdyQKhx
26+LJ0JxNH3b2JfxJaH8nV1R7oGlzy7DoMMmmkICSEJptKQGWIH2PyLenRuLNbkiMMMqMexmFJF5
a0KnrvTFt7yN0w5k3Fm6vXVsl3hAtWEUehI6j8Srd2XtwQ/OkCyIuhvuBhk2YZ7CFwFj9mtemjHE
FZ20g5q8vi1HRPB8V1/h/ocCzZU1xmbKQV9DpMI+giGofEtUIyIH6Y8aViqAEIMEQIyBKRmt0+t6
LgD65p8Nt9gx5eIPILn0p11goy+CdcOQEDXncSaPLu+XRlyg5CJD7JOd2M17b/+0Gr1UznF2g5C/
8pWJYCdQD9Ol+yVHbbL/fl919SBzs0I1YAmyiTQyYdS30b5H121xhCD6nqq8aiaJIaTrDRL6TEpk
I8cLaDtzX384TFJOFCyTxtxuuaXb3W5lTH40T1Qf3drPWPsgTg5Z3wc+oNOIEun1YbPXvdFGMx30
84fDTvi5O+/LgXA7clPCvsGEvKiBFAf4/u2BV50cox0Zi+YXGmecEJi3QxsZ/pYPEmrGkH9o657p
QAFsPyt8Pi9ZnnzH+0DZkWNpBvPAjFob2Rz8JA6cMMXfRAEHQp0BgRKR7SWm9nSAhsY3JekJKoCh
aL5oJxDuh43G1AmuTrrbg6Sj2cP0zw8+E/EmoiPa7o2tywFrtRiSEMJsViob4LOOcNGPKZuOdly+
prgY7ew2t7WdBPjYSMZcpZUy3fDkcRxYf9TiClprp0JpnuS90/+XY6RYjVBoJrjyQJr0uLMGeQ3O
DQAwCJhmQv7TtINJe8O9rhNKJbs7Mcvo+PF1xuxbgHa3WN/bSgHEjhNZdvmejVpM5GLkKYTsS2/A
gDtAwMS1h96crcr2p14RNHGqerH4/Jbmia637Xvg28Cp7A74eTCmlIrN5ImgL4tpbbZhePyax6wi
/mxS27Kn42jNF9XZMw64z63qb6q9ZfYNXEepJFUDTd5cwwyil01lpD9+//qZtcmm3glu+nXpiEMl
caFNSrqi0deouTcuCf8Tt4HYnpDyLh92VixB/lCwtfsTagVyT+WgmCIov2haILw9g6Djm5eKo6Iy
cD/5MQDOlJdkum5CwYzSoJ4iQyGQOQbWJgZXsD/qDbp/qd+XmhCKPgKpqK/RemWW5Ytu5CJSE9Qb
XZF1LlIaorhIcOEfUlyIqoIb9G4omwtTSmoWI1h9qjJD55XbwiHv/+GdZbDOUahchrZBJmf72QyR
cnZXKFRDgAXBvsQTnmPQLRjQrGVW9JWZzYg/7FqCPaMBCTAZj7vlUH5EImcmJJY21GkYQRO3Cde2
hFo3cIsN1X4OLgJjWHWtgJTjzpMAwk86syH3OEbmvawTSVUCqZF8wDZ69/sRXtiltH3nEqszaz6E
6Ip1qrx1uDnOKsCaS6L8EZa1t9ehPV29kWN81pj96Zvp4vcUiDiF3BQlpBVUh6UZzUCfmcGiOIpG
y6xORar+1XAZB2X2MWs4sUfC3oIq51C9qddHniF2cPwBtZnjdhlbRqlCdxC5aqEv9hooPQZNU5ft
IPowylvvOPLyRY1kxrPq5sNCcrNbEZQyzmwjYid10wzVcQjqBjx9+dgvBABKX5LBf2X1n/njmpck
hhHDjaiLOJV68kvoLwSynwWRoPjQwCtX2B2Y95tuPfx3dkhcyKirBRiM4MpLFNOe41OvGhqDhwhz
EcxRiHqCt9l4o5lVWbLoIIJm03hvlo6y5SEOJ96zrgP4VbufnAvONWz7T4LfAoZEFBoVNDGYkWeX
44HT56ggjUptcVlnCRAfdN2bn0WzCrBl2ftuTToWkBdRskRmaDSgTiwgoNW4+JAROFxeI/nPkJWG
gQfsMtIPWYLUnc7nWnnH/GN5Zvufu2YrFMsoosVQtWGBpAcoE4GfpSI3EeTfuEeAmBgUS/voz9AK
AXbadINeFrCZvE1dyxtzfJUAInQP1Btytfov8uzx4Va0HNyKNVtg1nX2922fRN6IE4fAFtSfENbm
IepNNT3k2v+CuJ2S73pG8N/7tg4ctuae+16t0YYyS4S6439YpgowxA5esY+JxDSP9AgggWs4Elcj
roQLAKn0MFhOFf/Vj00umr6SVpBwMgZP6MU/QQx9oLQgFTpv8vOpHqD4dT/Bs/iMMAOFuSRF9Yfy
CzLqPSYKitC6NsUww4Tg9Z7XX4/LiO2tJ//e0zvRZKblwSsGGZF0mtjeQQQ0Yp9EjikzewowlvWB
1IA5FplwZ7TFRsw2vILcDEvZcDE/X4zG68i3rHEdcuKI0WdHLcBYyTL2GrInTGEHFWWxx5skzbp6
dGDovkFOXdOQwlkr0WC/sf5TH76fdWUY4A3fmbBB9l1xhlKVpfl+TlvjSDVcM06T3yB+FNCy9Tzq
MOlDnvidvFJBweadQnswQ+fEiKNVd+DzickctFbXsXCIaB9JGSlYsDbs2umEghYtgQ7HAaZMDWJr
GW5HS1Amx7uDfqR9+bO09YOx5vMdOrUWyXXm3JIoVsCd5Vw2/vpH8uJDfD986hgFcilZZtUu0psS
zg8K5HU3jNgH/Rfy0UlFIatBmV9/qAbW2RfbZa7FBZTtgx14BQjTnf0lDHWrAaw16UlXCVMFC1A9
+18RF3gxSXKLg8tks1JV8HPwVoFgEDsx8xKjcjhdXhuBF/536olU58lQ7YLT/0a+rhwZBz75IEVd
AtCigcIqXB5F3gKGALWufkehmMVwMxtUvMCuY4HM8njddem5gGt7dPokdnSrYgjS52Q67cp9enQt
hWUimbOGG2wkucGbdUlX/n1OvNPFQ+hL0gRgs81Kr5Co/GSYru4eZbkfCLgQddElsZVCtWJL5wNn
/Fr4uGMIy5AWFe0wzPoXcULiZmSHgKNyIpVJ4s28+LevhBsBro18lBZhoRq+3DcVvyrtydeEQkKp
7Kwg1Y62C5awZp/kXTUyT5Poopezw/Y1yrMvQEtJ7QBq4kh7rkgXw60CgZSyUXITmGIrT7jZEoOz
uvN6hH4gd8TznytDu1vjHlKmVX4m2E30GWokW11W6qA/VyGpUnZgUoS6ZjFPwtFbChq5gGtuegNm
83CcdE4u3Yn9xLopiuax9Ozcdt4yD2TCEOPRhGyv6dyF4vAyd+otjIA9CMcgpvero0yXEYsWk3MF
3yFwTDh9sMw9r5LU7kNyu+SeHLYNK5OqNW1qQi9OZvsB4OHybIWW8IhlF4/kEdhfp4m2ppSh5wV5
BR8C2V9FPY+eTANNm10NWXBP8/5/G5gn+3IqHNnc8xyeHGuZzBw4JwFKD3NICdKrVv7EObDpxXpx
VxgbfsTpybj/KYKwcrxMb4ECQ52YSZnUHE4Qo+IHQlS4PGEPiXDdMlaDEJR2OP0mmhQVF8u9TscG
SGiI2bWtqIoU2skachj46T1NY+Rzj2+aasPaLnIr3JN4PBvoRAv1DqCgPY9pfyuGrJsqFMnADomN
PBiAFADZWx+92DLb5w0J771bsE/Iag433pzYq1UXCi9oztIuGjqgLD4bTaOayAYW7D8Dw8w7l3Zn
DE/KWXRzAu9XH0eNvLea6LpLMfcVy9gieWqoTPG94nQaJavqiGRuTq219l/kIow6fERRMZPZwODp
iHxmBM12wCcUyIK8BNH6nBQruM5NqBW25LcOJZBkOSTfLJA/oQEMOiPu/wY8sNUI+SuQI0N10eEA
Qk/eOiL6w2eOKx00yOCVYeXtAOqMRjCSsTa4rSV/MNIgxaUG8RqkcZF59jbitFGKEtjMCQj15xJh
8zvvo1Oj+BLOwpLr+JYcifjgD+T2pFJZFQxWOW+3VK/EYhzpGRlsZJ4E+GPGVOOOv6S1WLIVdr9X
2ELZo8vXYRBmKTYBb/Pdp/tpaT2HlOfM+NgLXWkjGcfuPy1jRjNjDudkXNjAReFmHpQ1OMH4uGfY
23qu6FlEQ0baMQ7SC6gCmcnHjv2siZ0MOWdyrcyaWk0+BTtYOpRcuz3R2y1j6S641t+zXvBp/DWg
Ijv+Z43vsGij0p9wh01uhYuAefEI1PW05HDwsA7G979VZP4VbojjzLu93eY5iJ3Kg3Bytk7GoR+r
IIHL2M1vETRCaLaVaxlSNm/JhUwtArn9PmF0aONKtPy7GBTNnRrgCEPCZGMolNm8DGrbS0valRfi
V8qcdbuAfpzw2BRzU74r2vWXBB3WlCqGluZhk6VU6sGzExDSaRAPAG4oBrmt+KwH6JwqbbZx96xA
V/G0Qv7ayDYC6d8d3gRs+es2JLdrPCYLdxIpV36HXpWWB3cCYmNJpOKwkFxy4kv2fDxByc/h8K0E
mHYCHh/+gEgVNoprt9+YZE+DSf0ytvc5CKmxMI0jDrNT8WKOhZHVAd64s8h9DddS1iGYqNji59mi
RxxrBJnjV+4P42D2UFfT+0YaltSz4izTbW/sGGPy+Iq/hwIsdNqvLEJqtowkk4/z+z/RzgTRLZ2F
YgtB/fBZ644EWkNUFUHmdCKMO7PtAiY35rPtnrD/K93CQ6gd9IGFH8VbldyJV8bT5LCBCdHKqjui
2SZ4oRbh9C+JJ6+uAnEPKHtygdER7osKtg5KUd3CdfzHRaTFW3NCtWiRCaYLJmEXmrpcR4VK+wBA
FI+9PctYhEcPv/Qacnw6tgxGA8las+CkvsMWkImgDoVaV7fCrmij0lZpY4MhffobDPH4jz1xQIQx
XDgUjnGnUs1MsK8udtVzfxy0tzg8WLdeOyBT4Zmqy2ohVyGyy1J22S08erWGPUYvmCO09AetW0LK
9T3iEWni6YCd7TJVNkeAh1IxA/7Tnx4ms+A9R4+dlAb9HEDLhILV87GbFsBGfkl4OzvFRf95TBfx
PuWmx5qnS2JazFTOB8NzJaarSmr1Ywc1WHCadhiJPTKQdP9l+WwfRSdUtgWE4MVtFgiGrOj8QVIn
oN4xvdTk6gklK9Xc6oZYbcgSEiGPJOHpjBDwt1Xsc/5rpzZafnJe8rAGs64Zs9COrMc1cYeJ8JgU
a20ubY4CQkidMauyi545LguXHEPERxmUvqHjIhNCKEQ6qnEpZx0Tnq28bVDqoywcgUdhk+ogmbxe
Zc0NoGNOFox4/XhoEKTXuGClBi0ivhKIXxmxWNsE7AP/Y3ukTuUwbN0fvVSNfJrq61WedrU3xwB/
Ydm4AaVXKnLlsial6KJen6AVgUN3fA+LrMqi8dwUjKpTplk24ZYHI2VNPcIVRoXtXWOCNNwFZC60
yQbOvZKoCp9/y4zHmkF9YC+WhjUL6M2Hs5MRqmFOSk8+b2qXnHX7F7u39Absw/43E2vdCjM3lkyC
sCQAyTNo3vMWgF3D68YKqW3m2U8njDaCdH8ZcE//ND/7ev4Fhl2izy8uPt7itY51EWvx5X8KWAiW
Og6CZHAew1pD5bDfjGp8sxF3OptjHcIAWjSJSQKDluHsypEn+FDOQQhQJtWhtwBzn7IbCcagb6pj
qz3GDvfgQhg3Ne32/u4LGWNWydCVWmUUWqvvA0jLAhhxinNp+9r7FrQV9nKp9tc8UeQeWE4aQH87
oA2LxRTWfeUu827WVxrBMANSkP5PWoyNlffRT7GjqLPYkx/3Q+8iFvVtJySS4Q4eSeWfO6TOfB6W
2vResyer6BQU6zUs0uM/twT1OB+5/S3BMGdliwwLzlRkEtS7NMJ1XHgF4OrJ4qHuz9KAanepHGfi
DsFffFTuGbYjq1d457/iXMTRkrQNyC0beX2jiZ2nuMUALOB1SfcDc6jMBJat3foomiAkN7WG3MIm
UvgI6z1pJ7OFJLZbAZv1kyvrDdvfo4dPz8wySaCGwBGM6kMEJMZihWy7s/lBKJMSncS9RCShtbA0
ca/5S3CVV77IGlFRHscglUFCKDMnHV9EuMnooacdBYeZg5ZYeYlvfJim/M0XO9ClcGlHP0JHeSOv
48tio3vgsrbPbTJWDfCvjbyIgPfg2ia4rLuLRNpJuJKun1O8W0nTW8r2JNgiyZ9MaSIArJCLeSPb
WXZKxqU6KK3NN+gl6jAFjr5kbQtiZpuV4L+m9r6Q05HsFxYC39FikcVtL8cF9ZsmhMbs4XF+BbOf
Lq0WUZw0dvH9BoBDztzmePMeJRvvlNWAfm5piHJSLSvKcSbyycZ/uHY/7p/Ya8MQs6N7ti5Xwq7j
dSUoGgwxPZ4N7I5Id39qlvpQo2DCf+MIWQd1ofB1v6eir5zlOVLzsMSimJPsgJT8K8xXHKN5p/Kx
V11p63i85ECPt0+CEtG7EVWZ7DfsG9pMOAMEDsUif+9Dd6eaWtXT6dkdvA2W7vhoqNtfWIHKNHVx
JIIdVnXr5KpeTCNsZWcxOM6QarGl2Lq86iloapOfSiD1y/KXLo5VBN+kEoQR8ypslCEtxNgKsts0
xOumJ3oJA5cj7n1CYhLwrYrxox0W2Z10qpGqzITp5yLJV2qYCCRVgtFCOwEAbBr8KMIX6/ZiVjED
kOTd+cC7xbyT7ZhOVcYophSgaJQbi6PWH56D/occiBUcpb09ASbqWtgSXVVVDJAONELKVUIam90Z
m4wpGnFYua1MnUS0z4sFr5FJfLmF9HBRGpKX3JPZGIwF5xhkVcegF7MWaH2HQ0HZU1kXoe/IDIDW
IBw233mlGWAFB+UApdUJiExFoZw/FNkQBRptmLYD7IA6o8kzLXeiJFi9c3jRIdyRWpvmWRTNY0sp
petQxjuR4Vl/RJZG19z8HJOYHlaLm1jR11ilISyYCKU0gYxecUx+gEEJvh7P65hNTE9Jq8dYU/4P
QOJh05YMKurgZjqmxHGligReboPzQGBcd8VlD9VzIw92wLm3Dr2mhEfAkiOPdDAjEju6O5jYwm9B
rVT1Uvmbvdodo72avdaFoTWj0fB9oYgzDlcg35V9Wxvs/nUMqnUtgNERmqCcVh/IE3/U5jQnETNN
Bv0nyORD+WfBrax0y33slaQu7v7D/xZU32ItDUdYMSb3HAtsjZ6+81ON4kHWsLKDCn74/UKyw0dV
PkNznOZidJw4Rk607xTOm1+802CxSZDpht2y+T4zB+yEsAgHGA4ECFEUWDd9RuN+cSyjNCj6H54x
JVJmcm5gvCi0xrqPL+BrmO9zODxhoikm2BXnZKUe1qu90gDQLmhqFIJmgkG5+XG5SzgMt2qArwR7
oOB8r1XrbhAHvZPI88yzmLmU54YRXjdkwnY6ayt5bw5P6Z+GoW7AlymAWvGduvLUs/6sNKbvWHk2
gVypmqCzqJWodSBW3gw7PA+IsWln72+93yYJZ+Gf2qRC9h5rAx0zu93Z0nN0h/ApydgSaUXLSPrr
eWQuTHFa7W3uY/dlITq4MmvyhFt+qUrsk/dVP9AJpxf/xtqdhrsYSpzwVxqkEDhOIg1AZCFL8TTa
XrZRgh9sj4JisaF1tVqaYexaDeOyvO4ktdiWSz46GjRi484t1JQ3bq1PIl6gFXc7Rz9soVAyu/+B
JY5GqQyuarT8AV0zY8o1SYngmH4gNZCu26Rmx2KZFNWfz3z1GeGPmrlfiexaDVNtvTGwA127RrcA
g+NxQ0JHnztNJ+gag5WxADIzwAP72mqFG71gNDvK3gCYPbcR30bX1Ov+I914jUdej3peCsi2N7uD
MqN6bUVDyLDIzyw2o0kCPS7OO/yIHJW5mC+3kE8FShdo53ebqOgy7XO2x06q64Yy7vHPU75FB4uQ
UgB9WdjWhHdYytngt/R4aZvtBCEMP/2Cp744xbHdbVeB0S9RGk3KX2jUWtbsXxmGQwkqyutwZTn8
KTMb6HWKKTP4uA0VpQajCKA7Gopnoipr37oGUueyOEDfc378ykeiR6vAJPw6cb868boF9uztAWKS
P7yjQAaO849Sdya3cd9KVO0uwxh+k+ltAZyIwqJU/FnRMvjGdLX4Rh4uUALNsjUWVPZw8AXTOsou
YSGO7WmWdpPCRwCXEm4sedXLE1rQSiyqheT3qyhp3hSvoSwA/pZdDUf3RGzsbkKiCEwdCKiShDLr
TbPo/Gz9FEVTtFZLM7W5zu7O6F6gB+KbN5k8Ui9JADr0J7AcbHWeneXVMXSrsxDiDGxCpBafHXrk
GjoixppXd5YXVZi0HVGFeJepBbRYDRyvFPTII4mMom8vIh2xZKdgKRvqSu3AbomNhem3ycXRgbbE
SGb3scbazN4jTLk4FXMjACYc1xCOP/5r6Yc5bYfnkecQE8+ID/GT8zViIpmmg5c1Opwz5josFejg
1R+nKfUTMGxAnA0Xqf8bvYLpT2qCA/h41Y+adcre6xDw4F12fTNLZCu93kCmLcmVWGyK0kjjUWj0
S3TaJrjowsIg/7UKPOTXfEdLeQunFjy9nNfcJLGvxenHIXW4TjUVAuv1xnJt/D94BeDN7hoyt0an
003P3p/aneVt/U/FnAOziud45NIqCAIZ3iPVA0oHYq2n4gJpfmorcKd3IF4tBLsDylfEt41KVp4h
4Ufy3vZt4iRaavD6EKFABZeEycfdL3MHO1YORFtTcK8degeprWMAGM+ATEm7LpjVC8YyiZNubf84
7wlyofahX8nzuCiU1tu4oOA/TB4ErwsK6pdeybgb8mzQe39hQUyXP4+GdOSdQxVGhc7v1+OnpUBz
6LdrW/hUC3Z+zBWjSTk+26GzD+LYlGCRR583bEZMfKXBIFEKwNWOChINtXoSvI/lEolWWHOnMvPn
uPK4gMy67QytuuxcvAjR4raRzazOXC5c00M/RYtGKkcmr9oB86j+ZqarCaStWmhSQehZuo7BIeO3
3g60ozJ8Y8ih6EzVB6ce7Vsolqdrciq+7wBZ2rY+Vtug637UaYzT0UiREdWLo6pKTv8R5nur8w8H
P/wOj1nCLiXaZ82zngaYUhw4ARQEWr3rO3diPSJTYA5kyBcZmk7tiQNdUb7gmTjr3MCkDKfrrYBE
csBDNulqiFtZ/xS6m1hyMwSZXZyDqGizlg3g9OBu82mv+lVOY7PDnWTKgsvgr79JYeTaOHx12fTY
LYtSz3WUihaWWE299jKAE4fXcDosLN8lcA6peyTbsZiRANeaSh0nQBl129Uzd4s61IY5kTRRS9JR
DnHBs6oiNFbu3ATdxyeiEtjpcFX3ZpCyisVOY0s0FqNjZkVqOBjtPJfyPT8sF7ANtbJXNQIHltP8
Dqu2Mmutfy55dvtbSuIpt2ql8OCatqa9wWbrcG7BCdhYeEhHyFUut7zi7YNm8DTiEL5b37lhZFxP
Wv4H3DXVTrSv8jXJBheIn5s7XXLRHXCfNfm2de0m6f0B9yq0YCY6g7KeH0ES8/A0GW+H+t0XK1GQ
ChBVfKuXYrmF6qSoex68rCnDgVb6WP1ezmhx7XLb6J2nxYOc+2FzY+NrziOUX2Ppj9PZy8Eg68JX
wOqcdV4370X8L2W8pHc7kZEVkkauDDZhbqfjBxvihkq+QAlN2AffkoQLNdMKOwV2+MuJtylTWPYk
L4zyK9M9hqNZTqr/cyQ7YLWkIWTGhXANXC7IReaaollB+J+E/7mKg8+AJixlGPpFz7DzX0TfYO/2
sapW9xkkmyPJESCP+uTqvpHD6nS15uo+ItfvzxitrC5At3e52PzrTor9hi55zYOu1bI4YIDSJthJ
eXFgSqkyx+wV+woTQLdCdfNUWKo34PcVeCXddTo9upTD1HTQdlwEMURXHj3dMU5lhwa6xfvyEzzc
+JAb2dTqRcQCQqCDJ9zX0l4ju4gYk18mTEGVi9eUkOj+eTXLgRfLWomn0j5jroizTrd/1JIKN6p1
a0qqxjn/MJ5sUdCC3Wz2j8zidzak7xxjbowzsG1K8lD2UzvUaUdwS08rpa23RxgHOmiuTD0SlVEb
GnlsT3xmoVSdusWGoObGlDMlafkrtL6MlR2cPYL8X9LXKZHXaAhJDQmlAykiV4JKa1nawJ7gpbrv
j5RPuoZ7Wqel5bJEK84scAZ3P19alUzSpeDVusRmi58xGXlgiMNXYb2mLC6dI4d0TAppU6w2+6At
yQyZ/gUWr/NhQSAYgOLQ1xIGbKL8mGxnVOftdKxp+rPADR4av2xKnl4KX8Ty+2xPr2BoKJTXGlXN
jBggPIiT1AJOI8LnUmd2GnxZpqp4GWi73JyRApJ0aN3e3Ec0DqU3zkJUmwxEqq9sOHqEZPMk5AA4
CVASUXzZJSkPGMs+uV3zfARPAqbHuPgPd9xi0JJQ2YK5RkgBIMgsEf+MVnr2UkFY9u40LxrF2wtJ
a/oXrLjoWvK7aJkOC+8e0pZifbPsewXnhizGVzNJ9tYmMLqCN7f+Gu/WNe4xgs66d2RoI9x6PgEq
iOBX9uEoQedOc82OejuMOPiUFxTs745XFvUrwWaQtcMHuribpdoZfmVy5ZU7rZH1tyjNUvKI+aiL
iQOKO0VQizFKk8C4VDIQRO+sI1M4phppfUBoqn9OKb/h/2MlHWoa2s1QL13tfHUt2js8pxSDsvpX
sYna52CZodXQiVKsGQuo77ryL6W1yJheKzbRTl5p9V3i5pr2sb+LU4c80/9Xrx5Rh0UslD35/rqT
fzw44ZuX0PznKm/XG2XPzCnAh1HzXtvbQD2buP+uFxET1cYFjPxfPNbCpZiU47RG2h+NrK8641KU
qK50X9dHza81Gndik5nHD2bGLwmU7RLuQDq34+bEa87YyP7LmB9SBW5rqlvSdTOfHL0WDk3mjEyJ
jNrMyZh75ABzMpKPSCH3T6BH7ArEb543Gfjl8O1adKSs0Xw4X4gKsDu8hQ3z89uodUETCHix+8jr
pdXlxZ9xy2JFHp9gco+xPrW5m0EosWrcB6EzM34RVFpBbkQnyx/VE0Wh5huMg3x2Lt9NSiPYpwQD
ctySTqVpL9kIb03GF895NCJL2lURjsYkreOscLPm3K0+3HYilVZHVu2pfhQRSKX6QrVNOdmuc7UF
gmog/o5TDkMunm5HAXbvqsWXJQJaYHIheQ0CSnO1mqE1jpBz9PYTbp/BnL59ObsOPklNsC/qGnhz
4OMCH3cKPqLgMm5aDFtw8B9PFXXoJN7w8LCuT4h3iqOKpMrwgJk0ouv2AUSPquhYR20+IrLMv7f3
AfOc/r4p7Vm89hWF+FOTEZ1jbf3D0+CrIPSSaRzLIp1+f8Ltv5xjGB9wNIpIMYhj7gB+hhT7lk3x
VhyuQEzVz8YQXuSkXVuOLizV/WT2s8jZwNytIGfwSiL0/MktxhgOjiI1XZmmSOlE5iTYzZvibq2N
7/iy8jgr51IJtV1xR2RKY41qAWO6KT9ghcQ465yuo1QIj5JjDWwgZZBiyhS2E00lFvwn8eNa+KkL
dAN7K9qcN0R2ZCX8Yy5RNWKTJD+Cahpa4T+ZBtn80T4cIzzSNbfnO3bMkwxAs1qjV2b36pN7l2Vj
inqglSqiS6TQCfo9QatOqRgfw3bo1m7e2vEZdgLJRAdqDE2OmBjt+Ll9o6FMg2z/o6vGluUFCju0
AYd58w8gMYopy7/mK29AGuYjQo0KPd5Llv2kbXAONRm8LZkxz1h472cxUpzmItUHbcRgpEHHlCfi
8lqWEa60TWeeulPhDm0LtLgDPHoakttrqxjnXy+thrW3pvL+gS6Uv242ih5dQuXELdIeW1Fn4St7
rZvMzVBzbIceIc2GalUQIXkM8DWU8iownnUE1kGILABFJgsnKULwENRn5zwfK2+mhaJ17c8vBjSU
VxtlEIRcTjXwSInjJIpJPFcVYd1AD5SSBO2c2riQ556/GwdYu9UvlNfMdScpkJkewnIVHCRlGxwE
C9zf4S6JKkvgsBXn+WEyd4qZbhuwG0XgwMWDmX5uYzic7MZH2DV2eshxQL/YRzkVK10rGdTECY+F
ts1gFwrKrWaX3NgIlbwpxpq1EOpA8fj2kIl+Wb+ilKRvf+PXlpg0Hz9pSXZQnbACmdq9Y+P9XtgE
t1Xpqv4QmlrK9S6Z7ktZWvs4PNOsUkJD31Td9VDU2ma18+yqngF0+wunO6bXgFgULwzP1DMlcZ0R
Ahu3wfJK1w97uht1n5fIrWjulMWvyV/RKL4n1m95WxcNOmtLtzXbX/FRo3hnRrPb+jyM6sWonO2p
f2PDC/B+sD4HoS4JMtUfGpsfozCTqDLjMsfHcHvOx/7PhB2y3DvfRjLxLTobJlOywUYehmVwX2ty
yqJoJecXIUHxR3V6oXzjQvKjZSiKZkTBFmC4ezX8oHvgSZxdNnJ7PVSOkW2ygqE1COOXPE6yKiEd
D1c/bZZwBslrLt6dgCeDDW4g8LYCqx+CUDwhpxC4KmoVT3GAwZY0qCXqQbjF/ghmqDT1ZHJn8vdU
nv+76tuzpVfgxfd1Wp1yJ1viilQKvZkW+H0d0oxP6De2AxYGH5VN3cucLIHE78mF8vafVHEC2bXX
ntIgohOaQP5Ai3vdY7ycKAn4O9JIVrySJztb4dzIQPz0pGkQVUsZHRp7BaUCtpvfJmKMX4btEd6N
IiYlQ2Y9DFTYLLyrGNvFpbgEbUFOr++XCauIotx0BbDyhrcXn+X3pvKycQbAG1LkROjOYebx9u8k
Yx4IUQKLSbIKLrcOBirei978yYbyM37sTKkYQ6LAsgxA2F1+1KEpwGIvcxoGZniCiiHaW6rayzRo
wU0XM7pWIc4vMkjW+ahnSzSt+iQdQ9erwsUtsPoEXKsqSLEBRNFLJnJOGqSzSYf631RwtDmErMgT
F+3xlFghEu0XQDlKau7ewB3an2UpfW39Pc9SxpYidkaVpXRMbGgGbJRuQp8bAbK0cuuwtwoJQ2M9
urftUZxsrens96+H9JT+FYzMrnWJG2hE8liWmVdVco16l8pRG+mBuXFzLYI8HhfHVhgy+xs1QmHj
iotYAB1GNkiGftpYrPE4otXG7iTUb+Ri6O9agLthhQjhXw1PiwDRe5Vwcdtl4UCX/Fic6gPeKQpr
qOaSfNGXcAtQQqyaiUm9v5zR00VYTnCFLfKxB9cQIpbC1c0duMXUv8gynd0749xH1jh9nugmUHgE
A62wXFvgq2+d4DlnNFUuHKQVsNs0hCe+ihPBCViodjoTP0sstngNT3nto+pIIAYljXY14MTykQTU
DglsQcygbTagqSFDKzQ2rKKI30OddWxQUsApeTcatwv1EyY5AXstAsnruRO8PQ/SE8nIcNdLe3WT
JN2bnFVfjyaH1XjGbptXcg/WBZ9oSajVsyr6ykbW5/eySV1xm+AjAweUFR3pYKetpyOWMbH7JUrW
peZzDSAOOJI/2leBVNEMWDe/OY4tYGyyqOXdlKbfkbIEm19860PK82pKmQSTTpWfUWe7fxex9/OD
XdkzGWaiT5daDvqGrCtOKYQR/2Jf262vpFexuJaFqG/9vFnh5YDZOL99Kg/htLgmWiIPdPM1OTyP
Wso/1iTM4AYUzyf/PsGtKfKbWZwFzuujZoLZJVhhx3BRfj7wwusbeC2KEl7q8prlkMk5Bk3LfbqR
FBIQigWJNLi2WSRE8LrdW12lvvoVu1L9osmZQWGd6nVD7NwjYwcVEyDWT45f0MOEWJYerK+L0lAm
TRXewQFGt2AyAAJHeGMY4n0IN7NfnhgzsjgiROB+WNyEeo3ofAXpbsBmo2s2SdvXWpQLU8kPtzeg
iko/V5ApUIV9WGAwmfodZ99/VFyVrEQu1mhmxUQnQgtAmMLFxim49lMQTsdaE3pfawRzM+VN2HOK
8HUUqR6J15LfYU/Fc4zhpBs2rVYVhruge0mmR8u6+LutZ1M/aMXiYxwse97dJudlgxWyX43i8Gjq
7XeBgBfvpu1a6lPPQoRP0cNjBHI4tp2UvApGAChLQZsrzWeuK6ci/B1qwQsnsCFQPhLw32SP2Zd5
g17SQU0Ll34ZNfl1NjdHTG0m7Xc0yu2dp6OTaf0Zpfvx39i4NaqwmgTshDrbZhvM+T89kJfJmAxb
gnLwXmnNHnAylEeQQp8fxi5W/bSnidf5PKxQjXcszxNPBHXW5wDDbpY1LFEOMQ5sRKdzC4DjEUys
o+ZlichVdNdAe6ur04khkHAmw/1MT8WEJ9wN55Cx9aRxaty/tCRemoLbNNZCbPA1WK2Xdyin+UCy
rBJhrYhlOuZpsKwjdX/ajcqkI41nQ3RKmjp6K2O4yfrjiE+gBILsEolUduNcuM7XGCR+oWZ1Lowy
XaGzeieNXXsivE8jkuIrIoMDWEdOAXPX3MB/+ZBbTerw9ml9+DDttyR/20J+/0HTe0AicakJEOPD
bLedbxwwUrIGpfM9kr7quzXzuNEgoqx+7jCHpofQxSaZXpmCJcdww4U8XzY1yD/PsYicWcznP7YX
iQ6Z1AqioGioYDHz7jMg7NBBvmL1HV9mEPks5OD1S+ccTPyLGOBWGAmU7/CWzdnfwoSxIAr9xjT/
fXYwla3DO0fZWa7NgoLwsC/XS5n5cufPdQwfjJn+P3ozSrbRGtB9EknuFXTnfXn25Nr8OqweCdOo
BkAsrXEqT6Y6dfhAoCpz8oANcju1L0+lqUxd3g16DnH3xbmY8XrTpjDAohK8UixQPShjw0xcc19m
dW6gM0Nk+cHzABZOtguXsIjYpDtivOm+Hza0wXCvI6J3p6M5g8CB+A99JcN6Yc1dWQMKhfCb9kZd
4hX7ld9flhcBqKMO3ypAR0DgOJ8Ftw+H4jIYk5eVZD70J5C9dTCL4V31lvoviQKNtogTil0TbxmS
bMn2a6U4zRguCHfUMOtcfE/ijTEGzQRncCUXM9LOy3uCN+pRY0lBePWOgEG/yvAjwfQ3/MYxVueS
wJ/bONCCa28Ublze9U3YLAokfUrP4RM8I+CD8+Z9ep41I11fjYPegWGtHre1RGqgdpdst9YpK2VD
aBBg11F8WKTggAGCNBeJohYoQgmxwNquIOhQciOQsxeYLUP3AyNobkyctg/3vkQZbEUY14eXN/p9
bU8dhG3nlGQ04qxpgx6cmVHiRbgtr3gJ/S6oVwT01foZqczJOmfhLsWrz254mqIkXEUyI6wD1qOF
+X2Qj5NAtkQfimxc/qIq4kY5fvDqhbsFGDBD+CKJs035NvBSc0z+UXYQYixid5auSJcScCclYQhI
k5vOCzSSbZ3g8xPOAnrtjJ3O6yTW+7pFZ4BaydJIrNH6FO8/g1IYfAcgYhDZbUymPqUxtTEXlTAV
VGNzQF/V8KFc5Ojg9jTUtS6DYUq3+4MeCcLkImHIIsfVn8VdSpkPgeDy+aZAhf/i4XKv52anWBOX
+BbpJiMabg3aaQhfq0FuOCVbHSrCOxcTR8VLtM/i8gqPmEcgiutNVQJqs1jqCOeAarVbfXSAevUu
fCeI7qDOyk9f26T5jcMFtGPsVSLpa0OIRmFjQdpsQIuAG9aqGOJYcKDz8+ECE9nPX9xuqDKCmSBJ
yrBqUWYb1muPc/KqyZ7nY/Xt1vFVrq3DGAD5SDrseAXQ9KbIRVzgnz/R0I1FZECHVjwrjHdDK0hj
HhH/RcPMIDmv/JMKhuGrO2Di6F/UFceZBmRYM6ORaSckShGFJX3lyDMPozLe4mnnJbsH0ubDHg2o
Xqh4DBbbRXu7Qgs0ybc+QTJA3dRuFLrY9oGRJhe49TpiI2eAovO0W7jAi3QN4D3+tK24MHiB1EAN
fPlVKMMLU6PbCbcmJCwLoWDBS3rp5yJ984gSwNGEWkgMBUse54nRcBatXJxEySllhuqk9/wr9CAY
TWSuKjI4Ko68SJ3iWMgNvzOVfR859iwlDuGDrrNtFmdsoVC0LpoK0H8g/eu0oRneI61gRsElem7J
twZjXUSFL2VJJcDNP6xa04z1jN4l7UlfuoEeRweUzWMessJ9V6wST61jEDNvUfoI+0az2VYcxNIO
oIxj+sM6pb+yBPRfTJISV3YfBYGikWt7rYe7Y2Rf/HTzNHJ3wl+b9dwM5YJDpKRo7jiURElG+dla
FeQA4Y4NzmLd8HmG73LfHaNIfWVFnpk+AkprUpkWMNR9d2mMO3Iwco36PsY4nUtb+1dbL5aM0dbz
kEywQrkmAn9uN8o2OxBQPIae3WXYsa5PD4tIVpqsGim24bIyWa+JomVUIZlr7gKQqEm+x1gOco8q
bXJt3uajf6DhLJztSquNpGkAXXZD9dFSLvCQoGwVpGQduRwBvBmt6RPvURLEjIaWFT0bBVXvrYgS
CfB/nBdD4tZ1cwufik6LglbkFBn8nrp34BXZVcDtJRbRPn5qzpMw8d3lPLzbISMCrpNQ7ZfenusE
MyE9iomXWrUEOxGFDustR84gEWJhSDXy4/uqf8JZkRUxFBP3e48sgQnkXFs8dFLSuCZsw32TWyG1
o0KtSHWjM8bOVNyViVkgw2uT2fIQLwuCR6NEW1kdU41Wn/pRKSuPoazm8/yhZXrPHVjfnGWzxW0z
qj5iEH9RnsQQUiB51N8kAyILYOgLYifd8ovXRxBZGe87HladkxAVdrum1ciVT0w15GjxtmewQwLh
7o7BxOFAHcrc1sY9sCYiwr3s6VByaY3ZjZ3hB/hz0mt0+W0dNHK0Mld7VaX05pbRvy0juIHuYSnb
2JLR9FcA9hrYRPKHqGMzPrw9Q3sD6YRJvhftt4wtLeHrsXkf5CI1AeyE1ipn1ldVEIc6Vh+habCL
oHB9UiODma9V2HzNoVCz2t6K6mguwg5yPUO3/Y5HknxQsv//JtQIGtFspP7vZKazFqtthvCMh1CM
f9oxJKbf5js9Ufzs229YqWNOaXuEmVq2jpMw79WfnL9TgTxfwN7eFEq0qhkUBWOZZkH7pnZcJgNT
5KVzudaVxF0RkQrz4EpnsKo9IRZnOVaT5M+xrjV2u8gBzjwShefrCIv4ZJT/glCW9eiqf8tDCeQ+
4tdUAvP1tkXhwz06qIXY5tZRJDZd7gpptjp7b9sHPEKnXC3oVpof9/d9H2DUzGTNBRZa7+RRLZVG
35v74boHWSAx+LOewAbdhpwr8pWBEegKtMZyg5xRRYLZJzr0bdlaKXLbcwkVkngxXv49KeA3160n
yXtML3f5id74vkoYNPZabemdmsZeGYC5pehiaJOtU4e4G6hnQ9P2xGYTwFyNMnp98CeP4+VkxBbM
/qCAQYcbAGkFhXC0vxxA3YwCKdDZzTgB5DLRyrUmCycwPeht5Ne2ZUzgbX918+183AykNY3wnMo9
H91vJEkseUBPo0b778/ERp+k5NAWLnl167/IeTWXHnFJAVrE7GlGcoMI10LSLvlkiHcCrLRuVn/O
5rBvYc8EDI0RzyfBiNNMAFvnLV27q672VO/0CMI2htTwbyoLOCcaEq/QsgZ4j4adbYqxD8m97ebJ
uO44h3VhHSGD5SVC9wznVuMtd6wwQMLLT+7eqZW77fkPwJpYhyxgfiyweKg4WKfgCeot/j51X0rQ
YhlXzEFVsk9WeLU2H8qSp681qUoJUeLvcJdiORg09xR6hdtqXwjs+cvgJLJuv9WrFXo5K0/XcjZP
1QSlbMCAWzShGrAW6LZzc0ntovhPxq5R/Zsw3ccrglnL9WfTyzAssuy1a4Etap9vUjAe10ALZ+6d
vp030pHBLeIaGbb5BNqMYqXaGPRFfNuATL2PXBt3hvMM7z0ezpPhOHurJnh7vkKrxFOQnqkThjn2
Lvc7xmTG+oQLb5j4I0WI2pQLXZ7JubWQgMGvwHPWS2PRn5B30zV3WkoeDITWW501IJlQTnCHpcv+
/hP2SiTRsnNmOIY8fBx5tCB71dkOtxlj81Fc1xiXPJADEkAi7Yzc4lFgn+gIVm5VDR1jM8F9PpTV
32bR8KcjGZErKUntcjrKyKv5Dws2Yurj4pvlR7bMXL212h7RB+RYgHUsjfoD+islB3kl0TD+hV4V
cPYSM0mBPWhOHn2q+DkPFPsNX/K4S9neVjxznJJ8MkA22DPUPIVHEcG3SNxMs+debE7A9smJ9dH8
uJgL22JwN8f8cJ+gwOy/fwgIl0CkZs4VCoSwVDZn5QsbnhyKkl0YKpD/mU4OkU7G7LU3zvkVyasF
HU/1DCX8hB6FWolGvS5cMAgfU0kih9dXR+Y22iZKl+jeF00RlKhJZjYzDkpD/+VP0werVe5DQZ6O
nlazMoDqVSJgMFff3pQuRas7uemOxkhqasv3SpRzXODuRruBl93DrdN3jd3Q/GTz7+c6LpD7yWwp
w0eVTnsg8XRuO433Cak9TyHx2qkuqBv7BuqVBYmF29H1cEA3Kq7d6P6NH1mbXj3qHzOUZhcTERht
ZEF82BaV8CAbh3NEbd4ANNpgPEfUmKw/Z4fxL3O/ajEDnS4b8P+Ei2ZxOJsVDFRirw/oP6pHMgDj
hl9GtwEmUrFy5vOHyW/2/ZhFrw3JqCydv0aC0K5VXOFjxe8RGkPpqwjGEHTB+JOVrbTEOPb8P5OA
4/Cn47bFPNdli/ctd8elUjOyHE40Sb90449kTUPjHLU7ME1sFpV+y+8SLsUrDhsEzssVLH4lGYSC
kIFsdaQ0qC0Sy9cT5UXrXdF/di6e5VgfKv4FPxTJtZMGYlmbQOImzx1PQmUeQYU7vCqjo9IkF3Rt
L5mkd4SaT3N1PSjoG1s6CrkfpEg+1JWViKr+RDDfyTXoC1WkJJ7QRAkvP88iPYyVKNrvaGWKy6eo
xX8ZIhmAYLGzPqtoTF9K55Foji2i7Jk8gMkyTTYRitMhLUgtX2x+tEF4M4IBsbY7OB1kMRxjJ393
QBkIyTKn9ia5HF4JUTFv5Y5XXWbWgPfWUVKuKgHIEsx+lFs7sjby7BxWUxZpPtR4cYNfw/Kgj46O
4zMhpGbjZm9D2nDvJYgnLD/ews1RGs9xrPgT94uPvrX+yv+IYPuaVroGoBI0oy+aAV3aaPX/iLXG
pLDrVf4Le6thXUcPCt0u9jKHiWsH3mbC0kfeohu7S9WM4ktH8oDmI8bLO0Fwl0v4vH8TjYLySaVA
B3I2vjMbiT4iZyG4KaE+YOu+UUJhVmHNrQ76c0AKnfVMtwS9yJ4cEDITP1InpXHJCY8XP3iFawqe
9eM9LTPvSHT5haKs/yzMu8L4xV8rzvPndQUGYat7DeKI+FbzKQ7rrggperCRLlIhmzQetM1gVROH
BioJ40RjaJCaip1DO6NePu9rA5QZtovj09gYAY67dy+r3m+rw5htkVCHhxgvvNimtnb2kwpgfVPJ
RVI7yvTvFeASUvb1eD9hQJJdN3CmTM+R7/ffdqkGgppA/rLeqwxJYDQHFaRjd6+9R3Jk+NEctQLt
gYFehnHLkPdTbGTdR0PCY5mDZNoGI9psNovZJXNeves3Kk1Mc1W9BQy/XpSyIzFbnYmy/WCWLMlE
BKgGwQCL4YjrIw+DV3kkZe9fNmlusRHjDqR/5hPLrUgGD2fwTM4qbeal2p62amUd7IsjCgrN3QUQ
PaJMZVPmXUJRVRH4tDXq+fA0cBvwXlgY9pnn1bUnPZZtt9FrPkTE804dMNmm0Nel5FknLENP6aPO
yiHY0Yeuh7o18ovYfvbJs5uajcZSCWybrmCeImMeBl1vcpVgidLjXxEUoPmG3Pl63+Hi5Q0EeiCq
/c+iR3bIR0zoPOd+tY7IirA3ftFIwiR6SxYpyGQM9sG6li1QfUIs2hJDZLluvjx/oOnUvNhRIolV
4b3dXAawsWy+cw+6zH6L5yy3AcIhX/Po08TpfuaWSf4Shecw2V9IJBry+EHj4o3+q64Bs1EsBzeV
hrkOgdtmIb1WIvDs5cpq+meW7jQ/wEKeq+GWFY/vJRBPeFQqotgm3GdZJJGBSKbAoXFI8OTgaXPn
ogSLQ59sUjl2Ik4zrp2nbdwnAdQdMKRhH9V7niLR5r71Bq98WAQ8T/4cHY5bCiiEYsvwWH09IvwO
fmh+lla4qTsqsSChYMLg31c6CzHAc+2fJ8J1xCbKCFHGA6jAWbl9O2IfKSC2x567QFGCiDSXOHjB
LwA5FZJNBdiqbzOsBCAqB+3E6esMDxhiLdCyy4ae6Hw27IKpCOuatvzTgsaY+BvebMjT0lWrH9qh
XToxA/Zf91lqwMvnO7WDmGOXSzA5mPYzXI7LzJIydSMKZ0S4a7Ybq/ubamNewsnAtbP2A08VSPFs
E/e0JOBTK3tR3D180gVioHw1QETT7mZaYyFuAUI9K/crd/qPS344y6BRjgAS9hFypC4SpkDlDHfm
BXHg2X8D5+2rS9980Zf9tLqG2srBIjYXP2ZLXBMxmvikdmwaS8W1z1PhctvAOGRa3HKEa17TJDo5
KnlBNF5yR++Wqye5G8w9MXgcfPo3Lg+cxoupaEetWteE4zFNwPS6OZF6zvCoQP5NA0dVuJb7bn7A
fJM8GG8mdUghOK12SMIKhpHd82fsmaGxNvLiu58i6rcnfdWxnVEkq/KdrM7TSR6FYjEUVkuGTzQJ
vFqw4gw2SHq8ua03FH7KOUuhKuFqilWCWH66zh3eBRi54QXLizOauJlVKJ4o6Dj0ll0U/D7BmR9r
JzUoVPVs6Xaxtysk2tuQb4D+JPp2UBeYbGPX3YHsWzHsedXbXs0FH8zxXjVIAD8y90RxYZDV1M72
61GyReqLJJ88vgphhTFOuDBw2/f5Umm4/04T72uNqlwmo2BCv+vpljbD+af6f7XXVFSYCG6JPXak
vZA2yWrKDvywa+Fx2DkdicMmm7GqjZSJH+Hox5xpAjkZk6crZ7dxD3i6Ojm/Kcvgsw8ceU4xHz5e
rOZYBvFa2PkmXtbfZ0jCI2SQ+MekfcQCOrrGX2pTH1qYmg8VrCsF3PsRN82EOjiyAuBilow/HlVX
D+9ilu3TJdZ1wmT5nB+XLqLtAiDReBJEJmax+cqs5axEbqGvibw9sLes/bpPt41DfHc21/h1QMU8
ptgqHLlSbcB5C8exLFBQwLVOMhFdxbREMPUrt2k+FFbbspvYPDLGzE2WHPc46b6+zAix2WTkFj4J
B70E8fpSWnrNi+og0mj0u3IO+oy/Q36J8GiZDsZY34Qw36MUG0t7UMFQXBT+PGbBrTRwXi/sG4zd
051aSwRiiGj8YuALhMyfBSLKKxXtQe9CRAxY1djIdrZ9H+DVDAjhaqjeno+KWj4AMRaiUxZ4C8Qa
Obz/WIFykQ0XmV/fNdtEnIFiKbsYcxja6skdSSdMmrlAAOviigx9XeNPfC8cDlK+PKcpAc1bE1rp
+aHXMtKTtlD+Cya3rEe4w6aAmM4IDu1llMn8ILxxP5PAhkgN+hbT3pxB65BQwvZ/tSgIqvk+Aka4
kTJgP0ONAX+Vx5YwM+prpvZkNQWS5n36s4OjrJ8cyuSFbpb+qQDD/vOLk0AVeNGwbQRZyFRnkuVH
xdB/n/MgjKOFsNzM3DKVpFMYvu0zN++aADeQw9H4W6lzDHrhgIU5vRoPD2yEzQ+XNqfgeRBHCKHW
WcFwMEns1aT/6EuY7i7lPXGDnzkLDgFJjHdmFFseTBvq/DKCBIOGb9cauUc8rgVBEWZpFWiuV/hP
BkC4IuShhegC36VCdygeVg8y74UIk4aYh+7aisnZ+WPoeNkz88TsGi2zeB4H1ib+RgPYbkVzMs7P
XQON0EaUKkVQBw7StSRw/ZkbFoBnHy5D4/L+uoVG4qMLKQ3i6z3JiVn+umSa2np/+Xv5ESIR5ftO
kICv+Yhg2DWpdi4FgcDJ9VrOAzpXrNsgFUPfUi+fN87a2dQNafe6Oo6fVa8ePKrpJnUgYZxUJH2T
6TiCmzqi36hFF1Qcl2cHrEIm/itRwaA63r5o5avqHg4WDpMhYSo0wN1qNK2N6xhIJHMiwpQLj3lN
T6mg7okN+8vtoRyBtTgITzGf7xOj/NotUvfOcxROVWLnjJfadCjXKINlpLg3ZuVh1Bo0DagY03Vg
0/w0jyapXjuI8JNH+6xH58LzsrKHnNE160aE0K92qNOvfukAJNauHxAZtL26+/rmVYoNa7/3ma7x
VM8fZO/LfNuzUi93Yw+QqloqYWuclsTIb2kq2oPoOgq6QE/zrdPj4RDBaO6y/lW0fq+ofazK3Nh8
EIo9UQtgVJlrrbR5cX50UKHvgubXlS/WSFduKHAS/LwE01bbeNVZqFWHPQhRXf4dhJlAk63Yneme
8R/BQv6K2eROwFh9hPRK3ET2Zms4x0MUVTVZaIQQxjixz2GP7+pUrochn6Aa0qShjgDKOEGdtMiy
YuMxiwYvb4X1UyfzvtDSN67bCvVqywWeAoTwK/GW/aYMsyUQbGJjoiT7g+RxD7sAbBBFSkOCvJ3b
Fac6qqtma0WrftIU52dlp8dZftzBr0uq3ZC+NJC92fk3mkNjVvIcSQp+xEf10/5qAXCgQWCj8CS+
qfj8OV5LlYRroPrILFDFlxnu0fRXEtG9YlSBktQVKyAOG//i41CUnbmVTj1S2GmtBhPlEvBNZnuO
WAe6+MKaBrsdz2WWijjiqLXrOC1i9/lTInOeBEWomaRoxylSTgIsCq7Qfuk+Lh8VS4uIh+Eg3oUs
WaBRBDiAramxzWv++/3fHQj5VBB5P/QSgVpRn5y+6sQRGFxK1Mwr3/alusgkU9i1lf5/MC2sCYkT
UtB+mmisxQVZrY+QFD3J23krhIsiIVaiDNnEuW2y45QnhUDMNQcte2KNbNoDyqNBMbwukHuvKLHL
6FDxf/e9i2bapvDETV7mXAc4+sBLIUeJaEDUtd8Im1eIet+g60roYHA9D40ObLq6VPYhdYl53aZX
cqV2ydirdoHDqXx+EOqw7l75i3ZYzuXVgFCTVG55edjGySkZmm2NjVLLAkmqsFjNZrJxCwDf49qW
RwQiCmR29vV9WPZZtdzJ6qn52vg03VL+KNuTjc98tthS9nuM8e0YrvsPMAn89QUgDuUoB9Z915Gw
XWtClPDXwq/0OUi3C4Zqtb2bY61ihUU76sB3tk0NGLPQ8Gd1qqGzFWOhY0c4v51jt+JOIZWHdTzb
kCfyTFIXSsXtm3sHS1e8Yv99Y8JqAIHyue3/lE+iZD/dntO/ogTjgj/rH+jUB8kBYTWWbYGFBkam
dS8XZ9D5p7Mp0/KtV4QcJBka2K23rhKYQxmFnLtdqirXJ9/Cn9UpQV3rWodYsptoCaBFkatO2/n1
ih5qrkOREa4a+1xOauZv9io64+P87Xc//LSjFf5kdHh0kgP8EoFcACy9htP5LfckAJ7aiNUGpYBj
cccGZltcFFsDif4joh8JXTLOdeQy2v0JzR+ZGcnSZ2RcL6UPp7n2xUrLcZ8c1nn1R7EvXFvTfC3A
Yp8BSRGuukslH28tyWo6mauWnOrD4VWrsuKi6dYbpTvpV0VIIklX/kjAedcZ8OrzJajDMVfrq86x
IOHuft3DOvAvMGfmed4Xv4+83UY4tQ+8iwtEab3xd/I3KsDd9paXmwAQZuna1xw2+iWT0lyutFBt
2wGn3dSDu7RbR3PQtDP6PiptF9zQ+gXzPWuGvymd2Up6slyFjj5oHWKjC0CXEZ+6ZEzA4L2RvoUy
DtCZcIz5C2I0p63ZOtOKTn9HYd+I3RycUk/CBD11ptCyGYxvm4wNJRlB+XxIVRraJA7yQeJrwaJu
3IMzgNT5KdAui5hZqpzDpJ7uTTj0VQjWN1RHGiT5ybncrRHu55lKM14U6i00UHIILOpXFM2UXPIh
AHSjyNJegusQ5WOh5tTii63lH0YeRHXyP450pq7Tjt80n36cPES1fagUiDTIiN65WeWv1VfZ96q8
joPiiQp4NDUhcFA2GZcYsJY0Z/vf2bD4xrG9+ROqz9izy4Wv8lYbm2Re0SmdAG28EjFzEWrF0FTM
E22sgE0srKBToAKy0R1Qrln/bacxoxbNqARBuD+P1iqiaOurqqsyDGyXHcnD5hO1fdxyvfWspN3z
GVKhevBczGdms1TsFD61ovK2Ag1BAcyqbRViXFsAogIx1+ZSPrYlDgpAwEf3fsqjOD6KHOn20DRk
vC/OY3XImWZFk6zK/LAeZjW8wZFfUnRTea+jsJ2S98/cWl9rVlEyAIV8yxCUtP9+P5yOYv9/zEhO
u8i76ZWBI8kYTwrVnFQzRw51zx3H3gh9rfTvL+fO8mcfBBKclC9PJvscpBUkNXSQnSJDI1BpdOdi
KVgXsZcdRrRZf2MDzip0eWDtc3kDJSLSn2ep1IWxcZbMou1WkY/37w7Sn1yzqcBLiEWKOvdCdNmy
LQA3KVGYH5lFAfEWZNCSAFllYumOCzkX/0q/le7EdLT6I6DoRfxmkwKo6CtbwDSxQTcCLeW79IQp
7KhuB4mvbR2AWLuwKvqvMKqAurGrfyfjRfw1Mx1DvFHRYbOFkzywVhuLH+BGCnSTWj+YHhYzHxo4
5t3KxgqPbO75S9/iUFee2pmXsQZQVkAuW4xRxEiXPg3MnZfZIFplrdeVpmbEzfKrAIOIQ6QabjCK
kXDWQuxrMl5Ms+cHdS4bv/C2877SU3Pbq3xY51JaVnkb/vDvkBCxtOpEKcFwmAtlb9MDqOvu573F
1HjBfuu7mXF2dei7Tm5/dgQEQHf7cqOSx+87xXouKNLMeDIc+mwLBW6DUb1ERcG+FHD10kJ8CS63
CYBKjYlwUo4J+aNnSdOd7hwUN7EunbiLozhpP2rosTEUQ8HRCvNiU83fQQSbj7OPb+1FNVBYnA3b
0d/kJ9rF1Wb/Ub6LnmJtel0ad6v8aYR4XkUEqL0tR6YNUW5xAvyxbsfPABE6BisruRnEKZa3Kh4l
XXQj4X/vXwLZFC6dLviGqH20kwBAPicnZ6C2f3lwQn7A5KcXHOxUWqwY0ShsrD8Oh7kRh12fMamJ
/5YuQ3RgdGgIkbsZG8aBBHk8DPil54yXa0r/JiefGIZYWv/XBCBXQ1oBaSSLgJlaoo5jhdtp9A0M
i61RBvkig7c8mEonIKkgLEZHQSIiOFlLPcjvrYBKzGKVyGok3T5zv1+2u84Jh/k4DwqqRXf9WPsR
A8dE5AIC4PzzU3lqpl2kmtq21QMeF7SAFdLFHQZZOUpd4GQH9inqeXlKKwsefXHwfrbx04dr2fLm
1KEfh8Malvp9LrZlGQVgOON69IPeo2nzvWq0bB1lszIGHjwAvq8DSwUwQ2FWk2pCkKM0K/lJ6fZQ
8REIE5F91azjekCazYYs3DQmRpVCLd4Ni85WxvRc3LHJQjVgMcrJ1xlTO6lu4mZ4PACnFukzqIG/
/6qioX0ecSYx2v7Tuz1RJCKjuYoD2zTs42VHT5c9Oz/BkbgY3+ILAqqf5Q2FxoAA9mAmQxExyQ0q
nMKgiECKr9kguN1M01pLVRafN7QY1pWQ938aPvzIwTHIIf5EyZs5OCcYFew3BA0h/q68hXf8YRws
RUsktNlY+fruPDMUOVbea2KxSXVowM6rk2vNMKDGH/UfXe2sFoSoZnS/s7ZiJKEb64RpsT5jnEaB
E/zU/3pTL8NuOk4iiIbSd8JtdzefJfZX2N7OfNXED9SrGT0V3NNOrsM9aCwQRU+UW8Lm6keKnBvx
dJWzlyoHF/408LEuJNtIIvXKnQ7LHBvSjkkzpnikfhvMsjYp3pmyFRwSazvdIhbGpn/VsWhQmJm0
ydJYy2uMGAjUX8T5iDGcFWtsg3aVniyom5ach27qj4LIouz1JYWjN44580N+k/V2zx18ImqLi29W
E5T4MXzuHwwRms8A6/28IZsXshWRra+a4pNYQywpmYGv5zc00sOo03F3V0PfLTFMCjeA9ikCIFCc
9Z0gDeuL1PZfGbsbn3+60YI6ebbdrZ+kOn4sK28yTgbpsQfzdrzoO9ijzpgWjgEbgh5W+9rWXsTR
OZV6J/iX6UAq3UA2wbq4HPdBGNSfTMntBvIxLv8AVRA7ZUtQb46WpqE7kFicuru96V2mlWzfNVI6
e8Lg957UhP4I0FWBRSsCpKXjN4gYMhaZI6KYDOl83FV6TirVA2lLaslkTvq5kBqYDa+tNxnxYtLd
E9hmAfv++fRW4hPPEs23V8yuDjHLWi1TCclX2YrS48R+6r9XIlziAJn4QYSFdAuIFnAzZ6HKt1Rx
UWJLBLnEyNccAA1AXhfpBKOMW6nEeCALWGMhuTqcqSlUA+Y7m8JUgZQnc5El2lWR7UJWnpKBwPwb
Y2liyUzVfS5rGyiAZzxZTvYPFv6LU4hXhQOpYK/BUhFX2Hv8v1/URoB4SYsX2+mmRWiW11WCyh8V
/EXxg9iqaUWMdiZUueJgtHiP5oK+fOozd9/BHu8FOZoziTLFff05n8s5ocTZoXBYGa79vz4fPlQK
9ktMLu/DHhN5FhT5kXHBKQVLn6a+rxZZJ6BLkoGC7zQTiLWt/TAh0CcUOtT6hgUx9WbMpnlgro42
XTmPPHZKIt3ifzrvQs7vQUwp2riMUYVJU3XqjCX72t8hF/Fo7v+Pq1r7dG2mKkyJwszIrcldI7Ey
3Tfl236YnMP5QMhjnJbsFFuzB52svTznpDlUlwwtfUB35v+IHaU8ge2zn30ZhRa3INNX1T9gQlEJ
Q5N2K5Uckli7aKfmCM/Y1vX/N0+vZWfnYjS7gd3L0nDBvpFMZ18F3fQxUj+8hht4pUuVDxhmGuFq
NEV8dyqPrK2rALNx2dcYdPJN+wyOcQSLsHFFY1pVVqPIqL6eqF9NFY17+UwHdVRyWAgrNRkb1SzT
V9uugZXN2LFMTJCT6dS6u3A4jQnTaSdJEoHZqJv60vL3sWah267vq24F6nhnTQ3HD2CpFCi5Cx8Q
Fon2O6nyx+yHNxHec6Vm9v9hmH+KwF5F/L1PT6fk8q0AEU3Y5qoJHLrMKG64/E8zSg/u0IZ08WYk
mHhsVZS4yA4OdLOR+UiRmriqqkEN3Z0HthoAp9VoT/rWzNgeU/96PHxcThP6UOa8LR3EItOD9psU
gEAnnFVlAPgswF3ihtkZ36pgwWNab46/h79I/gX7u0e5Z+T4cNRWKwzbp2jTqgeWCtC41PfRrsuH
JMj0pDcvBfwUesVSULnnpl4sQcCsISDIzsIUqI3DRM7q5MwqckW718C3Zkz+k7JxmO9PVS36pZAm
5oxE2nuBuz97CJBcxOSxi6YpLj/waHE4cRARp3tzfritE4nHM7U69FmQGQmocO7yltP2THc6UDTw
Di+qye6eYhE+nyED4BIf2rDSPWYPQrtGCcNmOsJN2Ttsl+ilM/K2sYd4ZMuZZjVAndl7LSVIkkXr
D7dvRZ/Gqwx/qpqcVNcvquExkDWrlHigXHLTaD/tg+8clZdvKP/cTNyUdAzpkvbEL0qN98+DxbD1
ySUFPD2ayKtrN4B436doBCPadBuM/jGPDcTeA9w83BgfPtNp5YTCMtOSFOYVsGSAoVlrXyuljnmw
l0pPPPO39WDwslyxUqQRuTwlO91m+NPWWTHNnyEHDsuV9HER39j5a/B98T42EIBtU7kJBkWmj22b
TfMSu0/EGssXWvpE9Vb8FcZiudchnrIgXV1V9vUEakQ50OgFMuIY9buJp7ZDUpSrgtRywqG+aaI9
sVrpTR9JOjfpv9bpH2ArTMvy7gjv0VUIw2k9rliE/UrUTAJGn4KqGIwQ6wiGQjUYe/8KDMCDlo8f
8gcwie3rhYQ67szLeN84vpTa+a2cRdlkYPHap0k8URZZ4jgl4rBlpXkEqxjm6ypaOa7TCE1ChzNl
tE2s+2KtpfUVgvIuFER7xN7Q76CfU8wKYMPsZSd7Ew/WhQv8OfndsntFMDOhNkk5sECEsKtlBa4N
j9YbjI3JPp0bIHDxrQVzZ7nxb+lseqKQsSfLoW0ETMP8pzczeLq8cSMf9atyWGvsbsC8nNR8s5ph
qzAIMaR780wUEI03RTQvxX7bJ8UDCGJ7iNV9RtwHhIoQ9qhMJU7ORYX0Fz3jn6u+cDlOrP7VsG7P
d01T7vuGSDM0AEaf/oUv10MuJDLuo2uqKdL5HQvIjOggz56hRQEliJC19xN4GjLU3qUCFyfcIWcq
53YHBBLbPRVi7wnykToTjPnVXqBw6OPKIsAfvSJOD+bXFtJgzfRNZYESgv/NzwAz3Iy3+9y2gTAi
ZG6RRhILfnS7yn7pBh5y3WaCGR4FFzriCN5mQZTuIuTSfnzRF2Wy3QiXguKzGRUW8Y23tsVbmwhv
pVT1HUZWxSd3BJVE9+0V10oZJvp9EyP4bNmVcUeOM/LlKV8eoz/kVPmfblG6pOMjsW88LKraB0ny
HdNNvhSq1tUn3BDIn4onXzn3sSO1dJdu8gHozvJauFA0LDAujolyHEpPuqO/TCkYa7IDAoykhoOJ
xlQkK9L5oqGPhlkC1Q/Ez8/UYtmocmdzOw9WSCqaNp5lJRumqcH34SewAjruiTdy2OS3r9fiN5mZ
NjVjQDEdApN/bHXRDZendruXYBfCdQPqlqkBFDsuJAlZSUyoLwemlDpw84H9ad7NyDHOJ/UwLB8X
U5RjqlHEDt6gL+hjTptOvc2k+1p/HztcpoaB3n112nA425+uTtgPcYeIpqZ35HvAN7CpiJFfpZok
hfRh8kP9MaqH47cSoCgnguGM3v4FGE+M6OBqOroClISLv2U9MgxFfq7yr+4dzGF2ANRX4aCUHu3c
Czh8r2kWVh+EOQDnrEg/5RWPaVjNLLN8aIjhQlrjdYa4vwmAdzPEWmdD5XRZjsa162AW0ocDfmgK
knhF6mcf+hSiIJIErnKtUWV21gYGbAbAnjqJNe2qb7FMj3PE9w4cJszJ32fDxwOPNDl/hl3iIJEp
OV5WkfzyGek4lBnLImk/HJ6q+OLQnulsPwwKm2e4lh1TENx4T30YZkmdTS7YYziktljAcWSpiBZ1
8kgwK8F1GAq+Qb/+Khvk6ORE588ze3FAATmkhrN1KSsLguJYYBt85A/i0A9RcWePN1ZvCrFemrG6
VznbH13R/ULXIQNbPqZ30V44nwZIsrDmL65Lf90iZw00
`protect end_protected
