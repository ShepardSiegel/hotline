`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dRuLvOpmlN2dQrSRZlqC5mOfVM12wVJTUhTjcenGXQUUpFy7pMT9SP0hEA/epXe4ZlkXb8zptfAu
HCChKoiERA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pe3AogxOT3xahWN6bXDHO7odE1ao0Q3ybAQ1OPHtv6f2AQCzlSr78LEUyH/Fu3XJeEWhU67y5Etz
V4GlImdpKtgK5fjV3sXtWQp27LyJARt9kJjdEUNf4zljpT6eYrn79/nV4q2goKb6hCJyRPmpqJPP
/wqnhFn2m0bPFfDYvKU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
zrikgGjCHFnPTJzhNAla6o0liuGdaM9PCMyNqoqubm77SRuHJX5oEqy50o8LaWoNmn9vcspbaJlk
kaKHTXgceASSioU7VMgFjSzVln35gtkRAJxSyCHcj8q0Oi63R5wdF4irzZwdgVxmbOP/S8qKcj1M
+wK40oI9yoS2PperB6uOUcNedZFeJl0dJK5Q1YkDQOBLt5wivgGsEwvtN1YBvpxLzK2U0Q8JXzwR
wrtf8HB55L2IrfYXgIt72GNZRefRpnqOyByuY/Dn82ceO2OWQ+HRJ6AfzuV6HhlbspS6nrIOUTvM
twOtSiqx8KLuzuzXCWnV8gzN3dWv5SfEpN0+JA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
USOWoBKGc5N7vY4U/TTebPlTsclEXWHxFARpCsXROJeOjVjnYE4fxmCTg3JpFyqqq/l0P+nqyH9d
Z7qkZoS6o6yJZlJoa9URolkeXWi2lmrv9+daqeQR3Ogr2PA42AGmO9eIGZRB2zMV1tychTLPnnEx
haJhcPb1xLbD4IoTssU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KwxfPHyVRDxW/5k5/AW85FbNmGQh2G07FFnXPTNHZu1WambBWiNmKDoUo52vdBcKnt1aTa+aKrWm
JUzIbPOJ1Nvxqw59pPhy4y5IcIRs64uR6626fTBf1ZCx7gnwK4axOMPkhg2UM5lwnHJU8yb1sZm8
4JuICg8b+i1MiBRYOK0uJeyBeeTnok9CoAdWJJgKFWH91CeuPO4n3Eufa3/e4QZfRBz4WEMhSniM
7Jm2rMFuwKk7oZ4uIsnvuSWrWBaPLhP8KSOEp3coWKd9k0CZthpxmITfX1mDCvf4eRS2PcJ6iwgL
FUyCw+uAF+7xdjAPw27k117x7faiCDGoZnHxsg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4928)
`protect data_block
LSzhzeyreRCKOkisOYge93wt4UdktHPFo4ERGrqyeLMs0qRoR2nSyZdZ4+71EJPvkBj4t4+aHEKr
FZ/xekzaPZkchNGDMTcPnBFbuH4Ux6sEeLQ29Qd2O7wEvkWuHVqB4Ldod1MYccEBowm+Yqm7aXdb
Ciw//OH/4B67mZn4PE+1u/TNHpYVfUUb5COUPMtGBjh7iJnF3Mn1izsQHjeGObwrFTQHC/E56L39
4PruQvhh43amYCbSpM6tGj9rCwIU8d3WO9vRNR1DALab75pELFbpPMiAevjiAgDfRG9hLXHCPsyV
/E7XX6EMAL5KNEzOW19N0v1KYXnoQuqHA0Mf965Fp1kpC5CYb6JctC+28+djD+lP88cz5dF83Bwb
/wt6qQI5vDFEUar/W6QxE1E04tQkx9656WQ2s1XO//ZnkRJW6EgtTOD0o6BaNiVmqTaNKxFOC1Y4
Ws0/uIvrzrsvFeu3Ct823I4nsOQGBApARcb4qOPDdjklep66+cpfbNg++k9eu6KkOXKSa1wkqPo9
YWOYQPAn4vrh9cBAPJcIEbm+fIHlprTkjiyYbgN5cS98cxtHsGz++Ew02H2knWFs0tBEW7m+ioVk
Iv4Hp43I4b7q5ygqHUwawuzsBxNk8IiP38n9KNSmdt+isc2xfQASvQKVsGTGxebOlhTwn9P1Od3k
1q8BM5jNV0DYVEIuqlFk7OVqbYSGid5kbQ1dEGL5esrXUX3mCfQQIQKm9XrUWewUgv1CzoPE1QWX
4mIUJdWAGNp10bR6Ia7IxteRzevxfRzpdXrFowIfYIJ7Z9Cm8h9Dam/wbluoBHpt07dpcJYCzr3l
iTW92m51VIGAb8wKFfXc4/+hTu0UdidDpD4n004xH7adVRYIh8y41zfP48kUV20VFTk7MyRL1xPL
JK3Xv95eXK1pWSbXKdGxTR0WocOjR0VWQnXHT5ZPjYrCQ4t3Xj6Ej9XRO1aqbAxv//w9QF/lcsgM
Tc2Hm87wrpPCOmRV148x2iu71f+qEsxCG7pynGgOrRPRbFCoXv90pwFTtxG8w+t4bPnRZSh2Y6fH
W1pnL+KrD2fTw1xENwAHu+4e53Y2OoSlk3tUhD5+hLRKJbdjOL32RLrRRG+NkaQ/i2bGRzl0pKJ3
G/vCyNeS5/zJy/KiiUqdXeEBd9MMGKFc+pUB9ypzMrlt00lX/X9d+TqTYgeI16ATKimHC8TZJD4B
HLYUREkDsGgvJQRQ5pswT2G4zXrmfVJwRnb/duIA9FOrLMV7SLQzaBir8UPh0Yb29PJiOJeoF03b
Sd2kAO5tY92VUEl3R4KcuZgjK1aZA1rLRmKXDDSk6kdFOiNRqOAqIhIu9piEt6cwPAK9X8A1/RPn
xyZ2TgOwV7lq5WFwIaU9yTX8rsiDrbhjk1yexgJLf/OvJTfbQmI59eGHBfjrWJMTI/iU8MG+BMjf
VW2mMrpTLZ9JP4/r+Jr98YMZPcNdqhaq4RuWlfCiuIlz+xVDww0SlvbmzWy2j25kIlswo+hH6Nnb
8m8UoPHGComQeyHW1zYty3lxm/ITUD5gGU1vawr5RogHJkxXXGrlI6sf/byfqnExSaf8bR9xChMg
8L76W0H9FdS6GBEX5xXZjG6Tjos4csFVtrodWWugNqov/bCsM3VWMjAlwK7ApD8Bx3mix6n8G9lr
J1Uz+2+anjGGX7UX3vXDWhUMuW7yBEIFnVsSgPZbjc3q+91LOtjhVZqjCj3q+OqIV25A8CooAeWy
BKJJboDLDy2eV/Bhb69XWN3m/ag4ec2Sec7XlWd8qz/xjiSbepp0h0RG8V5cv3DHTZ3/tbQi03i7
84qwE7rdXcRoi+KKyCNRUbBsSA0DP3l/3JMi2bOP6Y61F7xJkWO7GV2zmsvhUT+gDr9phwSKo8xQ
7gz3F231Fd+qBgXFfgcl4lT1MKJXv0f41vw5QE4ujXwykwjoenuZBjb4eKC6esgmH5YpGYIfjJMs
0qVIUsy1wGauoGo0R4y5VSUfB590WX5leXZW2S6H7iLLBRsMRsc+sTA9GxXs3nggtRMC6APzYTzo
4efj5gMuCoTr17qpsdHi1MiEujhJWLX9H8GemJ1wyJboG9ajvI0t4++XVOPwzyODsh9QvklZJW0E
o2oPNrVBbPWPNfLfqb7X9YejfEo45gtg1VAVrvOfAcbmX4SFMOQyp1fZtWDrdIJCfu87lqEN+xZA
ey6lKRqKZa+X8scpnIrTy0KNPIFu8YV1iF45w0U15CX6M3nUkq9Gaey6kOw2jIpITd9fX91hvX2S
fp13LBLzRWuu3OVgAlYY5UsSROzlwwGstfjbvspVmNi3Sg6Oa0Qqfh1iJFm1/VkPhugsTiiDHvwh
5O8LZr6DpstKzRNjvGc1JEokJSs3MMAx25fHlvMtO5/Bab/QhSp5cxUzpsIZ2sXzFUISlVK3UvUg
wnZTNsGg2cJjDYYj1jVcHwrIavryKlD/TAfVOf2FdwklgwmGe4KxvTCPi1vU9eELEeVZo39eiPhf
jeDANLo+dE9Uf1Wn/L6eVs6Ez4vBNTD9V+7PkBOqZidK5tVbEM1vtht5u8leYmBwtGJttygHcl6z
jCdTTo7uHFQHsTjy3dQXa2GsswWLaE3o7402nl3gt3v3hu81qOGM9Dve1PWqvXOCOXLMcZzSkCUq
jr1YAXZnAhsQbdfWdG3mw0BMCnWutHcAO1w0h6YNCFuooBNENXT5lq5m7W+QGFP783DkeQldOGjI
QC+oC1S/a/sRZnwcTEOCCu9NrYlV7tIN6OvEL2m5BhBJXWX5X30FDZUJ3LHMQbzNVGPl9dOL6t2h
P0VpPCpNJZoTw8ypUVG41w5eagQnTfIOq5ELTgIN2SP2iwq06jajsu3+bpPakNvcBCR4QDQQ6X9e
UK8/cIWenO/DbTAgTI5UNbLGh2Lrkc+bA2XxMci++DEeS6fcEE9Z/pVLFatZarigHa0toj1TZt2L
r2ujfUguVwPLk389dwqU7OcSEjtbl5SIWZCn3mjl5+Oa7PDSG2EOj1qxtt5gUlb9qSjF/brVxTxq
Oj0FrWf1fWQi89zRe0D1qXacElD6N6uY//krM+b6c/SKKzpF6n/d1iF0w3P5NiKeqNG5+qnfMinr
U5SxSTrKbNQJvwRuQA39omfVtWg0qcfowbxJGwDzHCOhM6muAaog8LPSC0EOLxt2cIln81+3DEpa
zunski9EMABQnRse6yKEkAhcDdcUTH4+kj/X0TWGL/NYsrm8nskFgAral7tX5nLsXjRoK9Hplhh8
jiDj/YEf2lkyvlytWtNSj+63R5GkwCn6PRhl2oxQHQo6hdZKqY9V65k0M16m3FmI6IXgve24eeMq
myANF8+0oW1fqzzbu6D+ZNEjINw8PWI9VxtZFtBXEuSzOq+WRUYKEbMddB12vPBVCsK9wf6aKOMe
QzWas3G+8GJvqJtkluAn3mLnkMYN7PGSW2xEyra1ZVYSClTzuaVqkiRhtJQiQuC4TThgJYlw3PX8
iHqtkn810ujtT4Xo+2j7nm/ALqbQ2NKzIVRLMr0ZtnTEbh5xWWi5kAtCTyDoX7ig+08KOwJslDrp
KCdWgxOon4DXwd+o68RLy/lvzdB4bpLtGzTquWDn2DYEwVZsvHd1/4lULJGDzjuVr/QgQIo0F7Si
UTBHKsVVvNjXvBrnUBvb+gITzlF31jSe6ukOIX5ZCz5gTJOTdRRBT+QT9vWw0NXcNnlAdFLruyxp
hziQcBX2b831RSsKsCRIbx5NirF4A484McTfotdq1E5RIirq8vrn2Ubam6megBDiHFslCsTy6zv+
tVpMiB5QUOzhsIb5ErfI4MQHmfWvEOlVTph3dpjxW6/unU55NeLaziWnRFCVAYHCpT0IkjYp5+Nu
o6SXzIIfncoCVPhW3KB/PpwQaDOsTd+4RwOeeQ3ZPtMrN3b9yklihdNnU8x4nRqNvDSsfQAS4Xci
nTHBvoKu8cG7zfqSMmNTXnl/F0F2VTRl0GMEKBq3uny7pfFtvh1FxfrUv0UsrU2ufDjG6dF4l/Ud
NPLEumirDauXtA934YoVtH0T3km4OdMcQbo8EHJfOOrU9OfulfXJV1Vi+7sECpTG4uakJYv/XD9J
KExuaGmME/KyW1x7YJDzloYMVjIz7EesKYTUbi3zDehXkYhriTjmBVaxfdSOiux739rmzjSP2Dnb
PyuWkYmu2n/FEvms0tDdKkDuQiKeVJ+UY6x6TOjQ6O9IqYXKWyU2ZL2EFwfsqFWxjYsJ2AGYnnB5
anVWPCxAAk5jcxRi9/lD2ptrOz7HrgNoU7Ca85epqEDyimcQEj3TlmNOefiWqhliSotr5D0tetfx
dZpltT29mbQPLje/Utebpqy5xD2QQUrEu1s6vVHz/2ytmZqVig+eaHzqTgCHafN++TBlmqEDqcbG
ing+JMZQht0cHORh5ZDKEyiT5VUeFjTdFTgh7kY2NF2tL5FxG1nelPQeJinYAMbPxIUVfmHfZ8ZZ
tVF5Fy9xrD7uFuVC4RglY0bErP9Zqb38UgSlQQiYdhHlRIOrB4XuMCytO+YB2+dxqXLCVTInVPV2
2XqGXvhRHd8346m4l7qDtJz+njI9Nmsbbtn2/73P3NfZR54d8HRNGxBnNPUcym9+W6CDH0Q9MN8S
pEWiQVboyrhyiUn1tCmyEaftpdoPY4jL1FIlPnjiXtVCB9PmFS0bYlK2PwmOI3Td61Em5xRMkSrS
smyyQYhW/UBjk4Z+F8poUcDfABKhoAASYBMXsxJ54Cu3pxM5oxCV4zGcMbTPwBlqOKxnZKmDZxao
sjZytVNTQy+64CqOZLjt3OFSq9xJPKsICdXJhjgrjVxBIH4RHmRHwSm8NOBurvgvlWFOb6Vph6N1
iD112Wgqo5rkkgo9sMEtPWUxF4R23yodXrxPd4t3CTTVjLQgGCkVfkiGDBoH9OkgyIsb7Tlgi7of
7Rt6W/xtZtQEwcTHSZb2ve2dkqIHiXUII6uc/i3FUKb5YCb/Rs7vv9Rb/JmQd1BImUTXuJ/r0s8/
lKehKFue3Vu5oFpPwX+oibQeiQCoa+CWXsPQTgdLcQWR0X8OketIp30U7LWl9DUSWCvheV6toaQS
8kbOvWweeEbvn+yi1YNRqoKVd7HyBvgYbTnn5syfUcjkB3NpfxSQsC0P7/UXL9zs9T5fEFz0e4Ol
jAN/cwsvDLtt/NVIIINaNwIPIU6ZYqSmomDb3J/uJn1IbAHbcO09greQ8JlvC+Lv/YgdWgr7VX+2
+wfvh6aVx7BCw1h8kO6bCyREuMcfjh0rxFWaNnfKM4nf/U2uv+KLqzf0C+d6b4231vHuXXzVQniu
Iws91rN4tIHV06+2117MQctwLnCam/SKjk6o1E35Bb0gT0B8HfmrAvqaFsUpGrx+AUbrgANjGVYS
xKnfM0NjjjnYZrjUfXHfzFjgleerRDDc8mMfzsVZLFhqPEaBdVgpIHWenUSrHScU5oSY0ZXmm1GI
K1wvJpIjrnCotpKWqy1FDIl99FHKHDwICaIJvFfJ9cKcxP0RbBHtzuEnJmONUel61Fivg6FJhrU8
tcyJbUV0+3bPRKLI5INYj5LYH6zf37nAgdBy3LzHEhUhsFL4KRznClPfDHB296melHyMRi1/Oqx9
B2gKZBz9NlyBQNnHWDTRNltbslRcSrrr9r8+jbWz07CX2EYxotkB/eMsdESi+CGgRZhbsgOK2/MM
DUvFhnOvTka+r9r7HYJcVxeGWeehc2UZWOlhbRd5bzGnhqlDyjQZoSXfcv9Nl4P+kik40IKAfdBo
YVnDwB+AM3VcmWpnWQF3LSPHW9puihEv1o/CLk7kHmVavLFhZ91VLi0iFULkEM45BiLEyyhd4v7D
EvAfhSv7OFv4l7ugMU3toJMOUuDz1yTatJ0CeMEbzx/0I6MwC4l24st085tr/nPXLtEIocqf46U6
Eg/gjIu6397CeQSUn9H83o7wpG3c9cdMKBsG0zRu5XT3y2D8wq3oAF5V4XZZ1kkJgKag+HpFHMMB
4bLGa6EBJEMm7fX3r62v6km9layLT3pWHhCRm3E4fek4FkVIbxxrDikOW6u57/17ymxO5TxeuZZX
UYwMBEArIlpYcOYjZK3iWjc3PBj2/GtCgJISK/hBMenE2ywfX+7Ps02eRU2wA599Axlrr97IZCt6
Y2/LBrc7uXovX38+TKe0dteJ1jxQVGwzMmdG5VtzCjvShMSU9ECIjYoUil18Xr/VrBadInHmnOxy
X9ILUZ7vj3JVx+N9uVR5OVqgVATiQknIwSo/2BR1sWGLBSo38zhCZl6ODtsG1vkR0wD9cj/FvTCD
cQnIG3XBczL1TWDh2UbObbvZeTyMlwFrYuQXMTpDlT2PRe8kFd2L1oynHGe4kDtLi7ahzCYqWygZ
xkL4JBa4fvUHmRZnrxaqzN51QnL5OxHb2V7bP/XLN14PYY7IQ2HZtYVfiu8Nl3atixAw32iWQa3r
MfglPbjVcUJon8P16VAZMyLtRCC25dXLKqaj5JcGIrQO5y8fSBCCeV2XsfXjAMbp+V72JCm0zyIx
HY+iVC8zLX6FdrSYrH4fI6TOi+BVOzPxNNU=
`protect end_protected
