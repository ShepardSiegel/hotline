`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RnMGIF3ERTqvR5TxUGvYx3StC189+fKVzuJ1bYZiu1p9MZ7Rh33qLi6gPqiBfiNwp3KbOSxSdXVJ
Vu7H+Npi8g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gVjpY2U7+ffzSXvV/5C6yAlxP8zlzdDDvW2ZwBcvyhEubZDiRs+OiyGMVqU3ajRoTp+BRM4/ODZs
7DkvfQkgm3eQj+NXwN/2wVJ9JkAALHeCeAcH9p4DbA0fXPLA44bqgdJWrwVRvMu5FyQNNAzZAuDF
34g00XpqfNT09euq/yg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
B7GmvIbKO1kclT9KqenLqTa/dTFxJFb+31BarIFbhk0u2JrEGkbUd7fH7Z9E57TxaaDBIZ8SPJ1j
1/ui5vg4D0pMjJbAIsn/4cWF4PZRQM4RkiNtHjq/XU0EjXgD1WJzGCzq1SOrV6yaEsBDR8vO6O0X
JQ4PWAifa7PQS2+hWJt1i00qVd9EM61cuu6MKoeg3UaZKazgOArJMozunkp7FQYFNz+TKY7xUu3J
fR4a/9Lbp0zCB0jvDbbBDufn3Ba5gmqNB+PZsNfYTrU33soV0BDe2Qp5CdmNWHEa0gHYS9nsJ2Im
V/KV14edjh+67dlFnBm6TCke3DCteVp//KLSRw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zcwDqRdLTH50uuPlo/Nk89wWJpG/AlixIkZKhznnyQVZVTAU2LmEde8WBRlqc6kIeXQ4eBusQ6rj
mXbNsmV/PEj3fqbbKDfa+6pPHflDmHm8VW+drKmZTCpgxfdYK9oAXg0E8HhUt0RE9ocBveBmXHV7
UAnmQdiq0IOO+TxGBRc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NAMW9kzQBuWj5sUIT/OPKdQr0EuPiLnrcPLSdWXm1UM2pdIdebhZsKrGg0XIv1SpYw6SVMf5eU2W
0HWSYrdNH9yPQYdS1qGDtKVLx8cL/EvOSTWxydUlYB6nNQEIHO0FUWai0EkslQK60mVRKXRAOPcJ
3WMndgoryv+Wei9wRApgFpIi+JU56hB0ira9HwIZpSPi7XaR0IaDLTJRuXhivjgukQuvUqFlHRa5
uBMR6XP5fojWdB1ys4jVP9Gd1DQufn0E6y6NztimMfnfXHCLTzYIaVEBxfN7szrIbgRnkzAbH6Gf
BskNVZIMTp7CEs476dFosRn5Yuz13WO3GH4TzA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10384)
`protect data_block
GGz+OFv2ZmlIqe3e/Rz+bgrj+5Tk1XLivltxOJAhIzCVnjjCQ/Hal4Zp6URX06ENYg2SSdH9gOUI
cIKVi3+rL5uW9xpHJGvwNzXXAzJ3kVUVquGOy7/nqEPm1LvPa0sx9x3O2PIEh0TRBgqOgwMiNxMU
C5bqAYB+2g3jYLB4Tq3iSLieRv13HvrVlNcLzS1KFpWVTT48LwwOXPub7XtyA5ThvdOCnmZSYkJD
dCv1SUK1KlTh7X5BtTQCKFvTw6vNDsGjWzMx/H83ScKg7D4wXKPaTh619i5dbwLcFS6sEM/Aa55H
7dLOIPOCvCptdVcbLwfY6sDGfpN6V6iZzmFrAZyh3iNhWS2J6wsGFIpqQ43MPG5Q7FXL9Q6II9+T
SZhr8n6ME4h5Pl2V57npKpp5n1B36ZWwt1duYUDeSd+1Qmmj9ttRwh2CjSsGtWxtelnsg3mhCW+e
rB9+Logy+ZQaY/RrYVnki3tgu5m1+XtfIbXGXX+nrbVqB3oH4HblSqW003ervgWNKn7/PVeMUdeu
UXhiYOShk4t9QfL1cwbi72iOP35lcYSkud9QRFE2fA4FwR6fnQGtnEUARovHpXUH9Zso9soqRBlr
DAltJohwoUIDnO2AnElcwxQYbMvDy1Sz99P7gfQnaEd4s12mcDyrl4/Y79KIBy9ui0X7gRJZ39ji
VkB8HWHVFqYiVw/00L6NJ9/5emwqafcb1FHi8PcqJ6ZQURWfKly5pBdFfhdLZ5pr8RlFYqCKOjhp
ptcZuDJfb5XsGAEHkEWr5Mvs+REkhrzBeHDQOaqV+Mf6DW++oorwLfTYQAIOV06FRjBKnvBLjG8z
jROlwPJTcbWE2PRoX3soMfBeaalGiydkSqNwkkOHo4ERU5TC6+Fgdy5NDmgIm6LzKtPxm+kSkHU5
/CGwCvSjjuCGFwAv2cH7efb8Y5jOEAPyNd0gIXapHdBlkMSEBJPqj/qG7wUTu6HBFEVve2/WQhe4
o6szYIOwRUDYGu5A33cxDi96e1YVCLrATKxlZ26tvt2w76HoCWTHIOKi27RfFjJco/gV1q/xJgFE
ql8I+8rmUKNMAXnl75/t5/y9gk2pidh0StGAmHmIvisTtsZ82Zna2I0CD+YyV7soj6NeXilx+peI
jZ4uyzp7oty+n56Qtp+H8GEwiTb/5xHgv/reGxzHDk5exuh+HX80ZYc2T1A1mQPiLNkQk48LvtUN
durwXjZcEmulkz6Rg6WyWAWXOLunGu++auxPyNAWvtaFfSDXEd8G9dGgcDJDtm2me6DnUpikE1P0
Lpa7KF7ZX1IjfzRoDS5TRpRyIkVBqYcI6rYV5vsck1SiWna6JilNCHO1I75ErDKxQNIrBlmopd6+
l4VmbXY8FL8B6a0HnJ25YyzL8ctMkLob2XgBkHwbkk/Oz751anH/ob0SkuR0TtXkrv5fAr9198qL
wXVnnknv/tezkMcH/0OtqmhppGRWfaHdeefI/H5cPO6qt/fg6Lca+/0fd7LY8CK0PkPI2ROU2VeY
N6QAIeCAldmhNmXUUXADJTGQ5ApLktPCASjfA4J8fKfypVN2zBzNoJtcrPpUzx71iy7fsCiMvVMK
r9Zu4O4Pti7w3b0DZUisjjNO5m7BvVCy6kMIp05w4P+XIpkMYn6iOsId63fn8lnh+73S0aj5G+Yh
96Y5R3V2Ot5KHAM3nnp9F2dpg02IQQ256cMzBX55LXDBC4eALb8ihaEu5PLBtSi7SFSpkYP9/Pqh
9PJ0eDwdzAHuQpY3oTnKCAIw8D2hgg8tLadcNo+G/oGWWk8gGYSZar82YBSmnp9CBUhUR4QyYW8s
1qIDUishvR/Qf5oFByrUJO3R1L7tbY8N8Bi1VjdgAHc2CvCAvT9zcdsAL4Rj1UtrqmAQDEKD1SWL
TFxRcV8ACU5GUT+yFW/RPD+0JpTETOyiVSMqeyCd4v5jKE/FJEV17iweBLdTJrWGPlJhTtyFH2Ol
ayIg7MtVDfNAslCEfrsEpcGKmToTt7R/UwcOq92v4AUT9pPpcQn7cayJdqHYfWYi7ttKB5xGzp/4
mhpn1BgkDf4HMIHAEaF6maYVj+KgyLskzTZlb09hlHNY6/4cUY+7xgOeHWt80jlaOCQh4b5drKOO
PKLDV8QNKGtt2wGrSMih5E+3PkMBx+Vv/8VAE2eE3WpJ9inc9zaBzDQJUTb92d1qzv9DsmQ0U0xQ
2djTqp5vhbYBnafeAd6RsEeRpqh7liuuRuasHO0y6nOxq5cY0qszsQx+ERL9pXhOmhY/40NDQz6M
4hxTEnPu1egj2Wj0eXfhjjiOieF/Nc7GrxK0RMlFlu0B9UFtZd1QXwCZH6OKhU1z6mZLIQhrS7br
0ONkYhWl1WUvfbkKWmlMsUJHMhE/jiCJPT84qvq/IQAbbPZs6BSJa53I8ZOUlZOyMHz2NBjCPbIS
oIQ2Qgkqg9fSTveXnltshwYPCoje0X0r3dDS4d7aWOK5SS46qirzBPcS+94G3hZ85Ygb93cC5W8b
t005SG8QVsFemIOixlG7F0ftHxomkj9HnlCKZKhMRUOE17MmPJvzpjtS2IRj0VvW9ITkpH4flu/H
dtxg2IL8YHmwpEGZe66vlQsyRsSdr6bhEi0Y8K4QThQNKnpAlUWTzuJG+dxRJVTK9hPHX9RxgiEq
HeYjPadPPHH2JhX1BaX3hAyZX8znBJNPMYKJR2WR97/CeXsnF9WfuSmJipdxcRpmPjblRuLJzxxV
s9FYAkiucwAlsILxx4BVjm1aWMi8RMoi1flWDo98AzkdfXGSxSyxc/kLJFFcaLXgbBILMYPHl1tF
HGWeTei9YBCkNxEv3DOetKydy0v40liovtF9XhrRaTuCs7Bw/qM3QUVhIPB0/WaRL/3heL39yfUf
CzOwxuuP+p1o1/LpiejNLjYoMsgtBjrWKmUFVKhCDLiw+U7ftbL7JHuBm6VJYvg94+Y7IGE0KmPo
UZbv6iPD9WN3YydRJSNiQS42vVh0wp0BWYLBLa/TbIKifYa6zaJ3a8Jo5HTF6VjcV0sf/WvsnJFo
DWMMlZ2oo0794YEFaRitaSzy19kyPAnsDOo7b7S4BBJox0NGGunhC0xYUG0BL6OfOUI9WLwOxs0L
2/RUiOscjTtVdINwrpL173X9my2ZyHd6LUs2DnVR/7LrDB35yBYl/5OxDbRN2wLzXukghjNUJXYo
o373+K4RdOnaAPgT5M6vnsm8z+4ClwXT08+jipzQKAcTzHKHFmKkWOvvDkO6lvv9SBtsSsnfrGUI
JeORRDqELfs95/Mg03Ub3jxtZRnGIRZ9mNXFUZTtDidN8JmbI3gBa2aK3oxxgKGjrf0GEwhaPCIa
lgx4meE/zzMRe5RIqXYtucj2hoMOuKwbcGjKbkxaTnCiEukJLsubFGY1/Ec8L17WRDGb+6xDv8Bg
rXxB4eEU6bMCCQGE4mWZjyh4ihYaZPG/AJGfTGKnFckhcPCRQSGxHbUW9M5j0ejsA6mva43wA72N
x+T4EFkxDPr+498Piugez8+MoncZcdG+9hblP8rBF7/XRyainoMLbksM6x/8oTgJnIyy6+hQ/YbX
QJB5VLtkYNesFog5hRYXkuZ309cw4OaL/nuEadtyPw4W5v3ZQ9z2rlsBppxkGPnaLE+Nu0+z85kY
6qbpdRUkwjbBuKIh1EfshvwxSAUpQ5+Vnmc/s6dV8vihCbTahVVF2YpZt2KbnfksOZNNKKtv2S6R
66Fdco3h1GXg91eIsau5STYEhG4S8JfrEO8faE+/oTWBhoqwkG2qfGQVmlWzvJP/WeSvcvLN+WM7
/EgyL/H7tsu7hxR3aNojiE6fSpSCbUn9IF5wC05ChS+iwAbcdz0ujxMj1lcqTdG7cwfzBE7ybkG8
ydZqCfW7lHOtTybNvbMnqRQHTOAZhTS0nZ/8lYbvvITo9ab6SZzyfJklnNwnj1kbTVMsUEqXVT/c
HW7aAhHZ5DMlvq8Znm2C8fecFX4x0LQk+cFfWagnO7wmPnapuaBqA5q0WywwgrKIXpHPwx+RRk2I
IyC6AneOiwOnRTq+lExs3dC7FQZ3JTTfX3GqhV5UC04tppIXA+fzVtdkEcX7hXIiOpSlLgrCAwFt
deT+s5eubqF5G9vEKiAgHRUpuXazoRz5+r9WYIDqjorSIlozZUr64YO+YMxSyexsNljwQNuAMoMi
bo1G2WrUZnLtskXET28e3COKIiTMD0kIozDj5z0yucKX2Fqc+/phJtYXbdhydLVan/xuD4u7UOW8
0KnKO0Em+fZjYGQ9tAQ2knR1A18rr5PtToBDfqCZgZBMTKYKIVh9rpo9oLqt4XA2oGQ9eqjTLi+U
uCw7NVRHvreNXGOl1IBwDuOZCHy5XIU+04vsrEQfiJJPVpfHCSVD/bA8ak6+YRMTEpVPG0YvCPDB
Dz3VWnBeqDUPV8Z6JcYG4VrTLYCyvPB7bAgqgYW0AslNyWEfQzllQnbrxt9lQkf/yrukcMCjAEoT
4Cpax0GUYjnz8ZVOa6swU7p/hP2lxb7nB12WF7zqcRjf0FReIXeJx/04vJA4LNTovrr0xeLLjJml
OIMllWyOp7B7vDICM4DGE+GGC9sf4lTVKc8GlgM8kIZFLX0GTE+2bTBRoDrhhL8L3/gQ565WKJWh
di2tkl9GQj9gU8dalEHc9rQ8WWXKp9RpoOzidIAGpPJ++tudongxhqF3JCn6USC8mU9y0xEJzlLK
qes/0caIacsutd5fn0GHY6elI5dqKzFmt+Z/tzcjJopU/yi+RBdWEmwZjqXb/VHaVcAd16lE/rHP
zKfQmQU6resBovQP8mkPsk7FFpuOjQbe6ztpcXKhBCjf8IqEELEidBmKKAW5a27etDPe5MMUkfnu
kAqgDQtiMDstYhAwYiB0+MEm7dqwrIKtZVbf5J7o4b+oDTQSpLMe6sRvS5zPV0hMATyM8CZhj6sz
eHYoxCL8AszgHkOEsVN3TO6hrRwA5pSP605/6F6M+PXGeldnaRJIdWb7ZG7/hfhH8+SzF8Y12t4q
2F48cUDpjVGYYOTOhEH1Wl3pt3yVt5v3IhtAqtS4F+OxLE6a0AwxPZoB2yRUIlN7vtZFZhFF3FZx
WJUeQn8mspSK9ZpOh2kAbkhoyeMLmSu8d6IuGNJ8jGjWRO/LiAM6S3dkRSy/kO9CnaMOs8DMeMaV
ySO8MTPZMyE6NB9z0CRUYO8B/Ksa+U6n2u5L/Kykf8iUnnhrNtdu01E9przRdUa4/vB+hqx2KJyQ
IfZIMQ9hF/1qyC/Ci7Cw1AmMlP8bkJ1RVXt7521pRaSXcCgOi1eLO8mZKL0gcajgCaG690+QBIf4
6OvKVHNuZHI75IvyczjEyxsFFBH9Z/9I8tegbUxnsVAgY8I7dNHc5PdPQif0Vx5s7EEJPUYgKiq7
WBuM05xVFWWnfh1/vACOwKPQ2cT/fn3bpyDhROXSAY+a5ej31NW7DeHL9TIQVlX1Pbvt73GPJ+RJ
3cwRuwEW9p+24gnTTF2KxZHEjrcBRvgTkKFzh8H0kqTGCgRRD+fOSFkVX/fFXUGVgGKvRYPooHxw
f6z9/YwxtwCrn9WQv20nsge1rr1WwNhaKA4STrLZ00l9loao0BuGDUXnC7dwAu4pBj+aa8VlYqLW
5juMSCmpKx39k91MOqUlah0kZFuzj4w3TuE/bJosC54JSGwdxhWstcHYrfsG7qJudkv3cErGBQRP
U7OtBX7YOJg7DVUPkiTJJiysxLdcwGC76bV1nAnSsdmv2Ax2UGczwan/EE92qQOdOOlb1ws/ogdM
SMUArWhnIzXpxHln1Fo4zY6XzNsb5aEtgdmxLTiaXnobpZ0Drp8NqDPVg4rcqFbV+FEssGXt6i3I
65hXqGrmEBH1cvMW/Sntyr6kESH7JYEZAaG0IMEc0E6Upp2EZclqm/1gjnNnpFPq9mhU5P5/YIi/
FSKvE+8iDKrg6ORvYHYwcWRlZj8LONa3C374nfg9WImjP4IPVgDTxbf/TlHH/gXEy8FW5pSLt1Hh
roD6I1yh9gNwghGJvq1Pkw8rTi7lB5PK7pRhjS5ZN8/gMVcs3cIzrfT/1tFdyxqWbFvbTGgytgOJ
BmpknNj9OQG+gjF+0+t55ZRAk03LPTXvRdiKuhFAy43nuUXfJHQ7GpTEt/CSKwJ1dzuOqrBqI1Gm
5y1NN8pLgrzTqGZ4s35o/1T/UoV2mxBQbqai3x4WaVd6UhoTpVcdQXCumuGSk35yGvufg1pOPfEo
bR6zpJzQujr4ULfRx03Dh6RbIGI2UPqOr5YGK4n4bv2u+/XK/U5QueFcbDU+FoXk6tKKg9q32IWB
6XrhXCJL0T1SkxCUUkkeYarCG3ZrxKqJ2VE+lHlcxTvKvuE7Zaxg75j7LL/xMfOWRg6v/oe2E8SZ
obromZY1zFYYJbJW1sRHW2JLPxijSIBe7AUk5FsPyx/5MnXfDMwQ089CExG8HMi5E5MNDO9XD4NR
9Ncix/r8/aXIV46Y9966UGOAKtpCjx17zDdLVmIqigVlJcBbRYd3e3Ka/ZxeiEs5ZB5p/enKb9aD
Yan8Zv0fJGTJSOf0PGRg0JI1V5+hTngH8JarBfyB/ZAy3i08ImN2/A/XjYzRPdJjFkB3rqprermn
U+troysnL+N5sylQ67E2rIIRknn0n2V8MJKKDJPjwpnJOEMPsA4CXnYdivlpIa2L7BEDpMAuFFiM
xFuqSQhyTjiAM4cIsvuN/kkP18QuIZROJ3T4LHzNF2Dmr7VBYYe71xyW8h/V5m88TI88vKP+JJnK
zwhhdpOETaYtPZltlvxv/B2KyMEGGQDTOY+ixW1525lJl+I6T9txQMmw8EkC0Attn43ScfhZtS2y
R7EK1i1sJa0vKZ7MSx8hRhz+zHTRCarx+QpP8lLaiTLTH08cfIFTsK4i+RDqCZfGFE4hvJwl8iil
2p1OEG5FNHliKoC87oSj/rUOjDBadsW7iCdXFpn8NOCL+RluTX8oCc97CjMPQoCYgG0Lcx3YSQQ9
V09TK7xOmZLNIQDdm2rH4NCKfrJe3vgwY2Kf8KT9kG+f98VkU5kHgh2OAT0T+/vg8/oYkeByUL6r
2txli/KaA3ZfHV0E79Phi96DOVxRDhcJDTZB9LhH1ZpejwiIUaAl8TsHbPDXPk3IsPRC4NrtoXY0
QCRGyKxYAw9HddvLlubbfycwjTOCzuaCG3pPl4FU5LHsO2RgRUUfxnv9hr7noO1EFuMKRDLF5u6z
l5N0CM8gY2A2zy5lpL9FemJIkF3Z9Ms7KgTthkYeWA9SylIxu2Enm06/PxHirrStCPqlUV72vNj2
w2XSEthJ4iTwk7Eesz+p+pip1wBM2AQFtVVerE3hirEnfef/py0ofvcoJGLhY9Dlrf8U+OCt04If
UgESHOlrICKTXaK9OJy05nDk43LRzL0WkxaYo3hjFsAI/8lPGxmU+91Pl71hhqK29aiNzwB/Djni
vcnBGV4Rf6+/nNhZw9J00UVsQlS9dRqfFw06zH8jA46077rqXtE9RQAGqRGDHsUta0yGSuz3asWT
q1Yr6jyyYEpIQVZAW+TNoF4KcI/wbJ2/1Xo8gQNFLj17MtPaLT9m/mE17rzjRhsHWQJ+Z591bQwF
XalRQUapjUge7GV2gjqITEeCxs5+LDs1r7vYkikaYN8J1PXlxKOYmGAXO7c7iYXlSZ9CXQ/b3EEp
gtAaWetI8E5oYq2ImWrMb0iRlUBa28UxeGvcs2du2Gf38cDrEig4Gju5s9Z2v6XVP5a5tyWBUEeX
S9Z2IRr/meGpJJq0b19JU3asqZnVFiknkrXYGCt4b9BZPUPWohhRMzRn9UwGufsXo1+9wgjeoa97
7n7e+tFZ1P/d44kBsnw69vuQTAXyyuBoiPgHkZYKjZs3IgbRcGxrA0wdifB9F2mKD/ewlaTsHDzD
4Jez5WNdq+Oj5/HZOo/jfA11lbJZ11k9l8PYWgirtBRNDyghAjGsgGuP1pu38rkWGIVdTGoLq/jr
paTLf9pLnsNBOt26XL8Mu5WSJPDqnm1UIGuIrOsLlW2r43pwnTm1vHOv3alEDdnSXRqjqle95DpX
Je/ra69of6kGGyzhJeD/+sAM5oCJYFMNzxm8kj0JH38YFIPKPcZeVhMEkpGtpJnj3k3ebqjMFBVR
fP2EQISgLl+NB6J3ydgx8YeJuPgp8aC9hbcJPndE50JBy0i/Jh7BknY26HUfRgYSRkRWr4uZu5Dg
W5xD84Q2wXLUaTxpQCTA9ttsn82kFgQ9RVPmRRga8jy6IOHgusFBFMtfglQvEslR0Z/gpwg6lrLa
ckRm7gTw1Uuq3lxPFtFpNBeredggqkbIlkUoIrkzp5jzEU7rRC4jj7fPA/Uu/KJ7j0fvVMxOHGp9
CmdOlMEdrdl1toDrjz92IqQqmBKa8JEv0VYc2JsAhvPzKrbCh0xSp4ayf65sxje0w+BgZVBT4MIf
umUkWjrP2Gr2HpWSNwuhBInBAJCy8mzN8sUH4GZhwcaW5AkEOOyoy2r3MUf/m7VBljiMqKQInBLl
3cmUmep14ZG0Jncgx5wst0D6iWG4WQloBnF6O0NT1nBMlfnZldVqM/W5PQgzfvBXvNs++7OuUoUN
/KNZsba0DniXQY6upP+kmz7Sk8F3OBgDkI3sCvGOm+XrBiC2I0bXW+L4mUOkmpSIpF0x5r15YW4k
Nus3hjLFP8El9Vp7O6WpOdtPTwR0tEHWTFmOGrdS2BgBUoI7MOfU5b8yFCN9+kLQtfSoLXurnZ2g
9zYAb/TXOBvAgE8/RbFwISQRT1Zq6K7QpYnIQFzt3Ygf9E337u9ma0iwaSPJO7LMZ9hSCD6YDHnD
ts3GIuL4KEmN1O+BL5C/W9dFdrpImucdVeUeP0Smi2Viab8WSSIOwwGi4z2wdIQHmWKkkS6yG4QW
QM8e+FBV2nLL5oe2zMUbPoWxrdEVkgRkxAzPva7Ww7sXWDLZJi/Y37YrA8PpVOgJ7OOyTroW4aUD
9LEJJ9oq+rJ6beDWxj/vleiumSYThuKUu5SbK7nrdr+pGnzjQwjCTxI31JLhGWSmt3j2EFlDkDaL
1td01hgLRKFAC5MFZ5H1SxRg3/XKRtFe1PYiM86vE3sTzSM6y96BWGDTIAOprKz85pG81oThEc6O
xAZGVdvsk/jqRNp1LJ1YrOCBokgj4sp3VzF+/QrnoHn1p2lHXbV1Gwf/rt9Q5XCRglYhbFLupXIa
f+19WxDzVgQtdvmBw70RC4XG1VyVUEuat1MZe2HTuUGqjKUYN6fjqbU70o0fInLyJQRGwxWZCSDa
T14iZ4BnIO83vse9LP1SdzqVqdetLGe1tG5VgPoU9OO4bFxLuW4TDFHnBjREtmafDf0mNRfkuCsL
Czh2Fw+YxNoW0ubwVqDHWqx6iA95pY6NrMqyD4N6oN0RUsBAILehlDYD05VFYakH8J1ByXKv4Dr8
flMM6NGshZ6+j6h4ANg0SJNOEGXrRcam4zQPhKcQ1x/NPWgremFXcKHm/Fgd9wbvEQN9sqZJ3rDm
I3tRZKngk/z0g0jkP4sMWIXywAGxHhub6XDZwnOFLKHxb0ZRm9cgLzeEkg4mYm5Bw+LN1Dft3+XF
L3LLLwI/iia+ECHJ6tIO/L7ELPC7qeX6AEWqblRQFhMF0GxIPZmolyQsse+d/1V83Ps7lz+2ViyB
hD4ItOs2gqqU0WnnrUsE8gzHAYgVlG+De1iremdSDy7ebAu7yceNchhM6YzkBsjcamd+YrKIxnFO
2U7ahNS7RvuQ4OrSfMD3zao1WPBT4gciKW28nLsvLGlU+2kSoTUCiFfSp9r0Tz/hkUt5b+xwv51F
EWgyPF+e74Ejg91rldZxLAlvZR9+Zdq75wsITVfh5oQ6+ND7ukT00F8z5Xz4cuTKjBJNQJEp7L/K
6AJt+/jRLGhyEx1MSG80dnofwma75jEWOAXJP9B0XfJqYzEbwzyoxjh60rzE1dyfk3sVLuZ9xN/n
YyLvRE6vPgZuSGCNda+sep3sY+iSh4uZw0MJK4796vD7CYewXvS7Zc6wLZ+8yXeLh4jcc+jUWBxu
L/Kd8JxyUd5HHoJLiIQ2K56CgOXPYSra2Xh0OUG/FNh6eDB31UMzHIz0z6CN7REJ6R1O7svb5qVK
PbctIo92andynhpCne4i+aRa77yPhWnpgF9WP6KcN7xA/ZzwTYTSA5833EmvLh195CUjLfg5IJ6l
7jNvYKkzst6+zsz8/mHEEI1YTkRCxUZLYL3oKX/8bxy4uq8V13qW1SO/Tgjp10d9SNk/PssfHtlV
G7q5gM9k5BZkAA/O8uOHAer3id72VmRjqRniayK/zJu0lafC5lbZTpSpxAsTp5HwUr0oBlmS8Wmg
rjcn2vfDev+W2noBQFPPHbVLXSVX7K4NY3gXlYQW7iaMH1nNtOHt52PD+cAZKkKlZ79yAfaTgd/j
8WdNFMCSukqdN8ANgHlHTM2kGSxwUrDuQ+FmNlHiq42MnOHYfyuPtN7SNu5GONQLRgo1HghYhlar
hL8iglc/tHlm85BP1z9zftsndRF+c4o5d6Q1T1MpOOac6UEl1tEAwKMN+Yq3n1bi1mx5SyEfWXVP
suYXaxJBEI6r8Xo3pbEkP6Q5n7DOhG3ZW712i88cM0M1yYEAJ2dSj81cSqlPdNlO9t+S3SDWyCPH
xPo+y2gsHw452pwuTbdA8cfG7sdH3UNNKUlEpgj3tXkishN9upQhBKohyVYfltUDNRsB+AKXEM5/
ow5pfZruWIjhnB3SlhGqjf5OIXYdtVHhFDlE/k1ntDeUUblQ5Csyc86OIHiH/pIw5pl9dA0TxYIi
WxrABcb3FzlVOHfwLejaqqnianJMI4vTYAkq/EB/gBy/ryisPNRpl4wWU7NAwlCfnZRFsXbrDUvD
Uu/gtCzs+HXfuajRG5qc6zfl11IlKz30x330Dlow+yw7rIkweiw9349pXblSV5RCQ/+qH8CZroM2
fOCwmdmingc5dwFgKwzv4y3qbrZUkTZ7AkuennD3LVcHezOF8L2oHFMSBSj1eBY9uUGzBDa6ZWWr
vvqqZld1cvAYAoh12+ogz/OL11lFDlye2QKvZdanK3t2xbMPqQQ9Qn/8kpja0UqVWFEVTwI1lroG
Su6GROggO/VW8OQEIvRMUpqUPkTwUNNL5QmFINy/uXUcAL1PjmPfPjenkvyxOar0d2Y3NK5BwKTX
s9U6EwK7oCrECfGam1R8dknUUor34atDTMzMhvr/LicxqtOkvJMAVxgSfBYK7GokiWRP1NtFiMLr
FN8lLXh5JAANVZSL+lyqOdfsERR+ngTb3Lz9hRse0P27CnpEL4vJ/sMcfbQcmmd8MI1nl+a+QEUS
jF2kKTxZSe9mQOtvua0z/Ikia7IQQMAX8tXwDIqsOcN8wNISiJYbgVIRCWXKdmksVYDMPTT9rJqn
YEsXk6Ey0Is1bqx3tUmF78gndGkaqjO7Jo7ayEBvTx9/ppkfwOIfnQRWwp8qDcYfXTXuMR6l01OR
+f/sHOqf4pXvRsakyuRFC6mVGVlSon+sveM0+k2HOmEWood9DXREmMiXSyN+DZTiPOfU7AkMzcqZ
yFrBG6O39/xfHDBC/ONyn7XfMN+Zj7Miwn8sbYOwQMnYryrdI+Y1r5mZ8VclkerZCY2CLeTUtoL4
Mu4ha6T+Zmcu/VYMDQ1eA6lfMrQuxQMQsBxS3GVIlHZ8SWWOcJaZumZRTDr4JKNf28YnVp/9pF1y
8qdamtRIvzrCeiJpF2p/mFtr8bwJz026vbqA6ziz8ZDuI6r+b2q3WFCPPKDNLEYu1sVxuVERSzjR
DT8eltsJxMwTS0wYkxvzP6IvHH1FfwVpeAPAhq6JVwFTsyFDE49DxBrcBUO929Kop3SmUA6ZaxVM
6JgPdsLrPcCaAZ2eS3YQEHplwD6F79ExC1e5a3niONkk214SVs3bC1kUpAd9G0agNsA4LdQ6moEf
bp47nBHB07lMsRDG8WJkwW05B1pmKez+H7TM0dG8gWYzZAKYo3PlNp2YkskKCoUMxCXgIcOyNUbr
Ev1TXym2GwjLO2oDpj5YWTuLXzF9h4vvYfoe9iK9O1vQYkjijYZRPebpA/QK+z4kh0WpNH+VEFVj
f9xOa9ArSZP45dOB5HEavrHXrsUXw360fZA1o2IL4Yt+yjIjMdNJafuOW7Sdm/236XSXh+iTWgW0
fxJKe4tUP6dnAkGlLd+Y17wQi3Jjv0loVi62+vK+pQKPcKHoLjBzEHgbmnUHZk21d3zYI/nBa95n
Jj3W9yLz5+agZ1OsSsiuKx7DeRzYP4a+5WLdDG4EYN9q0/NUlfzANnrPoDvmk/+4rIKI5LZH+zM3
+01KkMAS9FWEtgFpTaNj8KusDlkX8Gk6Qyk5h6XkFoZBdvu/ouKJlrCEZLfh2H2VBtk4AJsa2Jvv
3bs+zopWQnuDeWlMxkXcn5vketLGKhS+AqXXTuUW+dmDkyZ6dy/uWbhhXMEY1oxBfmLFSjopcSiu
9+NxDztNtQV30EOa3bJCCzWYR7Uk42oI5avlk/ADmdrvlHtqBb71D8LNH4iviMaO2uz3j+yuizqn
hbg0LEaUPWQ+i4Jzv4OEOoJhCXyns1CRJZuE3JjkQg1kgTgXUcLxZHlO7tcZFIUrWnlkt1XekYI1
QDAXf1GJzrsizI9aCdbBMm6TFQsSKlLrhP1bVACUtQVZ96Qh4pacKiPYAQ7HqOrb0IWWF/k64Lsk
6XSybT10SRitzzqMosP6lzk+k9R3/kZ5Z9ov1wfbLGAxjvT45o1VnN+EDgBQJ035x4WXAkC1RtKh
Mz4LjB3hg2I8J+sW6XS5MGDMRXAznmLmI3X3aqzVCORzd6XC2ctH4XEMX1eLrfCv3vHPqvJegH3d
HmpEYN/I+qKmP8sBLSZYgl3P1jIt21WdNZhiWV2yrRIVQPFSII9vWrSpgA6N0Jojtn37ljS7qL82
9VK1Tv/ks4ZIDqsJS7GdKpHEJjfYNZTICABGLqPdjDmHb0xowf1UHCmDPTrP2e9qW/zxJxDXzzyw
EuQ32Uq9kT0CikNtq+hBWpdw8YVDweeww7i+AZDUu09CMRhJcY9inw+e2GwPRvFCAX6LLihyO8da
doWJEE5YdeQGxdGl2JQnUDAkIgoBXr3qpPK/5BJcAFrqbWxUFzXRs4rDAkV6ELOrV4ugPLhwYHWD
T5vZcnr+27KmWkG3cMDLAzeXghdSdC9WGf7DiJZNHVt02FBHkp+8Y3FrCB7wKh2RYh+ISm9XAAns
8K6LZ9WIxkpUGiFgTqYETr75SZfU3Nzlh8eYD2gJU92Gp+macfjmlaQ0Zuz/rFUSuw83j4fwphwX
yf1d3BQcHwG4IjygTnTjNjqT/gVb3dxQRKzARds/oIDLy+f8yNWX1gWSOEgaeOoq7wBWTJcr5y7Q
9kZksUQ+iBMG6AvEHpRZrnvZ79s+OF8FDA5ePYsNVzcECU06nmGq/2OgWBUP3Llq4B1SdnZuBtFY
pnVUvb0s88WGxfTM0thPnGblfAtd/JcoH8yt/d/wKECUvkE2lB3Xv3UG9+QBxldl9BR67xxW/DUe
Z73Vr370+RkU57wUvmIqakql4dgqhC2i75eG1rcL10Ttq79g7ocI/a4btijxYop58cAguCESxHU4
v/5PacUNEHIXULls0RADjUTOSEHYHb4x9q9a/m4s5a8fpWCWXPPFFC/CBRuyB0BNuKJeDE1dwcJd
ZGz2HRhkDmksMiH1aQu8hETpcic/sSOXE9S1Lu3WfajlSLN29MJl67acmMCzScFLm5AsBmPmFfE1
a4f6czdbKKodEJwYN7TWI5mh3L3MggrNFyZZw+ecLqQqQPehgsg0D2469G1rUA4YbK5ctra6VO8P
jtTEaAIlEVH5DQ==
`protect end_protected
