`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ewftC88g/2hGiIYTKFto7eOuI0ifL/UD7rKxd6iuQ6uzv3tlBaHmbAzpLdJUzJoB+E8tZRZG7F9b
8zzxlzH8/g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UNLP06jKnjw1WzJvIp0YbuUcaUOi/3K7ZzDdegsT+KEOnI8FkJRlimLWR+48DYgQmQlpbtcfThoo
edJDqG8gRUli5QCgceWyYwDzK+YJu/XPvseMXI7IGd1UIfCuwAmdmfZPb6/RDo9Yr4FCU4h3nA4+
08SMGMcmlUtoVxElme8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Tn6ieaRN/rKnSb4GRHrfGvww4jqxnP66JjkVzrXdEoQVEJ8y2CBdzFjpfeizShntev/yWypeaBZO
Cop/Jhsnjk38RT50XcZ0pYFGnyK1GylL0VQpqXVJm6KC4/j6YaJSLbXwOMldosGVwaMaK1NVeE2a
85naCemgu/KZVJ+2E5ehN9VO3Mz1Ed41ZLpe8/Loz1b1FqBfSQ0n1UjeYlA2k9Idg7t7nDaELGyo
ulBjAjIJ4bZetVwKThlkRhPvtaXlkJBxnuUMnr7Pdho6J2NWlRe3g4n55wck2zd1VI6HoPRo4N/W
X3ylPiTXC1uQzw26XUaY9RJiwGvtm0IDkLcBTg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FnFP0UobP7+LyRFUFHIgC8AN+btvsw/FmHgtYFhXn2+uKF3owQSc0/5TjenOn3OIdy4r3vpUp8hi
QQgf78IxASAE/JPY3buuM8IsS2mTo2TxW3d45NocgJPusnu7NN/5OwO81/RkG0hpYZzBm7n6B2tU
5gxiB3qriyZ9dJTlQJA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eM7hmAyALOuU9skprUX4TJUaMOkyJFFybjEMrlgQY7eRTddh9A7GnseOD3RuV+HJ7zWiiERaZ3Dc
7lO2R5WZM63ATVx71//iGzZKwfH0n6q/IRl2BseRHKTKk2bW+ALQiSNEim4Me2zEXZaqHsYsEErI
343mUNBZ2Pd25YdNuulz4NABoLpBCHqPJxqy4Pz3XcPzlpPOk9BFkUrBBhHFsFF/2bWcxZ3eUFG0
JbXIhPNnSB5frF6w0Sj4HuFss4vfUZbcoZzw8YMX/aIbzu3SzE66FrrRq632TAglYYoJO12ZhrZh
+8Us47OSi8XOBsaGkhOuv94rNzlLmsjdcT1m0A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13632)
`protect data_block
Jd3+OvsnkpRTxF+k+F2CApbbQkPxuLLcsV2Mq3iiCRZlmb5/QlRuMRS4+XrqUoelCiNtq3YIO3YO
oauCzlTC7HJCPABCEDs3GX6uzTWV5dDBwgcaiaHZ1O6WGQSLyHC6D+InX1SQvzydULanl67WzPO7
5RUE781nMsFH8oW60gY3UC2Z7u2nG24+uguHjpawlpZTIZcCU3Yv3ILte3MDvdqD3aqOWzkGvx0r
o06obrRKGSgHTtJ/7RQBkugKNJcoyJmYSxQxFN/5jvuCjsrAMYDbdENCi2ypZMGKobulbpGAcYae
goNYo4ovU4V6BDJCtsB47R0OpGz1ARD/X4+QPjU6DZO5Eo/ilN77rAd3A4n2XUQtT5kbGzPNgo1d
wxZNlAdaP2D4eLkUsC1yRGbD/LsDERPDJPnOnOGcXvZNvt44J67KYrT1CT9Sp4zE9AFaRF8b4kee
N2bwLTuHGaKJ45nzzSsKp34+OHWIBnZSazsWraHijKQyerO0rcpLZlPasPd4PHvAepk2eVDsQLXB
VkpCH7lRnHQ/AZnIk7m1O2scEoBqrst+/OsgUvBU4ZbLldJoC25/Y6qat+39w/nVp9oATUWyCvGI
mGiervCqZgYrJrBEQWyVUsDccitg9om14UKNtZ5bpDTh7sqs89T87cAcG8w9bZ5g+4tFbywDls9+
+ivgLlt6dRDU8hKQmAixKRDVxmuXfWaHb/hDS0fhpJIjdxfutSuhWYCQl2vb+3r2bVCPGeH1hB22
y8QFzeH3tXf6s9sZ1F4QAgxJYPOJx+CCKzyv9iluNLH7B0nWWciD9o7qSSrPtCL7zV16PtAPDiGx
jUMD+AdSIVqABASMMMArPqZj2lvCIfk8kT9TKhGrha5NM8HUpB8eBQ/KnNlFS5tl8UKZzBrIpx6u
AWbvpqQISRoGAn7pqBx36ckETrDzw51OsmV4awMK0BMtdO/yEFKlV0THLZtWGRfvIY1xC9FNE2WM
J6iS/HP/U+yQBbYEGjJULRVvR1bvZzVOwpJsR+u2ib6Dj32AqHxx0thzGXs4FZEt4R7r7zoNnQd9
pHUv697devM2leZnjDa99ZxrRkEhrHOUgB9RtE5ekEvL4GBb95pYvHrZwNfZZb6ODQ50nl/DNjP0
mywxWbr5dluIP71772EdZTpZ6nAAOWLzZcVya4gZp+rPOyp4fdesgItI+DtyFydugn3jknk991K+
P8z4DSzL1xtxBrXwXVkjY856U8MfIUJquAGKOz9ChJgeWHXlORl33RDUZt1MkAzvCZvqVM/il4mQ
aqKmIfteeaXDl5jHrTC86ip/nLqd66HXhCeeU0hGqYrE2nGZat3Dzhfv8alUZncT1sJh/LIHue5h
257bw+gwAIS1wgGkTYk7CEyTxCKxM4xJuExzVAHon++XdeC3jDrn4ykSEMenrm/7LxOw+px2EAk5
HS72KcNSE1ZsLuLHgsaCcBVzAIOfedaPoTATYu4KajeFgx3tmG9Aun3ap6qy3hGRabsOr+YxpN7z
/imhAt9x8QZ1PfD+uehXAxiTVvZr1cRe0jSLKLpgeuTzQjos7NNBztOgih0KtWugRI1MNisdk8Tn
mix6Lu8h2OeWcTIfetl8RNmg7FAd0XisnGYsR09DVlYzjbxzjb8KJsqAODRW73KFCJBcxxZEKpt0
3E7UQZ3c/PX1NNQgAdirox5BJrid4vyWadp+aRAWrqKcFYhr5wvhS2WSFH5zCyQV+78LP2hatdSP
8d/51VyYZXTovGiH8bAWTxwoseMltGwY5NMq3kwrvquoZpQPrbSDrXNJ4of6Zhq8GvZ/4Yb5MOtW
eFGRZoUY+7gaEJFwt2LS3ZWSHeL/RdsA840pE/92b9HLs21XAl3Ptfg0W68qNwy/lpr/uoHnakLQ
RRGJdSuZjVkF+W9PssITDMbTbEPa1zWUIrHCFuNeOK+/IKlCN+uuOjimA1Ri3GoDzuiSOjOCqDvx
UdlNIQKMLfnt9Sgf/OPAK3jZiUl1OUx29ZQ0/ZZu68Aa68WKTmS15K1kHl5bea7s4WxCh1+FDv+D
VX/Jegcs7NatkTi02yresr62fr84Z9s0eY41FPcmG2NQV7jd+eGJ3YEDqKBK9hduwpZSe1un6Yum
xlxTvds95wiRwDKmJ2cuZzlkM1qjP9LQ5DNDvCpZ7++1rGXkznsrHu+lVjaYkNNtnszHqFmGQOaR
la694YSTKiRQXeMIskD18aJ1hCwsI5PjS1/lgUO0ZmhD2DFG4pVvchkgI1ax/mcYz10AbcRhJNjM
MZYHB2sibeSlVWsRauv9so0ZkUMrfnGYRaY6+Y8n0JotZ7VXJq2NA4m+yUhcg+TKxeHrs1L6DIGe
6j068xQ353ZeRYUjU4/xmdKCAv7o4ECqWwlgv+3DzcYrkJJOi9mIy7Sl+BIysOUMIFc8QfAc6w/w
Q27ztbTXJ05untNbci1ZbjlvTQ/WoXHLfBzE1XkOko/8LODJWuprnKTGIjU6jIQxTqwA5mNElsap
5+Q4syw9KkUqGdNDH57HdzX9y/q6CorrSnJbKEuKq9+U6Vlxu62VkG2CE6XVtq6YuW1IJUqB++lK
DSbtXPh5fKWR6EX+R9qDVzRiSFbeOu2sn/l4vf7FzOA1qNl8gOLwvOizMhIeCRIHsUp+NlRiD4TC
IsnTLEbIrr6eJCKf+m5tgUQGCrK17ClHKwwLuaLvWl5POfhpyMhoKl0YPsap4N0eA71/M18nwXQp
42a0YG2ud1wOV7bI+2gGPyz2IGbZVVcKwpnRM8TeZRQgZrgwr0TOFDAAdTEH9oRiw6F/bJGyEzp8
uNqE6F3LCXRcDlz2whJlhCar+ujRfaV2DWWeailsjiAMeADkG3ntWoCExRwj5Td9o9LHlDPFIVTB
AciX/kOwzVTvbIhpRn3Vnqx7C4eX+CnUGBAb6bPL9MBVtJkQx5TWR5c+WalCz7D3+d4YCcsf1Hqy
BSB+gAxlpKI1/LOqkiam/0dElV8FfFEDeCyiZB79wISRFqV/jYewsW9iClWplzaSnbiDwnj5SOTJ
Cafzus/j3I/xEeJjp0HgmUqcPPEUrHnMaOMKQopHzxdf4jQppjEaE6RfBUXRQqTZkXFdsXHI1hje
LkMP8Ok3N2EdUYdJypyghwZRUCPqB4h3PzqnRQ/QmO736VEVcpFpMB3Llm3StIrYzeREZrDyBBD4
GBhL5id/qHEzOfeIBdcgPr3Q2NhdazWgq9Jxksf9cofn9SFRa/kpcvrC/AyL7VYLBuzeZbGdbvGs
vXD9/MfH1/Dej0nIVqTSYaYjTzk3VaaXbNDK1oK8yKJbijtrOMWYuGOLpMnv/wK5H4HX4gJuXhUx
83+W7fvzCWvLoCcgq/h3T+U0gC1xTSeJcEGsoQIfaZoTxDmYpwuX21v50K5WiHFYfcFD15u3rPMa
B08qaejozWo+aU4ue/fYXN5b8na6dpyp1LmUUyNwuMV9h11dsbqcFU8a4ax00f+EZnW2TMOqjGkp
y3iZWGsFcyzwQwRaoaRndmVUmYl8sDNOQy5fVT5gZIpnh4RNjZOl3vLzEE2KT51xBmMuPSFGw2wT
W5KsIICrSr10qNwBUdA2UlzmvV2lLGaki6ExzEemD7GZrVE6eD8t6ENBwoFVt14kCx3rmrKArwNl
cP+ShwHhY1ulV0MU+yz+bZ87uy/iOJXTJPPvUWrIkohxsYxizhrLNuBAW+TBbVlLexKtC3tFN0qU
gvrP9eqDEuQtpvkFbxL4mMtLitbTLw2IMeIrMoEb0BR9NqvEvBV8Z7bDjK/QinlVYFOmJb2zzfOr
VuuEHYL8ZQF1d2Lx2WPArJwF4Kxzu0IdQsYPqShW06tIVVHOZXWKzDg3LZBGDnTQNxb/ouGgVBUk
WkAYhdaAnYVs6AaqrYvFbIy4vtR0EtWc8ZSQMQTgTQ3iT8E4yt3WVkQZsqkSkv/KPqaBHc+v5YY9
uxD6fmMd0N5mcyrRt9XHYQjOiflPyI6nyzyR4aqWu7GdUN9dnYDvGTy6ocr+VGfbMoijahMjwNm9
X8pxTtDIyuFzrjhhTrbnCrlQz3Ijt67Gdl4KIE3crV2a4uZLkMHaKpWtnVd5g+aWFiONilZ+Cvub
h8urOm2GI5a9yik4xh0E4tXodgBR5SsgmGOgWYOupsYeV3nYNI4p8MyOJqrOA3Iy5Ic06gnhiXhV
dxGKD8GWqaivIEFGRSX+7I7A15sc50gbHFY4pT1QL5+U2syhdgL2Hlv0jtReZoCAEXi4TwWPQv4+
Mi/+FNA0O+ri1kFcYk3iA0Mk1qVOJhSuGU/K94OhIddIawNZ+CJzzslp56qQJrBPZGOSDA54q69Z
qM+XshEBhWFtaeIUwaTn9nW73Aqd5QExjgDTAGZ1eEUBPWIhzXQEcE5o/sCG5KihffXODbqifx1M
Oy+IavUWUwH4DdNE6Axuh7Fks2imL66z+ZJ3uo3dZfpth9f+Aj0hMWZ9JJeVvxspKrAFod9Toh6j
2jBAGMjH52b8IcRJ7MZPOxcz9recGzcPFslnSL/X3O5enEZ+KWA/sG55LpMlfNXosUQpxfezqllg
XP/dTDa8tuTNl61o967tClsI8wGEENR0+idfc4RBqFSS0Z/Yl0NXKf+z6sUIzOfa0tZkAudT6XZL
z0bm2LsnWEzMAFC+TxERwAB+aaP/dMtQm2ZR2nAh2HYBF0jPI/aLzvHuarQ1he/47/2azxBeq8dG
S1ZpMvqf+i8bshSjf23a48Tthf5TFlD9eVQsjiSmhX7D/DHaKxRBU/PjlFu2vtkxBtWolj7qwugl
p8tNLdK3gIQ0r7hANJZ/zVZm9Qr+mUTEv9kuutZOa6/Tu7X079mz7Y6YaCjDMjVgjugzQG/H4yB+
I6wgrw/tvoTd6EQLd4wY2dgIJPxs5NzfluGALKNs1xniG/hAyGIfVVgqtFr2rg01RFkAt7vxyq3v
h1kAJqxGKWWON6kD0itjWx2KCctL7cnyY9xtjgdLYuNWzOP0J6locMNyqVJ0NHEN5uVVfWGgj5Zq
JCyFFvNfVcJKluN4GtjhVc3vK30Uk+UKiOBncq+bLJyClU7Hw01HDLJbmlFliGfImqEagX6FXCys
t7QXCeZUkxdbgx3/pMawen+haV2K2HRZm1TipTMfRiTmBs8DK5mHuqeqEr4fXfqUymScBbnDTtwx
dIAAl7GD2lZq1hdT30QjsCnroGUsGJu/M39tXrBmXs8za/L57WAK2FW04JN6qcbvuCcrVtsUDpbK
ioV44vo51fhgOYDDJmHE/CKna6s8f1kkXZougc353w9c5u8rYxaX6e8VEatnEA6PHcNz+XOckqlj
3untBSOdylQ+bCmR2SouNorkY654r+EI6fjweRwG7faMaADTyKwATvloJ5CBGACIBDC+2YzV8fXO
MuN0Tn1vDCSkdkO8RuMFsV1cfmcnS0KuTTH6vMacgJUJZbwqP+pxrBt52lEKd3jzsvyM3pv3zGPz
wKNG0sFLPke6RGjGAnlmN+PrkNr/WukS35lSuXLBpjvbpCKFNffJl5ltZ55yndsj42zy7J2ZNNrj
fBqCHhpHP505iK7fo8LO/tyPOF5P5/fwZLajYj8l4v3/PFhTV/vgVAwi87U4kvMNEfNIjLPzw+CX
mX+xs1Y+UPgXHwMsssKR7F6RZpyK1MH2wJGMGRZQzKMLkh2y6mtgoCw7aBOQTAeMA45PighOjyDV
oneppM8rQtAxUkCwrztp70F7QxCJhDlN1Dn0Pw/ZvNzx6kH7QCG0tMa5UMdqauH+8Z5hkIkCbrBw
go6ojQG85M8yGNZLkhsJ6YBMNLN2bon0dXgQKslbFrviXGa6PJiN6dShVeIAvHptpCTEDmj8a9mD
OGACB2gL0Cr0QTmZfUdwIW/HcidVGW86dz7RQPE9tKYewYFXRDc1ence9vcuu9MhvagQq7c2ZyZT
ye4kkCCW9eY8e4TRkRPuD/McjRzMxv0Hc5pG/xpCMcA2ORVYDCBEfU5QxTyowTXOcQ5pxUDubzkY
0PZf55VM8ctuxImd3qwMUgFDrBeyTbEroc9CBwFI4Vc75jes/pmVnM/1IzM752TWIaeHV1ffjpyA
eTCb52B9TqZPDbUW+yyrqpezAXHh5wepheL88ln8coXtS3IO8zCagcY6EECRmitpcMJqqjBNZGzo
MpPD2/Hik2Nou40v96FrZxq7dm8GjayK+NGYvkzKVb2B8IxzJ1fxVPopmnb2altbYr+8Q5tXoPMZ
6YQmYARPkA/f8rKS/lrhUDgjSs7EzH5N9ABKo0hMVhc+0keWhEo57wYDP9dhy9DkjrQb4glUHV6z
cvSwd+P8HI49EUeRy3r3Dg8arOpw6HmH2wwV3q9k7G2uyVOFKZ6WiV5W857ziYoRNhMS0eyvyzi4
EftNgiZazF33STn4yTXx1wXsNbKgEpbPXowyzwBJnF/GTweIeksNIIcVTMjpXml0VUQP9p8PuBns
RMu49baTZUAi+n3hnsLDbTS+UaIk9uYpq0e5elMW7G41N7NIFaB/iJxQZlxsdq9APRRmDNaTPqwN
U+bBW/D9OXoyYJjyxws3O2zufzMzl5HVIlv4nbgdqaXD03VLuiay5SAFmJnMjbkuuQGClJspJULJ
/HL6O3k4d8gLGD2kmWljEP1NPTEaYwgCn5exnKyTVSTd9RuM2HaNKjSFqLkSD/U2SXR/LiJvUXiE
K2jcGJBEXbrDBIjIlqMEBV/1PXwmtJ3WLOfQii7h9o2WxEwUCAk2+IlsahuoJ5/RkSXwsnp8lapl
X+rbIco02ZmZh+bnQ9IK2Op1w3Y3XBwv9yHYVxzG+7mAcUa0nI4GPMlVepguVF4IIosbtJvd5GgP
eQq10K3YPA+TM2BkHigbTJXZ1OLzKMCEdzMIxhGX16VHXBzBFF6Y6O4oENGI7Wspnbvbw8V/4YSJ
tFWZLvhIeCdW8LuxiPujCAGRNG65U0oEJQca0AKAOJlTxi07qsG6nQ82DnZcHgqE6pUng1wR8NIM
IMs7d3RTqP8kFST+7P/BJyakGkYJWcrVf9C4yRJ7OiX12X0nuSZnnAamv9XadhGnUj9szMPoUYo0
hGdZF0VHiMN5EJ4QkWhM9hWMxJl53C19NJqAaIgkglC2ETWEiYLKknG338P/H5z6+XC1r+mnKYa1
miwnF0JEL7i+SNSDwkNUh8OMgKlr6B71zr5gE6pZolY1KNpZlI3DwjmBTfYyLOcOdka0FnQQAWHQ
MqpeIaRN9VHE/VlFPYaBhJ6M5JR4qyuFZ4Z3KMvhd6+TSvmJIjN4hzQak7APl4X/+tjCRZORN04v
khNGNgoreJ7ZspLViLqKHS8gSjIOHQcPnnh8ElJWb1f7CrG/8Dn+zy17RFrHvQJz3yDALvJ3Oa3b
PdwRnRvLMAg9VwHCQC+XQ8OcL3JwC3g8zXEdis5B7XEOu4oH9OLosjcekHc6Fsr/jHnd4V04uXzP
vlh+NatuQRKLLykr9OkN9TzwNkr/wlUgzRJT1nawbzdEDcUH4NTmcahM15xOfD5mYwuPJ5c3vTrT
7GCsq1VQ4gJbn6IuZU/RrdcNTm5N5lWG3K3fHI4/Hqvtl/arezv4XCyF5uWMNma4wor3XuN4V5is
WWnXDovWDtViVoENHoWi3e1hjkjTgD/zj3ndmK2ILXHbRpKV8PrpvSInXZ9hdgZQXf/nSw5MkZry
yIqQJsqzCw4ezuEIEEP6o1wWE+KvtqQSdFwoyt3cVg+R5XOIcyj61EzF4h8fer3jZw5eIdTF9nbH
Q4PqXQ4TTeVjSzwKZYqyTG0cfvVZSuakmwgxH9+Py/QcwshWL8i/zsFBnBFtExdC84bwPyt1MvQ6
GWowGtHrSB61SqYdpOWWQ3FXil8Z9IoV6NIay/LRz9OvCscGJK/yhKBgtAlqAkN/GsxfAx39SY7Q
RtG3JDrjX6EmD2sa1McgtLrcqoOa6Y1ONn4JXSaGjcgx7WYOgSL/3zk5hTd32ISpPuzDpyvXK3Ov
LxTFlHfg59f36XFyInOT46jYH5rFcyKrb9Ngb654ricKH6Eq4opWBAMfnSWhtffH2pcizGSvLCIS
vVP3y+gAI3ynhTXez9VNuvHF3MLsupkDcFOFFJMnbeCxkjuZV0tefTt/Sn2RFH4Yf/4lNUJsBg+a
wBFvExKLDazFcJdoyIGCjmLq4F34bpYTqq+B1ZZNgdd5NXoEK0oseKZ3/wmIdiKzjmPkAuKTa1gu
R/hCQ6QHLrCFjBJbNUPpIoPuKyXTzo3cg/ioqjikkgHIf56jwhxJn1Rn9M0SZtZPhoXONknnj5cx
RI5vRzO7hnp+2VmM8XXTkC+3JYmfHPITeldbVQ4FoA8Z1pxbaaJdAxb0f0SIeW2cObOPzIcVesMF
NM1P3c4ADQHdMlpxPWhOZInMqDDjG0GfZJAECrHjzYh5eSxaAk9DaqhFNqv1CXT2rn+CKOIw3crs
8RuINLuNGO6xrNIQtAbtrbmpa7ZnEbdthlBwh96HeUbZvTbdv8oLG0cVMLG9oVhj2DdMdxOcOmtw
jh3BwuZ2hiu8d/Em82daRKa/tlDJ/RqgVCa1tEYrgqTuGCmwzq0krJsOoRUmsheMHIyp8gvpeLpG
p8KqvfDc24Nk5q/nEqxCv4uDB+yPWz0pBK/Ui61bksRnJUm103uvZbp0VDXK7rAbyk7rVhwOEDCZ
ujenOcOxHWt0ucra9klpuWr2sXhe9g5r2HR23Yv1IRyfUNMMFkj0ZP1ShYXiFO+XaEkMg4CUkdHz
cnHuc8HRuakoMpNSo/tRZjVBfm2CRksUB7uit9XlWtju7f5+sDt6k6KGhQ8heW6fFM/kCZMGZGPV
L9Xrp/QXlzziMxivEp71gioglQTHaC+lDipcxKGaqbDyN23XCTMCjSLgUdxnq3ZkQT9/IqIiZ+v4
2JrQXSwESe/lhzOny+n8t0BqBxIQlaPxqVl8OS4qEItWXMSIOvy1bsN/oxpp2AVk3hFuCoQgZmmn
IImYOXLmOBAiHG28CNnrONooiymMsYP1PLrP7l5YSJk7CEekv+GAomuqleU99KpONffVEf8Az1S/
OfPdZbf2X22GOccaVQWGHounyML5m5wuPUKMBmTUSBZ76yqssXOKIzfZCtHByXF777uMnrByTyhs
h41tytiHKoKk8B/oBsVYABfzsizi+Hgfbqx122IDaLWkA6ZHLc5aZem0hXnCdBVEBP6F/MPISJcz
L3GGj/SIuzGZQnD5IUu+e8lDsrbHOjchip/9oZxsQWQVO/BpRob0Of4xTWSpyBe4XMeVinTYVC2W
kh1HDjQYJpGt+oEth+dDHPEhLwuwkLvm6zpsXy6oC0+BzvYd2FJXCvaQVJeOz0owpID6FmgRoMsd
Tz7yhXWbsNnNg72wZSDDvmS0CLk7NRyB41DKNRf9Qst1Ojhna2v3oOtcFCDkZFBbOqGVLTP95dlZ
hydhvYhmyZaRpnVVv995ljDKoNL+HWlZjq2PQ7sM3BLwpvPGlXXI/CxZV07EBrA9/fBrhmmbAcE2
cZHxTc0PJ+zEPpF9PeLx4//R6KRwBq6Dj6cOIK7Le1gBeOJn2s2v+R8Qi9GTUQ6+TjrkpmXHMav6
MuvGYhKjwocIeq+NV1UQ5oPuEQsLBRIoEeqj5q+XGc1RupcD2q3fdzOUmlsNprrmGIbPwq96lApF
A6XbizjZ7jlUapgwK1+FAPLg2BHZapu4oouYkpoxcS4WylGHkGzdo5mJyAadWVNaNgKVzPDaAqC8
N1JrHx07T9FSZH1/nsrXoDD+mRezPAtRCQbXg2zD+l8+xcZgroIfK6OQ4toceK7mGuSSoaiaCDtL
R7dWMnvMVP4/k7eeVPVlFNzkDfhPRkH7s+qR2QAkRWU+y+SvRqw6VcRkD8fIMeaF2h6X5StUc4Ft
JJvQn5ae48CqKxC5n2zrydWJeJWheP1RoaJwAuTRGFXqGwcbl/9qxkjJ5OgjixDPieBn8e6cCw9h
WTHnVJiyy6VIB/hH3D96OtRvHpjmmnOgs/7waypfk1jPGnrG7we5dx7eQ+/pSKg19nFupnfkHFtP
ockrMnGj51Zup/HY+dt9lu6Ns12wOO8yfracRpQ8WIUj9vO3hgNohJGvIADj/up9wpDc8gMMDeDg
vMnhw3eCKtcpcMs0keedcDgTZ1y/EFT1dssQvfiOdzSW8SQqUYMkvFE6ntwG8eWKMjb6Gacn8xCw
+J/TAYp4Mzm8teIpTPSdTjJy/lpBsunIdnIIoiY3DV421mjPbG9WTw74NaAnymUAZAMNN9mk7dAw
WYeny5uCNtYLm49/2nnvG02rr5S77Vh8ouyu7YjdtL5JcSoMk13whZNhWtANknC9O3G6JYhHmvo3
9ZWGdV3GcgRX+cju6AWoTqtpFB+e+jw5dwnNS75lkPisLug+V1Vo4LS+dR0cextjcC2SnBwNi9kh
Jd7micrMcVJbjfPx6EB7zMqc9jE5QcjduCrjSrzO9MsUFZkJELAhSaCPFnMu7dRtdbhkWIAlc2XE
0hrSCvDp8+gct5/2XYDVt9D2wbmlPwTkjSxiqNaQxDq41C+liqPvtSI2saR4wzn40d/dPH3ZSLzL
ruGVgczI2BPFcbxTek/NHV8z72AbdNK6eICvBiytHBMqRo0WNx1tDqfdaHNLczjX5OSS4Gm4lQI7
nGRBUMHkxifFYoGS53duZvLnE5LlkK34ir1pZiwfsy3/Tiwvyj6J+eH1nsCrxMK+cTWsplkcr76Y
lix4yuOfLv3D2F6UOcoBVCBGKIubusVGgkwnxZqkqDU6pn3APUdGiHL93YtreAW7GdAPBMvm1ij5
jQo5Ro3I89x3HMzfwYKRWy4XGsDWgzucHPB4HYZUBEha/6QKugwOHP6jWUnXtvzwDH8H0bm3EuQo
v5jZFLyqnQDgtNwLLGSuM03rNb8p02QZoOOxrEDEVq9oV8Q0gbTQyK24SejxSx94hQH0bQLgjhgB
2ti4oxyyyU3OZLN27ZFyewXZKSDOzF8k+a2VYMeWCPITmvkPRsjKCf0oDDUJScnViG1oszN433v8
IXsmPxNUCEylOxI5mwzwvfPMY6EGYUjmvQSzorILSFqsJ1BD0ny1+uSir92nP9LOvmKX1GdtR4o8
+Iee5OOftYx/GoVs3gBhD9lPd5pG8EGPF7Us8xWpNZ6pMLDP+CfWc53Hxg2PM1WbMcqpXwDIH7lS
gYkuZiklMjAh0jUoH/9xAq//gCwSmQHuB43QGoZsaZfXt0YFXwcIYbQTmAXlAGSwA3+xSNE79xHj
imJnvyAknIlMQYQ9RNoHr/7N6C2+79gif6rCQ7aOi0c338j1Bm8gFsjBkWxbawek5ly77SEXLng5
/OqbmIAw+/Pf3H9i4vmposm5bD88IcpEyLMJ98fL4eKQM3o/JEvOd1qtA67AKGAHHeN9jdbs0dQa
/AbFtH9iIWAUjswrhxmyfNixOA4le0GgVaMEy3wxfbmaYbCF2YjDG5q+umichcw+HNZ8eFIPtth4
w7SyecL/oofObKIAlHFFC5neUpp7LkElpPWtx32aoz5tvCXWRbUfvrWiKGvNm5onW2utfW43+Yvq
IATubeLUde79HCEPBuFjIwf3shOuTm6o7n4fSybw07SDqEsea53ElMpjrDvys8UqMRuPaIV4YcID
9Lrf5RrsBppx4uREqeRBQzBjnlnT3li4zg1Xcj2j5HkeBKQyZ4dhNlPFAKH6E62HIfVEWrSFm1l9
eG8b9LD0bXzEQ2a2u6tJ3Aqym1Jhjic3S57jmlturkMS/zY+IADZnd8i4msNr3iP0+we3axDKlO2
ytY7HiXYzG8/+zJ0jyJhQSU3xHdoabAO+yUKgMUbmKV0TOt8tjpBdOvNzH/PrCni/SFM7KmfRmuF
Jd0vSbi4fnrCbJrwpGC/J1vbblAJXqpwoheizL6dMw5SrPXXg6NMXeULl/WnmDsH7sV+V13CHAal
9aaa+bJ/50RYJXI8dItibZuN5CsMbZEl773JNz9M/jeBAadzQbvuRjE0VMDm07xLIhO7lhJGy5hz
2/oPri8Dco/VHyzksWK1hG7+JM5d5GJPH6DOnNTuEWS+86RrTobH70JcLR0L1Ufr2+IlTj52eupB
T0/71nf6SRi+PN7aGDTGve38NuI8HzRxmSCLBJUFbsASpi6lcRulw39MFUao8DcF8DbZ1IcIZGsi
i8/LbIVz4N7U5/l0kyuLpT03ZnWpAlSuDlq2q2mbbKKuaLB4CIkU1kdhh542NvmrLB/dOes0yviK
dT99FiL2weskVtRE57SnYxWQgjOX7vnojGyJMkkdeV5M6p7fNyAlF3YE331aR/7sEsDYHxBWfsYF
aTabGaHOdvyt9iKQ6+pKk1MNc/061q2S6h1iDQKJm8Gw9Sy0yt2viBVrUNR02yzbusJ+egX9SLK2
yDwY9Lwoe+cI75xmCdMm/0N6moz74LhPKM2tpEDW0xJfY1ZVcaatOJ2zkKui4RbD7mJ2uHBIbD2C
uodeStnkVueUhaInqpkdGzrXujHxBS+2LUdbAmNXE/bN0d5fc4W/HUfMzzpYGkw5tdeFcui2pZSx
NStmVwYlpZq0nFPLM1JJVOa9pxn2kqJQ3Bcq60osPgtkfobr237DInBES+hx3Wc+dCFgzGIhYePm
63/q55HmavVANtEIPg9Y+7cnHEA2kAESOv0rWnYogek8mNWwgUC03Kf+2he1oOLWJlPzN4JnOUV3
bZq+91f2TKRFOGLRAjhzpo8XKl3mIXhxAzxVd4KK2t3UA1pjPt45P+mosyraR9QFMzzZWdU97YMp
FFTybKbVR9uiHjP+Q8jY+IHc7ObXszIujRi8Lok+8l6bzLa2VEMT6DKQUWd7oY60b+lU7IJirTVm
yEDG3ey6D3Nnc6hXyQaIQsqgLKjoez4JAHdfYMF6Fx7N8XYZl6utgOglvzE+w77+nOQ2w8OJAM0K
17W8oTtg2WFIZOK7hZcWHxvGO7othNAtXwUmK5dI5zRWXcWbFIbukPQpfKkRahVPekAGeVX72ySL
3xhV3SeSpsf8kXTVsvwhb4HWLSSKatS6i522Y3Ui2wTmleNF1jsWSme8RgfdjZqIdIOhcJFdj91p
ZQX4PIaFWmsckOXC4OKAkxRKNz20ZsOsMWa8csSS6YZvnXYYAAJdsLLXil4lbXDXUzh2dMW6iyCa
cyD/dvH+a8VIvE7y8bxkWNrls1310b5DkOySQCvgONj183tdOKG8rYrx3ViOUUoVu4WJzZ0s+xlS
yy1vdiqGmHeXlUs+c5+OW9SXZMpxMAhmU9oElHoWg2yVnPMXpaypJuQZDTpeRAW9z0CzwOuE+IVW
MOwgOAkBsjujllo5NAfaytSi9jOQN7OILvyF8aNNaq9p+iGko0LUuQFHGM3ej7/6oX7xqnfVqxB3
zx8AV6lfceg5MBoMr+ZHkP8I4fabSnVfNr244SAoYvVaCCC7EfYwzfJ3va+vXFWEzTxqCdNQbHP/
KeDIlIPDcGRdEicr4nUm1DFz3Xjl2MIYtjH1nRG60ygOuSolv8IICClsUIBps8Za1qlC0LyIa6cl
OD7RR2y1gGwnfeRsTPhJejhcVQSWayOtUrFd4fx1K6cvg+AMU5LpHB7pmKrSbPTqWvjgdGTUGxVu
/ZPjRlINJh7FvHFUcKFUQVlQtGaztB4r6WUZ99t9mJlbufuCsLdw1BD0oawG5LjJbWTPZLzEcdc6
4t/mBsXRK2GH6JbGlJv7UWSwiHfGur9S1Tz/KmkVHPN8bfycdgmX/8WsTYQshCpKQdRYPC/CjnZK
9DIiy7neNFvNbnkVoSP6DFZCYDLpMwuIPVt047EYxRJ93MlwQ8tSenqlZ4Q4TT9VVVLq5+1PkmE4
y8tlwz1aPR9gMNjrUcLvOcDTtOtF00FOyeH5QgpieLuQ9xX9yrnAv2YNieQX8CeiEycVvFh5XCOT
XolweW/XMPJ4scOlgpxRYpxZjJ7o9j6h9nv5c/OVB5xPk0rNSRHz16MOq7ceRTrOvnz7Pj+BsIui
ZPf9Pp5q/8tvaTGkVIioQRfrj2IrJa+bC4MWZadwaT5+Yf67LEkWjESut+dHnLXKRULIs6OKdWOo
3KFVz8WUjogvw08dxPmrqS2srqt3iljJoQ+DcSvdxBUgQnTW0tnJ/SqANdyG2WFZvnv1DIzx4dHB
f4wjwT1F6eOcMhfQzldVbvkMrTBEfASum8+tMNd+lHo5ozGkDWhd1mM3GoCYQHs8ZBvGqqgPAFHa
rIHpHjr+O3tEjstkZ7EhAnLFkXhtWA0wKnb/5vxxbzGhGqAzTOxlKF4kdbVpXG0SEFQ0bqOdiRXo
f1YM2yz9uxsFsEB0NIA7lBYTXXVIHjpZGXVBkxPwv5dw2F7ZhyksDFKqV8RzVamC/sSfM+o6DSPC
k+7BmD5C2QpXZ1kivymVGmUvw7HUUmbHVTq/lJACk4wY0Sjik1KjAPgh/Ai+PdRJuBNh6FnOPKuf
ZCecmgTl8qpxP6xaa0TEVQBhEUbmhG7H+VGcDnOZ0Q+UN6JUXeOV1xMwEBXzuskrwIDW1sxKouP6
vUHx57a4tLRRKePGXIcKh8LsF5N2llM37/PJblrW5kSFc8FWjd4UfdUvGPzW2130Yv6Zuk3kbp/y
gIwstAmtPU5c7YU7AW6MfUNppMM/TGpOwS/C0kI+ObS14fZR3n9MgaPW4g73y5J/P9AZL7juAAB2
Xa2jyuHIrkUKxxvAJeXDu0wNAaQboec9s0nbQVaYMruUxhJ+W7NtrhC4TrSEhfh5ShTRNFUXxlol
K58GbkhKn0UedxB+us/ceV+1LCm+zPOxbC/8JIEf1dtkPeKY7W9tNEp36Bmz9ntwPS7ij96JsgcN
INiJ7a7n5GeeAw/j61lwTQAO+FQ6trWEdX3vVOcYLHuDEvJNtnPpENNNycUpczMmZOZkCMvtrJRA
zxehLY7E9LSvbmXewijLASvCMiA3y5IQq1gEY6+j/8ANWe1eyPbZPCl1OvMFqxnYM5UQEiCnVz7M
Ykm3rFT5c+CcfxMbIWKHVS2/mascwLHA4lMluH6JCUx2XeENMTUXRQHG5ibhS7/Bi939sahF1Ci0
ZUIMY25f80HIS07tmx9ZuM4RRblQPOTwwAhBt4+ojvNZnrsrcRcB2pLPa3UfHFXGl62gsJH20VE9
+6lvcmuu0tcJfB2W2gyHopGktX3QJkB+jNT4cdGPahS2QzigOKsVxKNoFN60j71xxIv3fxDs/G0Y
UmaBgJ0/CHSlVXqqpT6v9Xc3q4qiokSTQglhhVsgxhFLD85YjOtqKiwC0BbfF2BikKtLrFuItCih
SciyCceicZQ/h6Kl0w/0Yo4J7Cs+ObPaM3jcVcYTFfW8mpKAGEEctBJWb5TALdWVWDoV+An+oJmy
RT79uvA2WC/Jtkrt01BDc1oewpHWFeImv7rWFeC0EKdcA3AP+wCU9L6Xub60jRwF2GPHIgsu6nNu
tpDIBnUsbulSDA0MdNA3iZXywQlF6kyzi7schfT7yd9Q0JqeryVsUK450j8S9SSwzEEBpDjdosat
7ejbtTmd2M9FpfxNnMB9hZNZpMqyes4CC5belIuFqkthAL3GORP9OdmCGqZ7uxzI15GKPd1x5pYE
bUfCgCRtGouN116tivwh0WOnZHQhYxVCacWl3kYYg4L5Uwird0Vcj0oBZ9hxfwgPhXJ2BG/BarQD
luLLPyhWsRCXhB+Q9dg58GPr7GMoh0N5BJiToRkByB+kmcbsgGTYhD89i+QGT9HOi2iMA/mvqB8W
VIUAMasEfqTCY9LJnYK58lct6tTVRQYXtLLSE6aB4ulyOPi5E3JMUDzn+WpEXgu0jRDl5P2OZa6F
1U6PTUxcxdK1Yrt3KK11ywc1u8A2dDOmJrDUF5zND4qymrQzfDPeCLZvlh7n/66iWfR4Qzfl1bNd
lA/mpK1snMAynpDggsSWvft+6KiWBiAVDtbdFUSGgGaNHJJC8HlEo+y2mNyBtXHSz0YzjQ5OInnT
DmguRjfXQMe5xGbia2H3FSUnf7p94B767M//w2BL+41L28mcM68m0cyAh7KQoB40k0IdWb55NBiN
oRXlemlNU86mW/wRZ/fBw6vu6Ot6VHsqLpB/8VwZI5TG2U5YI2FvaTkdaE7wuDSsFUVoD9C2d8JY
bourwwwkH14kv6pFZb3alRR22sHi5j+daUEDccOQpt0OAsFNuLAPYDRwt9REeQBkI40KXM2uRyU2
iHyUzf5WvC5fIWGyuQhWg10mT9ebhO4D5CULiIMHUvDU0uxZ1mawwc8K5W36YTEq21uhhjEqJe2c
t2TuI3PBxMN4ZxK6xoeBSkT4bXpiYypRSctQFUF2wsrdEvJM64ycldY4wlBrq62NidBjGhVtHW2U
j6JpnB6gA9xoLzGN3AJoEBWcrUczHjnXTwCq70K4y0t24rTetP1Na/AJmKDpN9A5M54lZaUR0Smv
B1eQ3+iL+GwdXdavhUBgrops/9QvCaHZQm7iJlAGbiga2r45o3oRPvepKlr/S2dzSK+w/hZ768wT
qitPXabPL+M2dLPZCa+bAP8FObQz+1PTFtptOtyJRGqGEj0qOv4fQXmYvMGQNfvQLCNEWNv2/frq
eqBVUGRv0/dusotThPzsXADSr/23gR3lY/7GoXfQWHtIrM2Q+Mv6xmcL3y7c/baNkw6K6PcXSpTb
snkUOqlfovq4Iml2ImO8NPdH+BUF7Jyc95f4sTyuWxjXz6DqHVciOLynl/FI3wKMTYaZ7YIdwmZR
7E+qsK7wpyy3y964vqHJpT0//hqy8S+zJpwR+WouY35WeHfF7t+CEL/KsI+brxeOtm4RIomr6rs9
d+aBkT581qGV388jnLnerTHjWN868R0HUrBgTL+Nheuw9Y+BLBbTAEAXDadr8MmKXvZiC4t1X1bC
k9/+to3TvTdJLJNNlm8fqocaW8Tpe5V+pH9Z1e/zxw+C5E0tGcGbx7Bye48OUE7nOG3elp1PAHsf
ioQWXyQ4Fh1WZGmkeiu6lbL/rWxrYxZ15tZ4BKOmijUHtb5rJccUf1EVfHPCOFsODPxkF1jzDW5N
1DpegHNylPWhnKdpaLDmc4yEGyBEXwLGZj42KUMSjxD5SrcIs/LZcstchzBpBZ1Vux1jXmK/gCyl
rsNvGCdTWBH1eswfltBvW6+lB+CrBXfIoPF5Xp1E47myMrWDlYqhrDduT2GQUeH5XKDMB40iB7Vh
GtXtWje/Uf0PE4xP+tbLbYq8C5f+uUrUjHlIPGFPKd/7pXteVYUK9N+71fmQTjE5YjqHIURWLZJ1
ul9ALQLnSfr7WN62X0OJzdZBTdsqJymOtPg9bUGzd8h3zk1dr+krgwCqd5ze4GQyZyOPUxWGVo3i
5GCCcV5j4C6Cfr0X+bO2QTyednEBZv8yfdJgOo/G0w4LnQX7BR2IBgmLl0xACPswPfdLRRvnwtEA
FFU0ufAIvEQq1YcUrT3sdO8hDeEhhgUPOEaY8331cubUK69B3pnA1GLlZrUboFFJiJKwtRrYM9bu
lVtoM0qDk/oEjgRmgitWsI9D/+8XlpV3zL/4jGEyxVrwwk9NhAC43PhtDryIODLvwAaBGAlZ8uC/
3OAZljGCKJpiMTAwZhRcCK3/M+pHv7GYYFPlunVWWJ3x7pA/MYANY8X/ZAIxPVdIXHZ/ERcYRq5u
mNVGyUAkk4KsRXQI67ByhS0THQ+fj7YTjMz09l7gKk9eLfH0YoDDLiZnfZ8JmPajZcuHZu0uGxJY
nfN0xfObBFASpHBVxoRrT6rMTqp3yupGL0L8jzlw3ZiQp7Pq6rW0cThXajaqBs3LRFMHiR8gwAlP
sr4N6XPsdClqbe0+pvL56eFP42f+Oddps6SKtF8fI0SXbqfZfngp3iGByolaD2oUOfh0l18txZqA
Jqji452CeVPXyBZnV5tFSsukzeJqIJ+1JVK22WKmvPyc1qrmJLYnV/iDocBLshtWK9tA3YvlLU3E
qlwBPtHNdy0iVYThvThn4lnyvNAjNCO2h15MeWa1NW9mO0T9ZqU3Go0fQtqMcpYI44R6IV9QXrql
n0TG9Agxb/B3ysNzTM+1yVE9s47FBRiRu0Bay+yudfZDbrJV/NPQrTlYpU/S/BQdB14Q+hBG+KJ9
8cCEXnAHlg3xYBiv9DUWVi0jLAoObJMQugNDa7UjgK91mc2oDwYaiGGo/S9DMWQGuJRQNmEFREJN
93MH61srE9vF
`protect end_protected
