`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
H6GIpIlG8r2FuAd8FgU+pkGot5FrvtlzFv9f9MlqpiJd8v1SI/WZDH5BuIeebblGi7Bhp0QVZRao
+GiEMOgBkw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BXI9wZIDMvc6kpapZ/GyUj62OKo3Zp0HT+XR/XYcpgo6uQCUokYHB+Vl7tRsiXKJs2dX0Tm1urtI
L4UiYrVRnMrZeoNz1Qtl54dLzTqrIx75cR3Ph1nOLb73oSr+lFls/LvOaXtYD2Nqg1ATtLISTjDx
SBftIZYeT2pGCGUV2Zk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jcaTTZsZ7pyJJ4NN/mHtelUICDg6kAC70u1BrFgqXWWrmNoP0HSXoJmY/Capbl05ifGuwtppx55E
ZYT/59pNcVZQLDmr/X8okXjOmJ/Bb0B9rZ2LXuXaJbI447PM1ZDK5qmWwADyAQO5HK1quwj3h2Es
P4I4nfHNQXCOwQ3skNRy9g3nCbiBUL082v/hORBIFtUjbaFrvY3mUKY7PDforCvZUcOdYJE8v60M
F5uSqswrQKn+/t9GJE7HgN+iUDW4nwuGl3S2jzWQg3PBbPzNCUUciZvtyg1BzoSHQmg2pJFx2MCw
FU25RRM7tUHVQwDT9ZO4flF2sGc8aL9CNvG5DA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
n7TjpsU7JP1Oa87aBcqfSTGkk/F9vtBsU1WgLbLqdQl95pWrBfUhkpr2CjIdDB/X7z0HQhzHoDe2
xrcM8+bGItZDTuc6p72MVofpV80Q58aEwYoQmvDdEDGgVJfBL6SWJNfK7d1r9V+eKRcS50tbHms0
4H1A/AS8CKZe9lRGjqc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TLp5LKB8++KrQBuJX5398jCga1STLFCflVIQgeAzSq/EggNtjbUhhtT+KnDh1A9lERtGUVFdIotX
Vfo+qg/zuwjtSVtHY9mWZLu2NS4rb9ZrklycQuMkHNTUML7Na/xrkJzE8jxGffEoKSBa/t/GhPah
6A6N4YzpofIDS2x+RBOoSbNszjmriBDBbfeVXy3kkoieYPdtDfzwKdoxbBg6GLQEkd7mTp+DlXG9
t1AercOvmEUaj47Cwuu30CgA5iTVqC6bRwsWCAHLaGV9cNEizxCo39GsJiFHOfPEsi7j7s4BBWpn
a6ib2I8lSbN1JM98xlEGZrv7hRiBnEsMnSQjTA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13344)
`protect data_block
IXnGg4iQgd5JpfJ1tTkkGNW/Reiq08pTEyFGtzVZiy5y3kFyY4KnRBHxBUgTJjxxyfvKoalGd4G3
ljFpz/N/3DK5ikIos8Zj16qFv4aBE2zkcZQCXtwUTuGDVOlB9OrRcNHbN/gpf+fmYZW65SlGy/ak
zO2m/oBQiy7Sw/Uf+wO4ZRZcWevCZUybChUMoMSVQ9rXEt7eEeucUea5n768lrBCnVHaZcqpJJt2
EAJ+8iqNCGqP/43xl4Dl4cB6lco1QS7DM2IsEDYVkEHXqxXWZeLGxCnWietkqplJe69aG7NUEtf4
+GZQMorxjpsYUOnbMvifzDLEZiPuAJNxV3yKX79JUfvuGNW9P/e++5awMpULrTBdAAb97HmVpn3W
yZ1qW35TaQc47FYnTA//BhaR9jyWv2SllgRG0AzNpj+VBKjkLpP3kuuKfM1lHAEZv9cBoMPM1tVH
1pp1AaNf6pFMLMaZ9C0qrE3WGA0XnP5xrV2u2tmCBI6c6FzkbP8Hh+owMMYfAKrV22nIKlRkD6FC
t/ULQArVtssYy59MompctwFARE8Gzwh1j/S9cfmzq9SL+FcIgS9YpVZWEi5r6cVojP3PGTS8wWzI
TZ1AJcnta5tXbgD6vboC3l5V889iVvuy1nYz0OyxmT4wxynQNRJwyqeaHDupvO8Vc4ih/JV44ANG
7yNcbaGbSRW2qAuFyuGAEFBc6PnjpmBO4eNaovFWCcXiyd7TP7fvWhyxvvD4T3QFlYlSZHsJ3x7u
rU9DX6iiGrMgLabP9+QgagB3sjJS2sY9ZwcjVwHxbmGnH9NXFxBHM7XetHcKixm9aGJz0xIakufH
twHKC4MDjR/AV5z8Z+x+I11FcOu5VFPbFx5iOm3GZ8zLLRXHg8bzN9jEDAHr5xA/3w1Z7NtEqd2i
OoHpFIVPrHgfm//AlPyIL4ZwQgGlwUVT6i5c7SyB/+oXbjnJMqM/N/NSKyfd31xEzlGx0QaRPavD
BOmI/HP80TuSKnuBvPjg8IG3MnkfGL7nyOsb/2wAq0m1Zcz6RJoPQn8mVR0IVYJL7APv1qRQfRqF
deQKNTp90ePaCNz7w802BXCZz36hfUYVBjbqVTEycV9Bqc5H35HHcp20Nxeds51e0pIaGR5Reec+
figPCPamrlrUj6bY64GLxmrbrut4tnI4PRgG1wEFFWBGcVcllYZsP49LmlcU9FRjfD2hfbKaBrXI
p2yd2GT7EFhknfi1eyA173Ucql8qZfJjPts9/wpamtRARJwZv5G415rPo2afyYKOnWMykOOf7Rmd
ng9wwpCVYGHfZtjWjmpffDQCKWvGVqrzJacMaxiAf2witgPiWyjQJ8X3bw3p23O+FRYJh4Irw5q7
eowXAjtZlMybFep7bczAzgQ37LdZi2amVvNevDg9pze+6j6t2L5giCHz4RsfuE42l2xWmuFu2ng8
yMP1P7hwcKfwBcG5GeOHE7tgPFm9HIjZXxbYbVPvVdPuJVrM798+tI/o5Ly4MNqp9MJfSg9gei7K
scrW5mODdlTbJ3rSdso+BGZMzkPTeJK/ofuFdBnFurpt7kNtLBT3nn60ZaHQy1TovoOQWtMhtpPS
AwXQgn0T07eiFWf59HJS9XD2XLmQUiQmHuBY84uHG4TCK2NTPnX64iDwR1xDtenkQj8Y/mphjh5s
o392BT3l3w/ibfBg/w5dQT0jmYscp+W1QsZ4pASASwvwE6s6rtZl8+6U/YFtVl04e2mK1MT3z/VT
bS0WUO43QyS6tgXPxlXGIOQaO3SkUwi6S3qwK7Q0limMvrmOddH6HKCSDdYmhPNcKNPYowUf4gNW
BN+jd6/rNhxkCcxSW2q26WLDTgiAQDUDTYYopicHiJIbE66r1X5eH1xg3v2h8iqSaogu2hscOUtM
kUybijQOO4krveubcrqoa8B+bL6Z3KyFbTC8Xgay21DZPTOfrO/viQnkXBmtsHyRYwvIdBR/xZLK
jE0+4HeaWfkvDAr0YsbLdHBpvxmCLwbR17Ye+/B3AGGg4iPdcUdOyB1SttP2LBNZjaYYR6xTWqvS
xxOZkGps/H3FJXaCqynsLmOZpFM8KlantRG3cL/JlmOvFrWSYZrwoODlM0eFtp7V0BEcXM68PZ8s
X920W42KdttvvXWTpyJOES3oiRTYNH24j2CRJ6CDT/fHOWvlb/Sf5QoO9Bm2YtAVRkZnvufc8VVi
vow6naSsjNo3JNKiDnBPfSjlIZtFidsy9HD4gUYDJaLVeAtbOh+9e8NHJaMIkskV6u9CxlNlbC7+
vat97FPnD3bVbPerUbptwK/0d+84zNfLThY0Onvlc6iCLHlS02AzYDUZ4Oo4CBpmcTio3nPVgaFA
6OcMEabfAyEt09ozXdjCMq0xuF7BB7U3L0IfAj+A3Rn6PBOvxMHpl+f/iceyxCAlUh1hs42ieyuR
DPqydPXstxY/XVyxiFJi8M9rYyIIcvfx3E1zrrZ7eVuBNTN0BbPWJy23xGHj8oWzG5acremv4kIg
ScAZ7PebeCrKzHl00/RSfD1wTcQnysXG1Eu2rdFtcoa3Zoxf5lJ17UM3pLLk3kI2+LBL8VT2vLwq
WbI2QMe+qEXGERlG82uP7XJigZ52OkUTAuId+bolz9WQ7UQKgw5XmWWBs0P2A9HaesD7PC6K+acG
FKjpxPopHy9eAsUMrQtH3hxaBeQVMajfr9HmH4Z+xYP33RJZXUhXFV3PrZ+D5kNQnXrefN+2G6PY
wcUNcIvksVkAk1eg5S7D6HHNEr51ECJcCMaVT+8FSOVndXV8nfYVRZ2dbMXqfmV7R6P2Z7eVLYdR
dUGXNBNIQE2U/E6EVJLCeAPZchO4EqgdBJ6Zv/4HnEOAqQCQW6UlUIl3dCxuBr3TBJQVStHsnPPD
HlzqYHuwQtR7+XW5WT+0WFBe/e3a3gvnDh1HMgRG6uqWV4ajnw8J04dN9MPVR3iSi1Q4+JfZh8SL
3ytUPWgHX5+etD1DBX2t7cxI9FbAkLAB9ah8Tlq7m99aqSZDFA1CltvAcRPV/wO6Yz0Q6qD//OpS
QM+LDAphi/nPfz2oZ3+akg+cOUM7Rg6BG6S2hmWT/wxXMchuCM4x2V86ATVZ86tZFKJJCZnHzAyG
rZ2BJDNl9IQjGNltkxVyZPIrbR96CUOrdK0BB61Jdf3/NXUKGjrdL3p9qhBzyaB49+2tD2ZTSVXo
PqdotPrCn9ovMWcfK13qZrGaGQsrsLX0eEZLNS5O3vV1HGlQfWevd++hS1mw7Pue9IIeGer8Jw/F
x1EKtA32+TdIVXhbBbye5RN8UtEnHBfi0vJjAGplS027Z+wPaXMpVHGSMbkC+KonSkb7BJU59j+s
SL6XDpWFQ64/GgeTRLxBFgfUtvjl4msrLIff3EFyTRelgVoaE/j3Uo5dVsoe82VcWB5nhjxGZTYz
dYtoor3o6e9yDuT2THBpnONfZzZ2yHlmgfHRuJI9DWgafh7Q5CHJXQjteyUnoDpsmSksKOW2G+SX
wez76/xGklgaFeLIzuZtwRy26cxo/AMxeCcmATTSXkftA1tI8qeyzx1jp20oAC6kwc1mqF+AWTx8
N7JB+s5MIxzW0nEyENA1k8wmXqS6k5s7w2plt9Auy/4Z4NYFsMbyKbyuvpunv4D5ZhaQjEzm76QI
neJjyR11qVzMAfuYdf0JVF01PbuIl/f/pUAoMO3OoKJUxsVRjnnWCE65I4sKfBnQF/6NHZo2wKi4
7U4x0upqdxWr4eTM2+A1MdsGsLyH44ocg/HZQ/vxAPZtXCPKEnNRlmRe5PYg44qjJ9v7MabqsYdi
Nj65tP50Ib8ECEXtLEO2A8SAQni9jlH0/UNcfP6e9mRv0BTbL2VEHBH2Yf68Fl0XERaNcCNvyjBb
PUjOU2AIm/rx2JE8cJvmbpu6LgW+Qc4QxgfVOIQGiCzuumuBH1EeLR4zX7l9zIOiyYbRqMxenmkY
F5TCa2cR2nH1YTRzGlGA+I7hCDA8t7iyqhEqb/Jx9xpES2jFOVzJq3Ol1SdBNYZ/2JjqpEcKLEa0
dhAgoxqx0y9/AziPltNpHhl8ugLDFVIm+B/8Z8nyFils0M/W2e4lz/ClH6fL4k+dpMmA2b5QFBti
ZwXDc6o9WMB/WX2gVR2u8Qb4lRA2XK2wBkiJUbB5NGcELaC9UV92SO77jS+f1Eze8UYT99Zmp/7L
uBImpWnlHYFH3Y8AhLQAix80C35SFKpgmco3CIZ8Id4TL5AhqTjm6unuaJ2xX/ppWdfJbgqnM9ys
zohgvwi7QoKztPA0/EEdleg6un6tbTwKWWOb+eiFc6fTdiFWXekbafsoCE4DkSwfUQVCDPgA0mkD
Whb8wOTMsZXmSQDHXerzqpoq43/pNh3aucg7l0cAtxLm1F8EiMGZxL3PcBVRyKJqlq0+MRHZuBK5
X2D6Wbxr01gvfHS9KzdJ7QJdTpP4TPrKcezDms/wzjn6x8omMGKnqCn9fXSQC9qfr5LGp8Q2HQ/f
Vf/aUFSScN4uJSlr8fU7ImLFLChBroMFFSacAJpqiRfZupnzjZ8cilWNyq2mL5PJ9uoUVuE3g1On
5B3goeEJxkCmanCvZSO3GFIP/y+Giv2YRBmTYIGPBWxy6OPT6Om9/+4svTWMmR+Ha9BfgdB98Bgf
Lm/nLILJneLAmD4eH1cSaRAQuWgC/SbUGsuJe7NoB1TjKN5vhMVFaod62U6ZjJLqXcF9ZTJThwCJ
pBtEYgVTBvkrA9D1PAv//gCyFMJDQ9Na6zxFwt0owoKP+ESPxiLlOzHTk1BR6attY+5pZT2uARrz
kab2lXMAIb1/WVuW9GDMEOvzdnpxEc22wOqffBtyzQfwJto9sAiOsEqPfc58iOwc+cuOsRZfguaI
jvoRs7w5oUUD/jC0gumypBxiwvAy4iqGA7d0ocogy/YBghfDelFOVg+0oeUqJcU2xsjlriXNL9Xk
q5uTyHGVj1lANyeoIZDSoZxvSvkLU8rnt3UY5fPwg+HgU68WnygcxfePd/BU8GEejdLbW2XD9lh2
6zJNxpbsc8SwBfAVSetD/GTDVrRqtE2/+9HP+G0tXE4/oJAkXxdieImuuhnfzkXRSaLosYebhIUm
54wm5r1/1ea+tu55MVa7ZbtLjviE3dVsbcP7lPGM8osS8jJQJot+xR9HCbbqGUeA714CCp4wU5My
vdCGFTVwXsjSQi9TuY2CUlCTlIBZ8HzsFXsCzM0stdBQcMXBEB4UBmM+rsPqgBRFji+85SqskrXz
aP0ZPoAgrdVNVdLecB9UWmSdrZrKDbKCEse0z73yhNDAGf9MDCtKn/9GeokosTlNTtHuW+TitU6P
nBK08HYqRf53WdPXEIGc9/qrHTwptaOCMH2vBGn/eiYkkk6P5T1n163IO7DAbbAC1+BBpRLnSWJ/
QesDwnB/ffIAtu0mTm1jtjP19CF3FzlAEbfuiUwWUyB42rnFaaJhVwqCmyAtHafBNIc313PbAmSa
iD+9O/bxNXm1EwaiN2JdhcYcQzHYdLMVRC6p/qfpTx2/uUanpML02uy4zC9INa5W693s2DlFjEe2
Y6/Xmi7JlUZPZP1fubaqCwHvK6Vnz9HY0E8uWlNkumLD7CK5oXCpVS/WZ384dT4OLBWwKLfAVn5f
A2lnMS+XaSjTEYjoeM8A3v20kVtDbheVvv51Z8MJW+qt6luJ8PBF6dZFGf0xLMXm1heFtwp/8ryd
vm682L51szzes9o9Xr6Bipp/s+ZfXg7kksf7L9f3n7cH81k7gF/PRUNN5Ow3mtL1x0GdFIn484uw
WW+0rwg4eKXEOOWx+YZMNblfsFbMAc6pQZAwsYKuWKPPJMkJD93B21MubhJTjWHnZ0wzVdom481J
SUXh8AYDGPgEnZgkoT400zlfX7FlNxboF8OXCZ48BTSfwb7k06IFejnC6XNyPWwzD3c50BBYKhP1
jfalN4evxlo3//8BrXTcH8gbdFsnsnBVUTmJBJsHH3NR8BukbAULGK+Js0Ep40OyFJwOnU++G2JI
TwxNkGRU4/6q+twcBfsJnFRCBthp72HUoCuka+guh9e7BzatLLnqVZ7ebZwWdCt05qizRgsPf93b
ujRqoAOolMVvUzeqGWAcuVuc/XF1BQQgEQFzDE3b/DNSY8sQF3gEsRW8l46L4lcmpfbbfB52G0zx
4OIa5b3ktaM2baqroUq3SyQ60vVWEK3fDNyD3Ye/6xJLyDASZRZ5P0eA30su2gx48qxRdNVHjbE1
TwEgi+cP7BzcBpR9pcWCjTcYRSrBc69Dqs1bKJYTsU+wwGGO46yImMeQHTDx6RxJcqZM3ra+4tIG
3N1XAh11iv1j0mHRunH5qXuZXtpXLf29aQzWZyWuX3E0Wg4EK1TRCEpFx0uIT4XXo3UwBFVY53cy
wqLu/9NCmBoVWvqy0pyXUjQOVSCPC8ThoMXR4qM2ypVsdWj+CDl1uVYfYDeNR+8bmErF97Jm76hC
tAnhPjDwueJufzXaWZmvmqPQAv4qQ5hHRzzZMkhkGtECwtpgwkDIo6U9cX5j41vXH/q73rsRZxd5
OSNYrnAgiIyl1r9Eg0ErOQ1X6CcWGysxYWTgVBmCQR6FGCqN7TVmw+IP1iI6WxG8QR5VQo9A/Urs
8THlpXRQAjyOkoyUzW1Zpd8uFG5fc47jLcSTpO8Y7mh90q0hzA7OzrAcagOL3cos577xuJSdvlLY
J61SAtKGfCoeoh/CGqRJwOonuZlpqA6K0czZyXoyYdnDmsgVqFBq9dpaeD/75Hgp3Hb03mLJZdoE
Tz+5yGTx2E5vLaDtHPmXrfvsINJP0hiObU3u5n6ixaNg8AjEz/gVwxTg9bikCkk4Bfoi3tgzp7XK
fv4NSM+mN2hlU6wI9B6/BGnmmwrPHHC/5e91XSwDCf7AbWEX3zQ8n5RgfUapANIH5fKGPIREJcag
WWYQdTLKVAhUWnFGwNwbIfudqPzAvgMRon8Hx0eOG8MS9luiAxYT1caRzyT/B5UMQm/bkzT5G0lH
nAbDCX/ZbAN7i72wdVk/FaaKw+cFEdSbwu6BTZLqEVN0w6vBnRsyPIvThJXd8vD4cKLgg5cJCh0U
8O4H9hxekoSPvMSA0xLi7pltZYgQjlpD5wJYf+7VlKzElJT6Btus4/ouuPXnr/FZ3iC2KKqOD78N
3dezduis64EMQxnCMvPGQYYQ22zFKvyZGBIvKPUGfiK5xs5ZOkj/NAgY3LXtZ1h0bgkcDeSj4QEQ
tx4NBDBlgoCTX6KZ09eU+9dVoleBpBb8Tqk4hSigZGsVO6k3nGUaDiLyT3FV937AL2oJWmVPMMfV
HZF0dTDqy5CouoKHGY76QyZKV0XskiBeZkvBZ/vqK4gO/2F/HiVaF/VRY7FEmB+7BmsmO4KcwPK0
Io+1SbHE0WqcIJM5bhiKz9IcVgKkr6BjGIQ6Ka+Ryz0ri4vHHog540Xl/OPVxiYUtMUpsqIQ9AQX
uI2ad6WGsM1RstQH8ywnFqq3vOGUX+UFsT4NtuWH43w5PNtM78iHeNSz/PJMVM9Jy4ZTrWLMEdMh
i0FPdTYoPV7cHsUcqBV7j6YV69LXkbh0WC4QRzob1o8xu+vkcaK+0UC8m9gNU1NgMjTxl6ji5U7d
r53vwyaVe9GfaPVDg7IzM9Or7G0Sj2QxnFuM33tRzK6oaSr+PAyZZ5i4WaKzxkWkkMJ1kMzdwjQV
I4fLPbYG/Tj0iubsFCNBCQDwUkNpZjKu9PQ3vYGiYQhhKZ2tYBn88vxprzel0YpJCge2EWNbBXfp
o3iMJrEfuQ2advTKJsHloU52ZHdN36TbM+bIH3LwKr7Al3jvu0qs5xiQPJSwH/1vo42xe4xn16th
nN/Ai0NXo9bTUrHF1QhRayHkVzlbdw5HKEK0RTxP+HP6oKslCMB44ifhwwlu1Aqodip6mMfN25xN
MvMmFQjlbF5Cawe/GoRnJi78cij+KtG4duWf0RUA29fklQuPn6imArQ9HyWyd3WiClRVgvxI+ZlQ
gP5ETut1iobSFp5wYkEKbaGAyCMlBf+2THHbfcCWHAo30fv9PKAeteVG4jfZZGKNX7D6S6vN9bli
b9Buq4UWpFI1jFrZtWBPRDR+v7Ed751itxepp/P5acip9rVUKdzAWAKYyxyAL9Xcon6Pad5RvUUx
RPEeSoIS+N9iU43vl0/uzee7mX/+7w9sC9vxESqvTZ+VyGKiPXWea52A9jisoLkvLQo3Ph6lr6S8
rN8Ri8Am9u7phb8DdT6FyZTYbxoXTuNRFIos0HoVQjBa3X9EoL7k0kqtZPznPE0QruPBNaE7oVXH
NS407cnk3yhwb0zBu29x0LkAKPMg5PDFCQYEE9Zqo0O3KLItNaBDiPHTWQggGqGn/cLQN1XmtEu6
4q25VwK/HSYBqMgQINdXJO/Ej7rAD51TrwrLgm6jtTaCR99YJapCb73eLGMxfhOuVc/prZ/FpMHj
EUBKMsi33LkSMDcjcaaZKvrOzC+wftZuCAp4Vwa32D8qLJtsYRcbDw4ws48UUm9kGry0e8sd2wiq
CzIhRRATaxSE8zb/MfkVLWMkqCSPuhdN/djrXq5l2MFn3Uk0yA08ccie9P4nbFVYOqFSPCI3R2Bk
AmlOrsEzS+VkPzDQS1ypIa5lqftt76tlo2vbF9EstFdsn27rBPyN7cMOiR+W1HwDy5ZbxGuuopnE
8I5Hb6ofLC+/vGI6brVRf1vjZtiXZMPLtNuhEY0pH8qFyMOZK6PyHusd8562OBTJfZH1vYZOhXnr
fgJdD9hJHKphBs8XRDvp75/7GKVHdIB46XmozodOYAbYtxf1qlNubOgqdOzihSS/ziTpo+tdTY9u
kfgFAniO7hXyhkQxecN2oIFY10ZYP5i6G0OzU/eMMIIIKEBRweFi4vwC/8DCNYqGp6doM3GnBi2G
CEbasOl3DW0VuPbVv81vCi+m67qk2Hw9tLMnAPvRAC7Bpm85glbPaCnX35/j4i8bKlBo4yxd6nXL
yo1DrBBLp8NeWWSZS7hpuywIUQpX+CtupE5aYFsX/ZNZDHFaM94R851w6m8hB9FVebmnU6MFba5s
jOkS+4vUDtVVQ1oPW94Fu0l7/NpnsGPQWXkUtzaz3GJlQzxciVUgr6tDleaT0aPoaeDmtPDgU3Qu
a2sbHvuW/q6dQNDeGi4kbz2hQeStF/H71pupZ/nQuQFku6D2KCAgI+TqoPAguzh7NUD0cxxgx6Yw
9cM1LcQCBMPXpvHW73BTxA6T9x6R9CaTJlHZX2SK2w3Kh6FhW91k1klA3keD/ikrSKMmw/urccuu
k3kcy+50Lu50K/k7bh1dhpcgQdPapm+IcZC0CBIS4YSfn2g0MtrpQ2GJUVRFqC4RrR5VZB4uU+YA
vzpVDML92+XH8InKsrSTsG2UWNjFzmcpS5foEuvNxy7DB8Nb4e0gzrV8oCPjx2pRxMn3ZlH1BKSU
iMe2P8CWL6qgMApELIPY9sU2cRZXH824Ljs8ft8si8nEswDwFps3nrvhrNmpnxw/4V6POPksGQMl
Kwlpa8NtFLBrsWvPoEF47t2QYDPg494XLlBv+MjK+ubdD2pNnjgS8DgPoRs2DT4+AkmNHrMD28zB
/yXo1FSmLD+XKBDQx0q/gFSo4apSMSR1z2v8hlsQQG4f1aKyZSNLYZGmsF2oVkNcqGImUosUrRoJ
MBCq+/jVSMOoLU597se6/6HII5HvACQvEbZ8JSq7nuFJvf6vzAEnyyK4Duyrw3DF0agPD0PWA9pV
ECUPQdYpih306eMI8X1auqoVnDDbw8Qhh4zZuliT6iyklz8jw2eBJzx4Z364wyY6FJxHYNFI9pjV
FOXxX+B3aJlYNVoCwmSfaeaO5RzOaOjL1R8wrswHndYdQcAeafT/w6CzXJIScMp9TYdvvKn0p9DX
PGsSuKveqKDf2HisHQvp5DrHAydNwBYQu+i8HTrHWQEJxZmugkgMOlzlKdT7DibsDPjt+t1+/N2b
3t1aLkZWbpF/rG+9OxdmQD2Cu8EkFThoTvrIAAV6GVTFbnk53ZfuCs6QXblNr3OoJo8gUiKUs2Z/
YF3anAmMbhANfh3AtfqpjjjFl2tKlYPTGqRdDiqdg/RX7htpsvCY8X7q586mL0bOvjuuKUbR0qK/
j1MTyRSNYfyqdcUUKtSBv9jky76Q+wp5rdyObdTUapXAXsFpcyyURrQCiSpIyXsjhDaFz80g3TcX
Vu9BuWu9SAi88+/KuTSej8Jh4XzQfaHGhBf28hd8gMRa4vHsrqcaOGhuYMYiFqDp0VUBszXvtdZM
5tZfhgxXLuypFi7L6COgrpafDgoxPAHYaUK5tZ6p/BNzmUQpkunoljmeDcuTIfTuYOmuXusgCz75
XCX3IHQ65xrjDLtAbV65/2l1THyop7GsKKF3mztsis3ZqE/Aa52fuNQFoWAf/LQ/sD9LmopNMDZG
HCGw9l2EM+FKtcf2Wqj8j9QHwozY7SAYfBr/DjRR+tFco3yV9+g1MIGOi0eamU6lx3SwH57pt3a4
8DqrMWEnj1xzMa/TMWIGw1cOJzaJhkWDA30NVW1TmwYFO/ekJQSuyec3EYiTQ+ZSeiFKaonA6FB5
iDrja0vvcb3vHGiA4n0qM9vQfM6EwNuc0Vp5XjasYiPpNKxx176c9zYHwqgMg4zHKUagXR5J6KxD
xEB+b8WdnaoFXcwx/vDIVGcvsKLu1I7npN2wC4uc+Myl8Fc8LURLF/BrQk4RqdkmupUcXmrhwMkz
7yF0igaRJTF/NMKBnlhV/yfmObcJxH4dp1ayr+6sMq4V7ph1M6A5wf8k+GMep5q96oun8eSzJZat
CoEoibbfT9dDgdV3j9VqJw+uulIfGKweEitjc658rbvoMz+qQhVH1856mo5CzzdB30Eiwie6WxOJ
CqWfS4KcLWOs12Og4eTlpFBdlxU5XZ0jTiy27LqUoAET9MGey3BWuwezcdqCFLnGz48JpWYRCf/o
BVzwwpq6cHW/+BM0DFA4k8HfmzMYQPRm9FC6O1+QRoVGGuNz9Cv3RESTvj2FgbHgt6q4nvYanY17
ZWADcVkZlnfS2fsYigfmURFmOsxb9F4v/7Jz6cpklpQK1RIubqWPgkmzWYVV72MkPCLCw5Dqi0T0
pPlJ5R+KxVz17KSASaEVeeNOdc5qGXI710WYYG56KSXF1zw7A/TeUaJrwfuWXuLaGQfXsnW8IKZm
QLHcg5mCsf/I89D6uVSbag02ExyXZv7VSzzS9cF9rE1meg4KDsieIiaKKB1CQe+jcFPS35dzeH1M
PRhk5XIwsGQqHK8l7x4pQQw844SHUPjYlmHSMEbSg1HEsk75tMqrYqVdF49L4eVWKJkjZupT9t/F
1KLuhG+j/RzCRSpt2IphqTl3xqyFvEVwQUMGhElflE40bN7L9cxqDFCLJ9yI9IjrX0TVn9Vpw+ZC
GngDI1o9X2TxUNOVsPYjtaFBYCvqu6nfMv6jrkRhKgwMGvnmhs4Ymk+WE67tcp31RqHoW//Cknom
nl6YU8Z8z6IUf+jTiVCNoRpfSpDPEsXRNbM4NA9O317U8DawIVSvh5jaoHTu8rsGu9EWs/snWW+8
gANjx2LV6vl1OajBosk2Mqlm+RRnjz29cAyn+Zh4C8hONMiQBZUYNWq5HaHqqV50WuapCHc/PiAi
iopgIZ5rsjEMt1sml3h9uTb4rkphzMSRctw17mRPio1tXiEiAZLARACI6IvhR4c9yDgfDW/kGIvi
TTMiISesecclR6YwfNdBbm+1ibLb//Ea4OsoqxYVDkAaV3kcSshH4lfZRmFj95IGzTQQnXeZtZmE
Ejya7ptwY6deFWSvfQ+DihZgXecCFaaa2xsgdL+2R4rmyqg+KlTju7m3ib/yI0U9PtjcTWUGmIxT
PPQQolpy7yj2uPAKheqmJknk4KjRUcBK7Y6c/Oc9zpvfjivs2wejg8ZX66GfI0LyVtFVBwmVGB0s
U2Wq9E2Ji+fvRQ/gWk2/a86/xf/grADEArilnqngaardmKDniDE0Pg5lvwhrcML5OM/F4/FQ18vh
kuQFpEomsgjlyBsqxe3PEQqzHlfNmlHuENgpu96vmNn+YXVsUgVd0b02g/T86w2lXOjke/e7axlt
5vXuJ6oy7+UwIal+qpUJEQsDWqUoH7SD6FoicC5m/hyL0CNBKhlSgLSJOuFD3hRK0kVfpy97pRqw
Z/HXC2KwNLvA7TOoNsl/SfgiV7IvZao6AOPEVbLRVIWdOnAU4QMqLhxSgIvmzDDYc25sy55GEE5W
/xxMdohVVHD9YNE5sFTbInzhsJjT4kLfNEI0mV2H0UW9LoNT6xv8ic6+aFCZsv/PIaFQiU7+lrDi
F/P7wvzpkGjY3lknEHA5LWsWmNznjlLaGuoErq6BtGrIAHLmIWlnGqFL+O5zsjfueqazZxY5saX5
gdzrE1lQH7mBuZ5wHz+571Y0C0Wq63Dxkik8AYX/tc3a8MRUqA3OdFJPhMhm10RFhMV1Bvbp0Mi2
bQSFsiFXi75Y3G6Hqz0Oix4UQIbBHQG1ugOo44O83inUHSzl02/0XSNBGDjcLt6yemIBx8LsgVyH
KSy2CDzp5fUveELP1F/pVlps9cAWi4RRC5Kgi3ocyS9ecIWBVJhRHYQQWBNvqOLJEHldSZePOOtc
0psSi7ifKoVJQy6Cw7ODMnCmyRDurWvOmwapAXggZffC/w4ob1uy5o0b17HuUOBlxJvHQm+x69Jn
k/7yJEWO+X/7RjIQ2elZiSqjcbF3kxjuzrW7qvHzL2JQZjwqzzspAjd7vb3PsjnwuuGY5MibDSpp
o93J1icMODTZnVdNAJeKUy0zjVl4Gd6ijyuTwKRdDCXWSOUO1oEhZ62FG7L+2IoBm2hMDMbxWj6R
mVkLXNN6NqMOhko+l0AjOO7s32k8OpYIb/3XelnRWmyng3lyKJXhufLIqxBv0wMMt9dRpi8d1aFk
+FWLwSHvfwS3bXHyLe4gNHfA5pqvKT9diSaP+StDiltTxQVxL23lc93Y/0DkTUrd2dc6DlH48sOL
ZLBzHMNGY8Vk/0mrLylC+v0dI1RHZX7N3kwserdE7xE6jFV83pw18olXHUozEXxb47UWAZwpwSMT
1+7XKKksKLBXLlUmATz/DahUH6JvIeJwtXN1AfsiYGPU18gMX9NUChtR78hOygaBr9kJNltjtsDB
ipqZcqNl76STLR9r7c9Fnr9/Z7JwfTZxZ6VKgpOjD6zqCkA4xswwyNWeQULmb190sw2ZUHpvXsYr
L/IoUmDbOeqWRueU/kxl8tJ5iLNwb/D0xlAtQxhmwm6iiwkfN4zc+Ujyd2fNxxg8nREUe+W2TnwN
KYandu+2EMNVS0Y569bxXokvnTXwQaC+XyuoR0vxAOXiaGu84/M7NneZKHs5Fxxo0yFkUJ+J18Ky
4/VzXBrFYKC0gAQRanu56977yMT2hVATNcn2ll8ekpdja73lnSWRaBGQSifQuaXb8ms5eZ+TxCyf
/RtbHIz5YWXSCN6HTZNjCiQPtHe3+cCiIK/6obqI6n6zuy/PaaFnviwGDDvZ7mdgt7/Hw77LHHYa
hWgHMiSyK6035H0rHt04gLmAmCP/exe5JTRQaix58qZ1mphKmn/snjPvLIrj+aLgu/GuXgpfnqBS
Exjs831fnWc7nFdX9fqDMlFm6Ka/g56YsYODlm14U6GypRA0WQ2E5ByBV+kYCNppUO2iKY7RfiVR
62PIYCJ+o7JVjQDbpwtjCAYYekfxxGxy9cobyp+MTQIKpGHdgXnLh+nXAptTpVfz8+6kLh/YAjZv
8VhOW9MB8XqSmfwOciZDywDXOyq+w+0K2UAYtFDbTZd2tAw9/qLv/9444SAzY4w8k4owwnP3cRyk
9rP3soV033tzRUfJaFrhGsGLdwCPszaS4wXU9QeP4XPX0GqAgPLAUfy7fxIh7rB4gS65t/HuFaY8
9lmg28iYDPc2Aaf9Idsjz7rVdOsW5xY6csdnOgfB6MP8Iqp5Qkk0zJ7Cq20QRJE2H8+WEZPAo36h
tf/pz9MaFDHf355dZhfZYAj2mKB4ELlhtXmXSDoj17L9ZZszjZrS2kKKRIdKxgah3T116+9xXNs8
naClZ5WrBdHTINadgP9C37x2cRUYb/Uc6K++d53H1t58nLxmUrCNgF4OOEvGFek+REnsqYLYxouU
e3h+ZHa2T3hSd+djQ8dHFHyCrdX+0vzgd1x/h+Ijk0EXRxVmWF9nei6BnQcwnnSP+k5vkNrlcajn
NkYaiEx9X0tX/UXEEJGLllAb1Mub+hnkI8ZkTZpFENbgOMPp38NJyAAL6Hw/7n2yjezPe+DCeP1u
UAWhNz6HAiBRvNEPP1lt8ofJ9ajumOsgWqTwsngIudoYRtBb5kiDywnb6Q2WWgGZLIvqhzKrhkm9
mPWHuQR0Grl2kNlii+0hwJzvt2KOtabZyDOg60P4nznr2TfII4tZZ6F5C2tL7J+jAgdZXMUqCxSS
CTgnSePqPeYYg8HZGFQLN+z6/d7bJrF59m2QkVjg3nxHyU1t1fvb0lTeOBEI3CMnt/9WqypipBud
RNnqKiMVWU8+9gxczn1Xvuwnb1p7AMyXtnffUouHZw08bwdrZPyTaLdkRlK5G1XKWTJ5GPCN6WOo
bYsH950QB3DEmo6LF+Di0w8yv0kgUsOE5PFaWhOFbZ4Tq8Lj9PCoDgv5DMo4BQ4QEweTV9QojZEH
SP91Ri9OGAko3aaVOs7XHfYqeQ/MLbtDdaPXTWSAKN7z72XDh1Y5xrcX48OeRKEUZ+SXEgBfvxEj
iXpTzTbVlv5SPlPKMHBXxOaKxCBWg1t1jTnhn92/uywsBTl1Ah9bwFr7ZNuiE/jYPbLPYEWykXWf
9AUsx/ZM4KGuxLbKO+oDqL0rUMca/fN01gsdKXv8eT6NvUDF8pt5gQ1CXFPVymE8hD6HGrmMwaT6
gAQKhyDrjFxGapZGWxP4wTCWIXABs2+IDpky7ad5l8EO0j4o+BMgiTfIYp8KDiL8PLvQbn2OGO2K
13/+aNWHSK2sxKidqUJKw7suLtWi2J+f9Gw6jYop0nfAI3CXd78hrSjyicmiKDQyg5p+JcpQVkIb
zPglAnSITAANJMmBkHga5DOyv/n8lJfqjoL8AQB83PuVkQ8iuqdiqO8zySoOJzMtYb8QKqK82PVS
PgnRAPfGRNxDekgbFmHbGN493sTlNT31tz4wXvj3XlRvg1LSdh7x/t+80vtdlkN2C4CX7oV/WB9d
6ManIQ40YznBG/Ny1pplsRM4uqWL+rg+wqPZTpTHsLtuK+VNWXR1iZ0L51OdsraV8rI2L75yCogA
9JrJLFaqi6K8m0lwDS94KspK66/DPNsKFy6HEHkpVQaif6ufOtKjL9FnJ9+aTsMsX81esf4bx2eM
jjYlq0NVZIOi0wzo+o0iBFcsyOABCdbq545OOViY1xZ8kuT3qKmKqkYOAqaOwtDRgobMDXp2JH9h
ExwOkyepG7032icYdRYKdUUYjDShTWD+DT0vZQkGEYxTStvfRpyi3Q+dT/fe9yCMBw2Yi2D7Ptxw
JTdKZmIv1GPMCBEpJ6WZ8ULmlcdMONiXTtJuuJzPR5CwRER3hjfZW0C7UnaprGDSne7KLiQQ/GpH
HGOmVQv8hTF4G209PZrZBgqWeGZOnhdKNCJxI7XCfhRMHPEmTqnpI0aAsJVSSIuRaAnuO2gbPdtz
XnIR+QXDgOpswuYfqU0496Stkc3m1I7/Qcfm9RNgxC4opzEP+6AH2NOuhpR03ZQz4T8huOhx9kAH
2ZBewqAhwch/eXeDasfoxsTJFTpcgCXiVyyNp2w9Z6v79ofvTcWEz6pmMKUJ78EvE/escLDaw9la
ATeNUTN4/vTmE+LgmRRTszu40GDPXkCBsCzlKQjG8LV4+N2G7QuP+s22qiJsax7calETEEaxnUo6
wkwINfJgd4mrccn9TfPGV4w9s+2bZBN2OUtFGY9s+mwCbsyk9in1it2PMwrJ/0xbg0WQtVfBA14s
j6xDK/c1dmeT02YIXudjOVPv5cVZBiAFv9mGghoIfW1+IvgWXIg4tSDoGoL6UW+J+nv9Ik2e8PHV
NEfhuejrr3zyMZX8OjV27JkuMAPPO3jLE7DdqQ0l7i9s+bxbSB2CXAEcV4TaW0PfTq0degI81YJM
eZlSqLnEHxBFzLlTHQHHFreapuJgmkJx/0n0QJs448fgUIfLOXvVWQKtWxVlf4ytSi6e7o5WRCx0
fdO4VRqhlQ6Wc5i1EXvxpri+fUtdCJdhE8cr4MXfLtCKXihU3dx4A9wi2ErCKM06dB/3Gwdz5B5I
k3PJ/2hM/99ps46ZE8lgO7x7/FlECisei6GQ7OW1X7K7ZCQQM6A9rMX7Wv8FLpJn2Tdjfe6VQjIq
7BWxnyEx7LmEim9lXhy7fQO050yDQPAejtYMQNceNbWC8lnKOe918MngJ/SY0sZ393qDCj67FTIy
GwvGW+riwewDo2kN+TDy3KYDs7BKdMO7RiE7gappLO6uYmiROjmNgGuaspCIv6IR8sCOw+C5dZ0z
8bBBqymuWZY9uDJphYLP3tviH5oV8IotjdoBfGJ3yQEe/90A00dDt1R+hpHp0bWTUE/ivDK16sG5
AqYLkebqCHZYYJRb9T33dmWSrBBNeKKMM74SHVr64hDBdQ986fe09lsjmp/duQL3LmhAOBDJBi8/
w+goAJpf0d1MfzudgHEftMLfN84vc4vDO+Hqmul8tA+Lf5u5gqeqdhMHTikWlyNXabh4SFPCZenX
CoFj0PIMq3HClSoH/pzGHwDy/TYBIASJ2+8EInhJcEizyCIijtWVPELvzlU0f+q09P08jDTR5OvM
dPdNf8nrxWFAhGrb0JEcDS2yq5kRYbXKDkHZmbahmsRPDU7Jbbro6zjqWJeduDGp9Je4UWzrufIo
oK59jdUZCaoOMgvB1CkZl74EMCp0JFQDNT+NeQM3xqcgnBA+Ia9E+3rjwXnKpnCbDVBMSDITSEh4
7ffhTSSibin2jqSK/Q1u0yo2pOrEuxnyXsy2w7wdAkJqlPYOJ8Lil1cAATjBaag6fUAt9Fz/85cU
neBOFEBlYPmXTk7Lhg9e+eQ/hKqQVg8sFFl78HKgZpn+QYgtR4xqamGCoLtN261cBBrCQ65tVSrp
Lu426l5OwS4BdBkyGEnG9rRDdb0p8GOlAqI9ObJH+sIm7RC2lc9J9i3KecrVwTvV2gZL1oXtjqqC
3+47sCe+2tJfVcyJMxW1fhlQcEXHdbWGqoEZELkYpYzB8Owi3DSH0VI1PY/3Ki/qhzP3Wg1dwNW/
5y5wEnY9fErr2pyLRyPyRFwu+96aby8MvSsqhaxT8lYNsqCH8Ch3iEAacVOYJEHi3zGwCGKM1eJu
8echTDZVYV4GNHjgbJgwrsqdU0kPyEC4uzdAmzY8v7QpwqDT8RuksI9Qu7tHRElTk7jPHfOywNQP
6h/feB7jtb3D30JvJg3GNGZKRN1voB5L8leEkhEXqcYB95Ocm2doTicx4MsGWy64wztTueW+Hx7Y
Cfv8tQ75qzu3JHBJK33Yy8K2KrWF5jGEDNtLA7mCLSpdOyLS5y0hO00C6QXrESAb06iJhYGlmHnB
6DtoPCYjVGa/8mqZ0grpZUHOKrZSkrFxunSMYiiw392IbZ2CquYYVypO3J7u7awUQzSCD/ikb4+0
m0ToIMOFmMh346Pymc161rs/9ajiZPZxCpQ5bUnaMJnFrCqOF4H9zweAw+QZCEYVIJS2HMKIuU1t
rQy+zw/z2mU0xQmhODMBCmn1N6/XsLHBoLQlcXZOUXZqUjSEz5DrnrKnTe2Jwx6KUUE77Bm5J5Dg
KxYUcxtd
`protect end_protected
