`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UHQziLg/+oANwvV4Dwg31oc0UVeW3GKWqPV6GFpq2bqJdM7fFZvUqE5BdIM4YQ7/vDqpSpAm20Vl
bab1EU4hIQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JmWujGCy0NHz0xO5s+3XY+zXzGHxI6nRAyOs0IYWHluxxYor8ffMio0URuru6tZY41gqwreRMcVB
VblhG/vydvV9WUG7TWXh5uP4O5/srUx+n+tmlkRtJhXbDcyYitNQqzw6Lvt/0QzFuErkGuiK0Pif
FHZvvwih/lSE0lQ5J1w=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YE8pnDRRJQmAAgdHZ0se3zAjBnlFCxrxgycQL5XaHOZRrhSqIoHcbzCjx/l/0uODTO08xSYL2Erx
IbmQ/u077WzW5l37/NrkpBcrLcxQqVAv+L6Y9m6/LeEdDn13ZPwGXiTwP6l/z/9Tw3XHDhFbLd/N
iW5hr6+qsbipmTyA2UkDAyIkyhXuY9Ws8ZYQbXk3Af1s1XBf399BSIlJUPO+5IFmSixuFJNxrewf
+8CGzS8sYsfacRs17XLD2BL3TkN7LJolMcPo5gaEPcG5ABuvzcUuFcZSw91drVNbe82pzBVPIQYA
m6gc+CPOtdaPAruGBLCCCfHlOfZPlgKKPux9hg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yjFyJI8StX7GAKaWiGnTzBJ19p+jknaPne/1PUVYyaxgHPmYcpdpDfR0YLzFyHUsCMqa5s6XGk+2
Rq5YhK94U3PfH/UWLZKHVn9smqRoDICWr5sJxNGwkGOLwSz2wm6GcQibvg4FFnb/KRT28Ghw04TR
pX+aeZZ2llkZHq6BnpE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SrmpT5iGhuawUHWW3q4EqipmZxi9YJYJoTDR97ey8V7VPwtG4XSVeTRqK32Gl/WlGI2wM/taPNo2
+0eDVZJUYLTBMxYeuZawTDebbeKogOz3VJc9pOrT+vYWTQBe4ZV7cL0Q84QirUI75VLWFG9kWQRa
jo/Fvs4OCgQcUmttYORY8TsUhussnXVavkxgghB+qt610WpL8gtkpG4bkCQTEl+DV7UxRX2slEWN
zMibD0nb+NR3YNSBc26xzJ5BbpGpjfAelYSQiE4cuRW8/zw2sWmec8RELgI+V7VGR64L60Kbu9H/
UDenqEsBAZRQV5dKPQyZBW4X5KhNXwtZNb9zCA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 36928)
`protect data_block
moKReIqzIL42xhqt7IP/q7K/oIRP1zuN0DfZy6xK/bfzR8xMGToBtj7DzSUUWu2PFpbgeVlfnLg6
1Y4yLdO5eAyLxZ1h/JLY2BEHJY3UJMElZkAHzwo1Dk7uYRThkGIHlQGs854wjb3ewwfhVNPITpki
imZzcPlDc5TrlJIk16Fmc+sBDl3UUr8FSSk+n1SYr3d0FMvGbXN7HFIAMEDowwesE0p5ffTxyS2h
EKl4xHnZiEtypKxQkDftVsG5d/u1sIupxa3BlJdBkfTGVHA82Ql8Tg4rISExojr/iZVmcSv81Zcb
dFVtw6o1MynU4xYy0m2wpsOEMoydEn4muuERLcA7XUDQ/sfQRrgOawpFThNHyumcDuXqilL0wFKq
8pakP+X05r1kOoZGJWFLULB8SEp5Lo6UX/EWhWriPdUnvTCl+P/Vekv4ro3YotqGYywzT73BIARH
CcRCeR1WvPKDmrYZlHlvQ1hGs/bRGxoefvOexN4zePEDJ6GxZ5Gkwm0pRMNXyD8paf1edD7iNQ2Q
q6WIsbtkH7q4QqxwtsThe5S+mKtiRISXfq1cZRkFtABZV/n/ZI+JQoqEw/u2NXFbHL9JdCzgEe1t
CEP8TZRzKILOziPJrZQ2Y2VYrNAXXfl2wdFnoyH6nj6D0Mo/d6OuCMo28wgoVt39PrlGAIkInbch
dACoEnZSFb9X/gUGCuALntNNfJakNE1WdZXVo9OOdqHGzPB9ZZcdbV2hVJ9VrRIAhhPscU2446Aw
dkrpuXFtYOD4HMUg5IpimLwN73nhwvaHVTbrVtSt/OhYReyhjawGdpBcO+tcQnM0eLeCjp2mS8fk
zEZHDuncvzch3VKgrkR+vSTfxMvsTFhvKnta6zbDkmA9Li5HaZspnskQtiLNbMOy9L0BOuG52E+E
sA2RpFOQ3gsQrt0t4ir+OdBxD/hk0AkV9ErhxGthaW0bKtkBe6u7wFw1vttqEUn/VlCvttTAVLCP
w+1HqlXkoy7/HFTprtU+4OrDzvebIyPUh++7Y/DGm+hUd7VOLfiic4uDgaTrZVncoElc2tHgv9c8
Pnv5rhpmXbTwcyo+h27a6ZCe+NRCVscK2MCR/+qGM0bNVyRlhGtRtQ/iQH3KF6da5I8VsBzVnDrS
1nriJm+xrARoTbMU2Ily7rZLK8z35ytcV+XditzJ+LwZesDcyAH46giQxIiET3jiqu74F+igx2Ix
9Z1tycWM41CObd59C+2tS01VuG+4abzVy0WgtCPOnyPW8XoZ2zbcymIGBZxZULquNBGnwcWkrqKo
mww4FnY8UIOXUgMvRW79jcCPTHYYLsszMaIwYR73dnnkmMsf4uPmwZIv1B7Sa7sNRsNSi8/H1sKM
53JMRxlojK/PzwQIUWnh6+Ufs4r0CN1oKhOWQ24f+vsrwTc/RlZFCI/59i16kyT/5E7j5qwtKEmp
0KgfUra0pz2nNA8DUpmecKxFjZuSa2WFX/WzpMGI0PGa4f818375tJH16wXn1DlmoCIcVGPviVD9
LdHqQi66a7ZlMHpFWmjPr7jBAG8jzi7ZXWKaaWMENrTrcAsajuk+TpFTKABU6irsY1D4aunW2SJ6
e8M3LJSmGP5HJXn2CfGqyTgp8QerymkJCaL+8edahYZtoW1IJUW1CojAVipKasYKp+XK4AqdqedR
fmAhdbamzTVUjewVhTyhPagqbRI9E9SDjGnbD/aJCGfx7I5G3Nza3SKOs0j44vDr1k67ajUn4SBi
TbDiMEHF2O4ZUrcRk8YAJ7lQ4BEeCwQ6rvJGLfCXRyXxMCVO9RQnZWvM7rSJl4zXV5iV+d6W9twd
bdQdUDqzQqacjHeBhrN+oY17hpH/w2ucydaLuc49jXaZJ1NMDSRYYTz5r5EZwvwy5axm8mseDgwP
6MtNGGq0hGAM33rztbAyyX52oc0Ie0FoKDOhmQ2fDPjNSlbvx5sJnpSI471doziLZlPcjBNDgJvL
7aSx7yS4XdXgqab3D8xcC2TxbxzLZNeHH+WZ9PwEX6TNTKkqoos7X4cvtGiauA0jpQKF/PK4Lwyk
0ueyMStpPQryOkL2hwDcQZ5ui8QPLJr+PRT5GuwB1f1U6WaSwjWhppZBjw88L67rND0V/KZv+hM5
hGAD4R1kPFpeuSUt+QAsq3yLYh3WtS1rw3arajHF7e0UnCLpN0IdIqA5iL3igxrMQLNwdUmvv6Ja
xczqjeJkxxp/WhL/Qmtahzix7EGLzWeZG/E5iffvoKVcDVa3DHuLpx6bVG9iOG2vksHA81CYAgnW
uS09ivDnm2hVK1qXjCevL7iIcBHBolQ0no5IBiXNr20xUMfymbW1Z95EU0KyIdOTCGeG16J8CQCy
U44VeTLvnrsvk7Xu1hJ2gbZnofAJkH9lwhtM/4xNDdxRwDsMMw5QDZ5CD/fC6d5xya9/kXncVAe6
O7sl1CAoolpY9K4JyOTGheJVPvqg7z+Avwgv0ayMb4zPtrx6GLPFCRooHF3DQ5UovXZZJy/SerA8
StvFkE9ZEjNfC7tr2Fgfr0lIZpUqP6whM9pJKXI05g+OXq6ZC4rxlROC5Q1nEu6tcBrMWG0w3ZRy
7Jop//ip/jaD191+NP43sb0k0uq5TYhPmG1bsrHsU79OB5NRc+1DGvTNykboMX2/3IWHTfTgrRE1
5TDg3QT3iH8aOnr5yB6rfYW255tjwAJIh0eyjLj57aVCGzmcZXn/gTVxd5dMyIIKOMf8vY65P64Z
PDwewzRNMnYAS/wwoZ5o38uq2YJl7cY3uXOGNAkMtb6cQbPV0/wXsHpH2h1SB2UtARYaw76LC7eM
6EWGPv0aCLXB/IY06xIP6X7TFb7G/g9bcWZlxRYAdqLhCDm+ymJj56zFTAFyD2nQB88XCIX1o+CC
WTBHeRgP/fS079XoTFvJtIft8K3H5dT3mEgq+DaDcvHdNpc+IIfWB3faux685u1l+5PSJ9W2fjIG
7umyEIdQBkBchBY6953AR9TKqPfy+q5fc40C46n5Xr96p2kyAwq8akwwxnV9muB/195Wpy3RIhj1
btGeBm0T6V9ijUmo2NDlg8WG80u2WMFLc/oEtBJhz7oJcubsg6blOp0VLBK0gqQjsScI0ngBD8P2
p99L3SxNV04LIlkG/5lL1eWKyUD0kO4dL0M2qA0t2W1gCSbTt46zgYNPMx5prpKQ8o0LtIvNE0jO
pKBKxQj+1MDbl0jzFfG9wBWwsV3mDWO6n1q0g3Vgu0K72kKgD8LtmFiQ3NVRD3zO/CtuKSMInRuP
t1YskVKQhOWpmtHmK7LWaAFMGdwWXKuYedp42fPpMk6Ypw/6lVx3ZeZQkQfvx6oW++mV/gXyy9/O
owMFQeobB5E41HdExonRlylSAbTcMPHfQ/0rmu42dR7wjqVqTeS8bnebfsvh2D+MQq/9oBi/Y3X8
5jgQV1Xnrl/cJjUzLWmvUXne7MTu+NAhcfTrz+z+3eNDEU++4BzwmG8ZXWc1seFyY1UojdqUD0kW
pGA5vJdadkBgId0JhafI6lXHYDyWHGfV28ak23DuZuFi+rNiwJBFVeMaqW4DsoXNFE4YvuM3gCp2
QQWInBWzh4EJZLl4uhEwjHUD2kdfSqgz6KBvhL4dwFVhcVPQqC2eJS1hq0s5yTsg0a6LS+VEfR6S
CwTCLOQqZUdax/J7A1WGmnrAMk7+yHZ8Z5souD1L96s/xYyfmWaQeKW6UTKSdWv23xk/1V2OXL38
RlAPzo4prUsXP2Kl5ZkWMdFEF/R0/P8V1tUDIZ4h7areuVI45wB3XSWO4B1yK0krMH3EU1Tiyk3p
BQphSfXBzk7ASV9GpffRkbeqim3o/llAut0DlSCOn/H2tIXupMyWA3qJiX34sKyRnIvv2NjebyE5
de0Q/cQzHGbLVGcx3exn3ozOJVB7BGb7ZAfp2JL1+QuAZd6JriYBLougqYlGDVWrt354BxPDzqV9
FrO5HDNn9syOFMYp2qx/PwEBd6xSKo8o2KYCK6Gm3EPqiFbv53YIVJ4ikcQyJpZRl2PVawC9uk8I
tGxN5u24uH0CLiMlthglPOLlPzEMHZv4zwqScGA/JcZV7tpLFMEIupzZiH0xrsITZJA71gh45e6w
RUd8BhKrTErtN16MoLW+Tj7yM5jUGmJHErLysCnRNLoawryIuhZJShyoYzngJDVu5hlrgk++dshp
FO56RwfWXvH5m16QthjzItsO9qs1L/QPOkzrtdMSz/1MB/hN/zbbj4iE4PyYazuQ0aBpnvmkvZ4P
lrDj4/PJC406yZwm7U1/486mG9VB5OBkiziYwJaYi1xyLQAmDgD995Jw6m6eh8k2GNMJfIwK5bPt
TivBOeB8/CGkWcK0qoS+tKxH+dPHAkyX9ILNTahIgZT6qJmgrAHzG/QDo211OGCu/VAqajVyIgMk
6Wxw7rXO3F9MYRtyTALynUNMgQfpcw/rSHrOAtJgMZgksjti/HV8+emjXQqzOjCJfi8xDLx8IEtv
SxqoSOnOvwKqr4q4bAaYUUoxp1MM81kte5ocYrAnEO+WV+51FXLpPGHvkP1C3JO7IfQsY+hr/Qsu
LZQsyx9+iztBASc3Qfzz7xjEvk/sOy217+EUgquzGu4NRRp+8xRf5jaDGDeW2nL4jHjyXllHHFn+
+2PysK2UlTOssm2vNayr0oypw0nEIiYHO0baYvAkB3hGeK1CVNnzHHx6Q+/t8MGnuIIH0XBIMPhn
X0+qXyNEHq0vnPlDhF7iX3Wlmj5Uhx0ad3QKt9AmzQTqJgSR57nqdiiseUPI2k8BYAGqFTsv9JTV
sn3kyIzMSVxUWzn6qCys1r2btPJfVNb6ltVBAOaVWpQzW+ZcWNJOqNFM9WluyOfGu5l4eMN5seea
tMVcdihXoU0xMm9yNHLo/M4QYSSR4wTwsAdoKRzZ/wW+XnHDe3zU+u4+OXXKI95pDWH1UC3WeR7e
4QVZjCG3TpYFlsFRT9Y+LUDvydZTrlres+WwQg34sg5X5Fy2cTn+YQKP/MbXjaRmMSnnlOK3b8zM
TZ/BLdMUl7JQXDlTryzntoSUH7NVvFbdsgzAk7yrz7G0H4V1lWdHHB/qIyEMASKdAvyGEpkY2ztd
u0cOkFqTIaJKmNWXKiUD9H2luKYEhQ000YVDIKlHoiwfK0fYDa1URxgmoiIphrMP+Axmb0ee0DDp
oiEp6/RDgd40MuKQMmWba1/lSUSWoJOpltaY0WdNagZd24A9rzhV8Ybwh6TzOsDpgzg2EVOhzWr0
QwFq+baI7DRu3rK4rhVQfjafaBnsdKCj4iJ/vPZq3sTj7wt+hf+id/mGWZS0CXfhPH7q+ldbzJwm
aKfjdoN0AROlJxq8xeRkBVthcgK3h+DITeXSp2YOutr++9Q02s7tUh6AcN1WNPEcN+klB8CMepiU
CS97mirtY7IYiw5Kjoef9idECcpA9IvNdge9fzZI0iwn7hTZQsAFghVxG+SUeYIgh0DCxP16SCQM
KQC02CDZKu88+ZbRZFn40q4b7w/B1fo/2NF/MNGBDsJJvn3blF6Sn1lvpHsOmK2XRCFOjxTQu//J
ce+JXb0vZcHGkvpdh41daTotpo/FxSuKa+OAYHdvhXoVZ6wxbamTwLdscGxfroXnnD2lG0cGjqig
dZEGndfea7ahje5tOHguS2QSRo2eZuvFMm/Iw1TMSHvh8kKEStP9mo6S5T4MrXs+fxhRGLjFJWLI
e6w2eN0nQn+AMhxWbRGGeEk/2JRg5GPlZy7ZibpACPZQNVjrtc9zNKAAM1O2qNi08vNffGp5hwXD
PEhLbv8Za1MtHOFfX5X+f2iHlyWrHUgQ4UIJ/oelayaczPavXafLQQvdPwokk2thsp1fQ8VsnFHH
NMMqkMvEJbH5aL5MGhkGROS1f+XoHpP26LILwI1Mj2ed/+tlo94LbAzRlsjauqeASJOnKzKSwHps
+9A4Xb2AV7I6YbWwS4IzhWxWrGxBWPPqhKk3CiuSjBRZI5/p4N9ua/xQH528xX29p7izyDHjyvA1
lJ5MEtG7U/2/8h+P5AgB2YoRN5zSlZYEwvkSAaBMoqNh9McO/N1I4UIfs53dX8qWMU+xVAudAlO9
0OABTUiZKa2CDqhC9VQ3NxXcGD7Dlvse01v9sDok/uUuMlPsYvGMy40S40eBeEGGj+u0DxUOEpgr
kN6AiN75zcruwyW+zlBSyzEkXLouOv8NeczvQ9j7kMawacWAfzZLb8D2Czn54KFxZZg+RJiE+B5Q
s30nKbopiKhxF+7FYShBK+p9X2aIDtuMBkmnsIdvZdNqHfbgFDVX/9HGToZutqbe9LyOKSCbqxnb
78AxsVEEhGFrUfdJoLCQPZlTSonJ7MD20ls0rf+nUezN3j9fWXslUXCQ/aJDoh9GnhCzrDT1rDxI
bgUbGSRyBcKqET4xwLSRkYUukqZnOvCo5h3wNztriG1HDy472OruEYI4HkJNafXJYmHb9V1rIxr6
WYYTHdl6MDKxQ2eMnLV6Q381B9iLJUWii0qS/29Zz4Zsi7Wb8+PfPpdoft0r4Tm8tHdgxdMudRBJ
uHgIoL2IA/d7m4aCkqrRb3MnGyuA7pNjo+U3lH1bRTDXHgyMXCyBRtIDlLXgwr63yw5fP/pV1ELr
gds4p9aXNPxu+JqiNIM4Px/WPlf5O1cp7wuGECGGjHlU9PxdlgNZMGlaUptoeZPJYwF+PoaLabRZ
lxpg5Uejxo/+Ku25wvNtJgYzoKNl4eDPCfAruqyoWf1KciJBjpuFdNwG3Q8W0znPsse910Tp5iS4
P9wi9Dk4UwOITEmXdj1v2huZrkeeGX2Y0Bly6N8XK7E5BS5K9W0SPDxqwHJyPAJy7wFYwq8Vs5Kr
0F6SF8hyBMWaLzZ2atIsOLYJzYdnkDUudiCmgb/rZcP0IeVodxUxu3eRb6JH3xpeh/vLfayLhViQ
yFUsQbyVcX58bEeXaJdW0llQjccaLgx7dl82O9YetxWsEH6K/qs7vTHRYT3xs4HY88qejM8v10Js
fCkFuEi1dekWOXwDeqCz1FvCNa9RYTJ6v4mkfPk/K+aAgIzfrfL9wrg4tnuWzai95H/ZxtVT63VL
mUQz5jrTZMm774eXsdZbt7rmqukMR7J7KX8hPoq+IiGSGKtJguPlfq0ONbEns2x6jFNBbI4mlyU5
skzZj6Mg+qsiEbFAPNJE5krkSZICFmmM2XJbwpJvkyuxtoo2xFbJZCzuxLuFL4MC7JmOX/soiABC
5xTvlG5KQ+rl5fwxN9ZT/2XzTQKe5g213NoKRjmuDRidbHhq1RgctXia2FvV0Gd9wFh5AHfHLHjj
3AgPq8/Vow1YZwwcwunR+SP3pzFU2sBWZP/1vD58jWmx8i2dryiXDgsDDTJLT2zAo+4h6YlmMfAW
+yIxAE29DjRPWi05JmDIS2M4CtUHI6ZPnaJvNIUKtsCivzYbwkN4L3JcSJzTb0z8bLa8ivRg/kUT
MEdoPM9EwHJP3XV8X7+VARTcjrsS/taV+j325gJqlRHXmUKk+Y6gyQ/JKthad6lJhTjz8osBBqb+
ESDcSo6dRKx+XYXaSyleel6CcaFZq3pcm03n6DEXBhfhBE0jS+YC/acGPBmaCP+A1hgYVfz/AGas
SQL307SdQu9DlJQh/xX+kVZvLSS1MjWbmQ3YBaYkmM7fxVIsf6TSCDv3+fgwd5FWIDKmD0f429YV
isovN8Xs01BpR2B2N+r0CKWfnG5tSf6HAjz0vcyKvRNU36umO6NE9s32q88VwNLfLCRA0Fis7mrN
+vy+dMX0fBkAdu2wSCsFiLofQ3bYcar4KGYVncEDT8RgirdtMf3bKvdPAWUcKaCIyliqyIioLo7F
mGGbdIR0stoBd23yU+NjWXTq268XtLZzV0q2OYlcaXc5jN3kBkCE6sdmfUC2H4h2C1NGvDyEhk7s
rNVCMhU0H+MbNwS9BpYm+vVpkseZGoBakthM8cnmQGv+CNcA8cTPx3ZlkzobVIzPn1X6juEc6GLN
1HjcLBdvzlBApMBvr5/uRNiqdxhcoGx8IDMdoBxxuJaWShdlciAiPFf/Ap0s4KCiKku/YNp5ERPL
DgBNtxsMf3d65uH4eQKYdRR7pjc8TyRJ7cgtsKL7GNkLbArll1fxloftQEQ0NsJ/HcOMFWIPyYle
5bB1EmF8P9fqxNZuIPdPUCiSrXuJ6ZUBejqfPTo4xjnCdLI4NxCa2TjjgpSNk60iYCWBPaoephml
c0Wt2FqfhiHlCHoF8T0TQOpUOnaZZS1eEZ+SejOgzkvWHAwuKFViFL/0IKpECWTavvNjeBHdqFRn
UbN8b6+9DSJ4XYMNln2wWhfVPDq0dZs+FHJmgBSqCTbQZvsC7kKWAyAbr6b2Xi1LO36iVcLKH3ef
Ncub5JMvP6/x01tcBe8x6ROihsSt3q4zv9IpmcGH0m5KsAvls+I2d3KQc9qfBG000CTODPqKkYo0
EuN68O7ajv9vk3cdn1EUhanPa0v4NVaq8tcYle/FzWgObyScSGX6rNHwwbwa94OxDu2qU+fVnoHB
emy0dG8CvN4jeMliKqAM+y0L30XAd+/7fHb4OCiYPedLGDqEZ3KIKHylACz0XvIf8qaofnNpLXRh
ViKMG5/Eelguq6bQDze0RkfAVyOdAWOCoiHaAMcDb3dEYU8bGeXY9VtboW47L3SyC0qJoo5fBgdx
wYvI/4iOfg0HUQ73zjxl7S49MlVfPNsGzhw9KA5LjEQIq5clz4dHxabYNVUXLqnNQVfWekQIINej
PsbMvIO9ig1wLIBVCIe7C3zqyGjzv2KU54wBD9h1rOxTbcm6Jyyebo5g4uAfGw1T9MlJqmrXEL5C
dn5GgUBYaJxuwTqLsEWWOANOKUOGTw6A+juEldFjikJB2ZCKTHIu7uMEvKyyvRiiMHbSKbhGci6t
Qrspm7m/oIAQEAwMHgVqLcUxETtCragBzTEJormydTewqGWBf/auiBrAFwK39gT/jM02w0cFtiba
XmORJOYxbBNOzJDeLw2J55JiPSUgnLWCFhbusFKmNc40HNPl1FtfpJcspjjC3mu6/FW3W0oPeVqc
TyKZI5yeDYTPfJeJ/P+c2g52Az427JiFnakdnsY9pX/fyBQPP8Wi2ocP5kGnsQJA4tZddpIQk1ZU
e+e/bWZGdf00/6oHjr00wenl+wLe+5SB0Rx3VwVMD8p7hPnidhNZ6YsMhSLQI+hpQHAYjdwSloaI
r1Pdt9JMJqXSO8LW1T7+EF7w34R3OkkStejAs8VlEzBtJk1f+ciWcESAnq36lyjdD2nA5/OtbjUz
F3BrScvjoTdBW08+PVJLlCWVdDm+due4bnGeruTuMmjOg8UysAGJJU6TL6F2cJ2RTX6ATacZqS47
iqn0DWBn5On3QFkI0qjlSC1oUkQ3z/61PYTHFuDRn1g/OHp/5DS4Ml7I5abfql5m49syIl3SZDV0
46CJlp0mi5Dou637tmgykNbtnGIp8dsunieinHAQyv3Mgy1PoSRb9GJxrdvY+XiuPuHtb+YxZkDF
nlBJzpQdLEzb8sbLglHFuRuQLMmEXJVH4ITCO2hjDM7lrAFiVqtpojqDSloKrFnfACIz7a0Jw/7m
SlfYLARTcF2JtGl1n3g2hS57mAsO9jhWknvTnUvBZPyQdF2VYdaIsnJYBA0Wm6pwk1HYQQOlCvtp
rXl1GVnIKaEqO0SlWV6dIEk2dk+v09FSrsxtJxeH/scFCX/Gr43DgwZJbAk9zncPpVkOLFywVUE1
hJCVcuOHjGDTslsB6GHsQbMaK4QaOSymWO2QrdDPWIJL3OcNh4HnAFK38qLgrZBsQuf2F5a1sbPp
RYNgdxKphi/w6ty8FBXAkYfLHLeOK7rBQTYiYD14GaE+fhiwz49KBGc6IesTO2nTh5Uv7uymf3e2
sZi/qo9SHTy0qr4Wjb+dblTRHqspfZigoePEFwjpVwlGIvzBm1qLwDQuNv+snUDjolh47wjPNUkJ
eTH7/F3s5RI9/AjUZCFBDzvFm1SjW/dwtsam3gBsGbPb8mKQp6KC7i5SuuhJx+LGGgNmRBlwCwdC
gklig8c5TEkLxqRE/9j/VPm0seibRX65+9+GHRyF8WJxXk9vw8AU40XphAy71q5cIQTYnkjlGko2
CtFkU/DmaZzl78utXeS02EwG34jzX5RHqRtnt61e7WGoQ3sLV3E2j6zkO9KvL10PuwH/59A297tV
fDwNSZDZbtFTSRsKq+spn8QhGKDUxlNleylVXWdrEbuHBTMbP87wew0ggRVWsLVPRu7W/cgVG3S8
C5IFx1//0xHcX7DLuOkKlv+Kz2hGzbgVtPgLq71P4L0gZWvTpqbOp2sWXQW+LCsq30Wok4ZZcoOG
VQWrTrBJb2mPB2+StvhyVVVDgTAiQUT6G1XsyTq2xNGkQ2mBGHS1dVNrDAQOJTOGPyl/RxVx6d9T
aqEtv0/BssNQlt79haiOG2BXM+kXnwX2clgXNFO24U1ZN82ooFI6pbejn4e1HEXLHIty2hl8T67B
vZ1rdG9vdcbtClbv47zhjFJx4J6t+ng0N03KSxOT5JSnFlc6DyKEpbFRnBXeR5+iFOEvMIOSHG8b
DhM3DsNDVnj9QPjTrAfCEGodhNvi5DEzH0Wzx+5XspQYxmmDfsGOQcdSLjO/Cb4+lSIkvZhW0J3+
k/oHtDMD6UxKvp3WI/ZYZtrzQ4t06qK1tXy9U2dNL6NxISqCMbc+JTIE60ZuINwal0hAgKva/CAT
cfOQ0qqZEN+I79AcZ4y0+f33VhpEtwALyQQdzjJU43QZ0iXLsJ0VrCuVrpxMNZMYhUI2nLiEiQfp
VsGpHZaXGWz8aKSU24L9rmmtWlXJSnOvXv9ho5QIRKHXqwKXG98KdftnBpq433QnmLfr5lzoMF45
pqHAe/pe8ovYAkHgr+E8GVJmIKDu6iUyicLs9bbh0v5N8JO/teBRr26KeRm9rpGU1yJdmafUmxDT
5HbKJim7c868fQzolBnKHQyze7hc1CqCB2xKESFEoeSnqIs0i9k1YxJd8v7fywRYlvOptp3G5b5u
0PLg6dkAFLq4N9ogMiBA3/1v2aKY61JFMawmXcm92kDVkVxiykRCo+lCBUxT1uyNoDpj2F9t6GGt
S+1OxE39gPoAk2JPVxI5EwtSzeJKbL1+4poORXRF0J/1Lgk31VZ/55FrF0nr2zE4ZE7pLanR8WY5
uhCSzMU2dOxgDnbSMlbyFi0ARKakztT5eocWGVOY9C6RGLZLmR2vyWgmuWCN3R6laAPT5IC6mbzl
qVU1EQIOJweqfVjlvLZvXYiOeAr8PBVRmcvNPYHig38db3OwIqS+G1hi/aQiM6mgW5N3302NgR5i
QNq9H6f9fUXZb/7+AhIVxnaN2DLr/CGNSsB3d49bU7pf9A8Zh8eaSbOzKuN1Exh7LChpOaOvc0g5
Iupm//3XLbouzgPsJPNF4am9L3qPwFRXzX1gVwdLaLqWaFsoM3ZNkwxI9oprk7mSzAmHXyNgeceg
9Izpn+UIdY+FiyBUeezUYBxHDq736h/PoDmlyyTjvUxcNNUfRxhMllW/IUXMkbTBCnsXu0TFiJ19
wKKSb48stMm32z0nOIwyMFAMI2667fJOW3TgiEWqUTTZeU+7UYdPGYw1wogmvVZ7h8/1cjhe5qkZ
O/f1iIf0/JODUoNws0LlIHGNYoDgJaxuRBvz54MzU4NxIKQN4cwtg2JE7fStTOoS1Asw5M/A6f70
OgZlb7CEOHo8ZGySJm9z564yitpR+IkQbMnJs3aVaRRrusItYJhnfeQ57cp5vv+RLFB5dgUs6cPw
DshB77yKmsRqyrVkKiHvHN9JLWHicZhOcKD6sJ29H4sOfO81F12YomucnofpL5iQv4bpt7LI81Mw
BT4lzHK4ufUGF0Nh6CK4gcQmAbKYVJoRr7AjsvchwtoZyrOdIVrVR0RIRi7RVcCONYE2P9ZpH3Dn
GaQ2kixazY5WCzMRiy99Ai8BeD4Cx8TbGCsKALKaogpuATHSGUW8C5VifEl3OeyrKM3vZk+apm5u
j5mZddmObyATdbmbL2TjrAAmOY7xFASKmaBJETjgDpGxNf57K1YrnFq5w9dQOz44ii5Tai0qhvuB
XquheSjW5teB8FwoKKTMaBdhJWV+faFqJ6+E4qr0R7m9kDYip+7ZqQLZzCQAFp8XtQip2ry5Hek+
PdctmQDX8eCM9BAUFBMtFkGO1QpHZU68z5+ZpS4CLivlGxcVrp+8Y9U+icSe4hLpdVqjL8iJxguE
Fzp23f36I41FXGc2ZMNlomR3eUUs6VQsXmrnUSlxlxBk2bQFLslaPT7nkRfSq3Vm0OyzC7zsa1bS
Dik8S9uwe6D4/DqKXg5VIayzTTJs5jDdwP/6ojCJ8B3wjTC0xcclndMlMWfWRIIOzXz9H+RvYpUc
1czicKeJqOsTuJuEd1csmyEl4LbHLB8Rbumw768lnrJFNGoBR47WREg2N2ET95jBGmxXMvr69xOm
84cCH7H3e5vGPRUpRaL5oRAVXIzEt9sY3u1J0wgntfo5GQybKLpBls/ppEQKWUSrYpZ8grKcqopQ
TwCDboB0Gsep3Icyd01kKUH62b0RJqeLrBKyupxSEtLK0rqO2lDnbrY7iIKNZRL5m2ubsoUFrWKj
N4QkGdOXiGMN6T2gyQAYCzV0eFl0I6T6BiMSHsE4Ekx9351Xkz1TFu2gJZ7tTnwzDEdURF72Ih6f
WeREjGVRPq/WuRAnpc6vXx2ggcaV7o1nSFsv5UmoNRVM6ZhyI0Ns3jrnAZrhu3RX9qTHx1Sgo293
bqK9g2l1YrY8KH/bkUoCVLuSzzjwnvpsK2lEYfjlOOvpv33PO7fN9n2nUhW/8l38jhCSjUJvbVHG
nKnhp25XCNsX3/e0BYeoPSuWMlnPK0g8dDTHwq81h8Y5/rSMj1iVwdaexMOeksNxricEsykVD3MZ
NM7OXyYJ2BUFvFXjpCDJM6BoGasJMvFkQBK7VPyPzM/Pub3awqOMWXhm10fHbemQFmYoPnzfWZAd
YiiIOthgORItP2cBHWTPjANP9BMhSUkIfGXfsNrZ9FRUzhAGFMkDQkw5UhUp1CFiDhldSOSFpvrN
v8rH6SNecXJMn0zhVCH4Nc5/l6rCrTUD5wB1FOrm3dbYPugTzJz45niN632Cv82ZlYzE5oMwVn7Q
UZ6uj0827E31VxoSXRvBNaKzM3khgovBe38LsQVGKSIIrVfHa1ivFAoUaFkmeQ6fO/a5HdPUzrcm
mFNiVJx0eIzgqUVlrzRCZ9SmQL0lfyJ7sB2P2dAkqcSbIIx+mKw3AkF6HUAHvlwJPZClWuuCP0Tm
xX7P6L1NuhLX0U6qwqva+MqBrawgGQ7C/oj8bMSYN95Bg4fjCn2jHmwKZnRSRN3pt1e6gxJnssRM
kk4QDFhWAtBrkdUCeH26zy/LVCmgcKN3dbZ4LdA9xoyWNYBFCF02W3t06uweTeYa73ltfqm8tuBV
RoiYmhwjoxK985OfDud05PvGBp/6Otqy3TTKh/VGigiGp0HySOgPvq2AFQDn1oJB7npQz5hZwUKI
xt92sHyuHzLubvONECrg9NGtUh7GSzpdb443YDlEPkMLijHNPjq/YEmg3PT9WGddm0yzezGnjqRB
tEhQNOk+dz8bdpPXyj3bnL+NBbHxlBUMDjn/9uQ90KZhcb94P3khQZ5Ovc6ytMt/fSMdy7Qgq0r0
cE7SwDWXu1V249KSRyO4ju7mc7A/iT2g8yO56y67TUtgaMGX8SiZp++Kh6LYj02p+N71CBPWcl49
ZC2/RJTmC5kBmwCoXQO14GbucUkGqmo7ofi4845TSjMlfA/sMia54PWQ9XooneZoaMvdy5DGOKwU
Dws42yQ+xR6x+fCxEgYz54eOI1vvriq47BPi+dvQGKlOWKQMyoZ+K6GHjr9U0eQ4KpmRNX9lyXqP
Lh6tr+PYlECkHt+Mb95/Qw+fw2G0OcIRyncYnSY5JVc1WR5PzloZw5ZE1T2jE2t8SJnZIY54DmDG
zW78mp0vl0pRWlDyvn5tRmwLZWFMlo9wyjFMaz51rmEr0SAl9f/gunV8CXixFtgbPpZMP+DC9AmF
FTqxqeuT1Hw3AzMVem2SPyJe0zPcadnsUhJ7VGu6qA4U701VfvYLiY0fR+T6YVmZUfcJLUuR7BgH
DZdlSVubnpP9I6pCWe41FzvFmNdqhrsvgwt55sOf+wWMvIYHzFjkURa2BTtRL+9G5xGYjKKyAnQm
8Sb+fX/0wVSiITxgyuqHvB3sDGQNWk+h8DDTy8DuCqyvk5lHDETT6z3GOAffBst0AlV5uKaUM5IU
qwCx97L9mFSREFM84R2NJOu1s9hWN38X9zbuLPkYdDwIf4QVDZ2ohrsoml8GhBVQDFJJVNrFL4sD
WuYyk9HIOD0KLH+XXi2xH8QsAKIODhfVLO/65bNvFeKARV9J+qXr3NwbO/WhKRZ8kPwd6t7nAMAV
1r1ZTG+VBmUPFCKxYg5B7rMCjbxTCFiaPS7803r5v/JSRECmyRYF9pLZJ8E0PxWcFoi2E3vz+ZNU
TqgP6SnI+QLenIB4uXb5fDIgDrMIuYtykdfOudG1yrdhmQy4psRgSVrnWzr32227eax2vx2KrxeG
UGis5yTUooAfUSdcCZHpp8YBEmt87erlZZrB1sJIW8kuf6ivHnZ5htsRuKJexDY0ge4GDHHDTjdm
OMnyNryWdWtQRDGUeMFvMjx6nEDj30NM/s5lqexrdLdDEk81qtLJ+gCd0p3KfmFdzb/dU77bgypi
JTt3KtEQ1TcKy9lvMcH9lmZZFujKB+a6stH/E3PGsTwjQ/fSjqvo7ScypV88V93u0kk2tRGloH6t
ijdZ/LEtuHvNcT6xuJbA3WGzeYWjWl1cpr3Dt4yta5Kcxrs7vdJ0CdPYQq61fIaUQMBhOKUjpBWH
XndTTMI0aSIm85TtyAFqzo5WBXv8GYSvQrNofsSDAyxVkOM2Z0M65DE/7VD5ugTVgla0zFmUJciS
uvuOwSgq6HaAUq7V/zdfgF7nxTZCKDMu48aGNsoi504kIjIaK1VINKlJxXqQYAhStHdAiUCTiOr9
HGsPK2ky8o43CqCFDkQhSc0qE1ZbYL0st+aK0tt3mhHSVyQI43/C5Wwzaw8ETz0zchG571rO00db
mJ+LJddLIQ/kPRe2FEGTgcPLcgvWr8dwb2y5Abr2+133LbkLvoeovBp/9pL4vJaRGxtgiA5+yJJs
L7j21VhdJho2Mmpgm5/o3BOpvJOmr6o7wkalJUyA6uTQwnUcW8VqViK4wX+cnw52dy05LoWJcMBS
Vs5zO8mJ/7beRBCceui6+7hEyUmAABG6nCXJKFktSzZrRq8IUPlkEFyqSMXXL4eJlHU8weBqX2tp
FZYFG3SgC074wxzZVJYClWGXLJj4pngE1avyRGiAvFfpxNAqRcGiLj3WeGBCEZMOyuHQjuBKPikD
gGW3nm7DNJ54n5Gs8kAuvSCl5gala7VSmb1msBAdWQRnrcIdlQfJvuJyPRkpEYPe+h8igct7QA4M
dVXJYejLOOWfOEcUXb7imEAP8/hsRdv8kzrtLHCC0ArBRkamQ6zR2xosoYTbBDTCX516UphnZZ4c
RrzIzxOmc16JPPuAPzf4FA6jcECzuCbaUpRuBjRw6O7M4M0K9HuJU3XAfXEyZ9JdUYX56CnwBplT
J4/hLg7liStTHm6A8xCtr7TgS+yXBUJbWsc6O+GcayOwF01WMvqtEnUypTvUG/1NstSi449U6wDT
13UY9HFMUxCo046uaBl/8eT5iGTIKfyA6ZM7ScPViVtpn6fbqeEMfRD5lJjDT6i26MlyIt+0fS7S
jPrZkYRmWHlWOnSW8J73nm2cqTfd2kh0K5jp/FSjOi/hmTuCySH23B3AawnTe+6/hApvfYm2113d
f2RLyCJT+JLfkrzJ/WBAJ3xclHsPVLLyjNTscY/F1l4HA83sD61chd2h3ANUraeWgKQlfNQQRiHh
BjgK3kyk5hIWK8fBhc+/e5HTI+hLLRabI1v0nETC0hKAM+FUlsQvAS7w/aUZumIsuuLr6foK6Hdt
cNCVRzGODZsn/GJqKZP9130BwP7+hQocujlJvujf12063SGvJq+lahs86ubxM7/6r0+XdYqN58jw
cEVwTlqUgGIWc8+Uj1BWGs8yiLxfz+0qNsT7iXc7HffzX/0hMPVCrbhGFx58Jj6zAXgiPjcw7dmW
BQwpynM/snIbj1tJUREtOaB/ftcI5cpOXBtWMVyKEJHwcjy84BpK0NX+khfY4HJIRfajKM3tLhai
fNC324R9IOnx75Q1n7IVlgRtWx0ZjAnBuw2PgoBnJ2HKXMuirztCFipbpk+WBHmVrySncJzI4MZ2
spNKM7w0MAGJVPQcvajJswuyzSzjUScYuW/xebw3/BIbRWMg0UawSSxHAJbf3JC7CU+NmSXYC4IU
4VisZ+8sQgKU7BKUQ7uHx6vqJ4z43LqfHoMTDrbO8PbomUjopScu+m7Qmbd4zVISnHeHDUMldwZq
MPjYFjVm+DLu6UuJYnBZqOvHRqsxdU+dVW4s2tjATj9sLPrQLAUQd3A8Badq1Epg/a9dJKhyh0RB
iqhpz78eP4p5fTcLbZyzhMUpT6x3IXV2TKT1GYqoneM6kG//7MnuNIS3NbsCNsjhZkHj9xQmzdem
mdx7D46/zUsXFxDox/SjEUvrF5mgz7K7Sa0MOZv2OinDTs+aOrMYmexLA+TZXCr9ZV6Ry+tz/8xz
fCNQapl8hPhRHP5nQqIYaOFkOI2Cymh9zTWr8NJ1mV798YjOfjySnfsvgaZj2PcU9aMu/3/sFrpz
RIrT73Q0vbR/IwCC+gV4isNiDA4DwNhDMqiPMYXFB0tenu4TdpNWF+4/4J0HGZDivgPAkQ2fjh1u
8bJipWo3vUJ01SvaWySzie/+6dMJAfDeqU6F6cDRGEbSD4Xz/rIY1O+xgfgXuZeH3yg42sKTSd7k
pyStMHqXDf9jr+A5zaURcwS2q+71JM4twZOcFN/jT+laElLGoi1Eam5JySTtn7I3dn1CNYN0yadQ
dFROV4hM0Z+pmIWh7pqaoPcutesj91FeMMlRSIlHmV4BTxb5cdfsQopFslKp6ol2hQAZNjYlYHNS
R+iKinzHzYpHyVgTbdNS5zMab3LeO/XP54dG8sZGbPffybxPwpYAhzrMSf1+ketxi7bQYbMnksnl
DbpXH3nWHFCw1/PHqz9Z7IC3kjqNAe7hVADqgTfTTxM6QUl8p/dr6e6K01VkVJBq1TAuBnsmRRnn
szRV3uBQIFBC1ZN88txg2aMQTHF4VBn2BWLzvlLqdh++4hLUrGM+KC4G8dgoM+KsDRcD6RO3Gpfi
yBznVqOL3QRCxqEumYk+rrUnZd99hoZTH85r9KClo7qAZSOKeS/meF1gpGni+WWZ2zaO+BMlw+4V
LFPTxlQTlpzTT0h7T/VgkJ4QtNPYv32giLnIhJGdfYaRA0jeHCqnCGM/SCRB2GcOl2aKC2xbKt4I
IgZ1xP9YjIl2AigvipR+XMsqKWYJZdJCN/57mOt+VppfaV5cBfYtz8hNSCPPf9Eg5Xz7B09U05sg
+tQv+ssao/qmssb44KIoyejTWAM2ybfeHnVcTnPEvd2rNxnlcCmRQ0PlpUSz4CHO48KLLu+ETlQ0
k5KNw4KCBzMqc6udGrv4MRtRNVOpP/IC+7xcZF3RXRKZ9I4XldPwUjb5wiiPMSMZo6/IWlBGwX2j
1TzQZQfasWMZnkToqg8nzltegj5Rl2oQtKSH/i2A/O3a6+NvskAn2sJpBOQmwsS9P5POLT601BJ7
li2o54P6DTk3Lgf1aPKBQ3aYykWahRSfBG+2EAsr2BaR818To9mj2Y1eXHAnVUpDYlKDrR9vO1WB
JLmouRdJxIY3aaDZZedsqQaFBu/g29B8qa14j2TgHspr3DQNNv1FSmjNsjRvT4vsPL3vLEeSnORC
VT6LCRCheaUcyrE8TCZf/AaainzuRKbx5UDOuqRqkEScvyupQuwEMD1bFWVNrRthMufCKscJu6FA
Y22uvoywXi9VZvTfle7ogTd+YCdns7aPSp955YTR5aTydSWyLZd8X13kKU31h8yA9e6GnWPBwpdu
Tzkka30vdW8tUxzlnjrEy9OhOAyYlOaKI3fYLQgnZwWgV3eZhVxYjXhTThc+WqCetmy/AKoZmAD1
3Y1R4WpMdV7kQOde7DhYZg44RhP9mSaRetvAvRAIbVqncVFva6wR7lve6f6nqN4W9e8j+1S8k2Kj
haXpE66Eu9rEWehJcgYsTNprJV54MW9Qt8C+0ltVCs550tnfsQB//dqklkB7kTE1+1aVyl/M+PW1
HN29bMhmFhisysz2rjJxf8kwJG/caUptniDXuYy8rK7TN29wuBmpaHSV7TknQuE6azVbdIAKQcHW
U8xB5ApDT+NoROv+J75BduLixRpjCiPXHGMxCV5Tf2ZC20nbq4NXZkSG9CJDVadoq/zFZhU8bdqS
IGqdqy0vCu+ekLvvxjf1uc2cMZOShfXOGSqktp4dwFqRZEUvulRSDwlMpQZ8ToOQzPRntRIO1/SL
DCRbPiIElIfScDgNjVxwAtq71nWWNxMf0UMG2N5o9Qp42RoGwn+t/q1BJimhOwMwTGxTQnK0hdwK
OuMwJQ+GLfMkqcV+d9m7uVzpyRCiEaIv4rdWHO9Q7ptmLAvqd+zT22GBn1Ahzv3LGzac0rGpeMCs
izGW32Mfye93B3NsqeYIcPh4tUceA7GVrygDsOPQn28tpLV9hsHEEUO2GL/7thtPHnil9b6Mv4C6
2YfJy5UzVPuvxOgW+Csc+IVmzcjRh5MFL50d1gQ4WHbuyYuf0Yz2s4a0rWwW3J1Jr92XOlHRGCqX
l5Y8EF/oLGR8YGOTS4jjzLBxoR372yrpb6JQ1Bbqp6EClaYyY6Vpia8XXNzG8aU5f0gM2EhPAz1W
QFrVlfv1G08PMLrfAlsFQLQz/vnGoiZr0w+9nyIxz9eFztOlSoHVkC8Tn2ylnQR5A7BGKoKj0FuZ
VR5APiFwfaJxBwMXG6D09no1+LDWlHvfo7FGHiJmUQtI+zPEBjXNu4H2Cf/7P2p6gp+QmimOn6mV
tS57/ekKcBWt9hlCuNF/hqWrGwx5LiNbleNYFESBUSlU3dpDVRE4pTKiIyGpqqJJ58L4WDNcGyaC
INRMLxqs+Rp75GKzJ37S+d5yPlbeaPhMOSEwFRAqjdOAmJL5LNtZohhICvX47i74wifQZdunG29e
0n/CM6zeihyHeZTC94tqmUVwMNjS7QZkh7HNA5/+IhrdwEjzUzVjjqJcUR0X8esArJu3Kih5he7H
vr/134rgHRkx0W/MpkkrJppgisT56ctQYvRUJTWcDUF7xxBxTMJ2LZRt6XevgSHX/vRABkvM4z1q
LuKqykarjUWbREPaNaU76XA8D0jKevYgRqhDRJxe/7Lm7BRruK86IsqicftuEDImHdbQ46ubS0Or
Bl9dNxwTUUI6oyn3u/VFPmN3UmsX4JIos9W/lzuiyVPwFVgPEQNyXGAxcaYbGx1okoK2Gk4U9ivV
ED8C6r/he8OCkbdlqxExtmskDRDtxSTJKBzFQoJvdtZQx++chqWciMdRphF3g2hpAxKrEex/EMTn
plIzVZb9l6s8XwTz7hVBggI3L/bggVH3+aWxsFslppq8qZYaUpc2UV8640yy8uh6FPiNZiyJmDDm
t5e4NCC28KxKqm7mdKjo6dLcB5O5wdGX7X/ye6xGn+K6vkcUaALM7NoKPI3tDvTFKexP6yR7pOrV
QXBjbiDbKSv/Q7YXb/IWn6cpqjapvZgmC/jxhc+jyUd17GjMQUshwneuDpmYUYTE3qmwZQN6PAaI
8LR2KvskohFyMRWEQa6z45kZ+LHrJs80jTGUXRPJzp+DyCUSau3z+A2UeXsf8RYfAzf0BfiDlF8k
lx+xc8LNsUzNnZdj8hpGnn0XjwP4Ok0kFIBLmzlDkMOu60RTsRT/BS/IRf/99/LvZc+/ySJJ2/sG
a7C492VZmlyXOIKBMdVrqYPmC/cfIHNRiZJtztC4DC/XWbNXOD2uusMbw1ai9iiXmxFzcLq6QUA+
hP27Va2u/mC+R0yPEpjKyHMwM4gwrBxhfiP85BWqoevULDEjGCqGiysiMVGO9R4xSFRPmSSIA0vs
WZDml5eDZeTpgDoJwZixtdDV9UFGRsD5v+Gk5gc286uJ2fx0lV+YxYRKgT8irgh/EQjo0OUhJM3/
Rf+NENZSVzGfkvdXrxJyeo8u2mc+7W6XQd/ft+2YqAMMihBkNrjjGgN2y2Qstlq1FrAwkZQq3kLe
6dv1Yi/G059o1LonOaUAfAK33K+gzoLMI2dsezUlvf1AcxXsHEH7tTO9pVQUEOVlvRZC5MboUMs/
gyKfmr6q6t3Suy6sUorSwh2WNIPSJt/6ZjQ7zRucoU/gL5P3+nXee3toTbu83HQegV4O59IBunhj
opr8M0lvot6eE6ocG/4kv9ziqrpQadosV9yGNdQvFrS/5Yz7ir/Ld1LaBj54UeJqHDcYVuQft3hc
DGEjkzYRKTwhKgXIDGAccXkKS4uT075ORjPjK9s5QRajte6Hx5we6QhUids069ShGOCi1mr9bVUj
v9WZwGuMLwg92HwztHydz0lA8t8rhBmk2gj2mM31GviqolOiBrcjLVhdAivQe1YZPKLDK6kcgO+M
dh6Z989aLtY511zY0YkzGt3dUCxCyzZusAlysiljUxBgDYYAdFnUBF/Kq+Mod9Yii5DzFC9Wzhmp
8ty1n/yz8y4zOYOktl0NW6tWD5jUHC3GyJWl0IoSRCPVcXUxoqG7DMEemAjHPRtN+wdCaaFHdcIG
XcW23ijKDSZu0nzJjvNRMhYTlA9io9eE08cvWj4JT3LmShX9xQew948luJbf0hKhCLvnRqkymGeQ
qJetSL6dsocCWckIKsqs4cH1wuFDPRve8Ca9y0hKmMhumvQ6GvIOmLkn4CWNYJhLeZYUx/o+PfWm
bshMlN91o43x2H3ClgaHsNEVcHaxrmAAv+zZqXzpgk+RETqzBQD+yWOOQYd/TwLU0j+E/Ojb/MWE
JYOhxaLAWZm6HNfGQW2Nb5YhnIrKgPqc+XgkI6GqCeWl2yhfmjujWy6g+8c+sWKnVZU8urN/lHgP
WrSy6wImuI6DLSv680Wv7VxzfW15O+bAU0eUEL79VO9TwXLAUoUI4MgbBQsgJUECjiqMN3iD5Nmu
DL5G6lIsNKbPEWBHs2YyLx1unZBsam+fT7AmXhFTAAZwj2mlCo7+AFDy5YDyQ2ntY9qpBl5doxHi
UUze45Z2Z4t2k/8X4zDsIzhHnnGFIvXfLWqCOi+LkfCP7kL22A6Osb6BfMPuWdzzfjT3MsJSctBy
p4WgBKw8IA9ZaAERslsM8YKPcrP6f3DdQy3iJdO8EncpE57nS4updN+6W6RJdJTYJvmELH78bMxm
9jvZXBt2eu5ycPLMfdMwlJ1KCn+P2e5U4wOha7L0jtnWP2XXSmO8IidX8K90GbzOTN2IOSsbagsH
ONZZIkx5sGWCDIM3zLdCNnGd5m/cnLowiF8aMMjy6tvsrrnYEPMTr4DuXWbIFeoII53i3VWHLmxQ
v8WjCFtNO5BxUJ6t2+9KDQbq1X3Rh8F4zFjyKUuF8TNrgYZ78hiEuOyRssdAS6yaIrM4o6Z1/DVd
+MZXgTJBLdc23j0PvShEUv5ydUm0QggWWHfV93wev/z9g3BdNeSlAnzQAJdyXWdW90iZRWRzVMnM
o5xrtuRfm/MGQzEGh3bHRvXIzxBDvWic1LzDSJn9ZxVtsVXb4cX1QEIkfcxst4PCfYgJEEP5D9wU
8IahVgxecsh/eZFBC+bvzUmKW5Fp3fXtTzZg6Q29FgPwSuUjpaDF7ruwvLSD+BVPjRjCnuBaPgcr
qO5LsOPN+S0XjWrNSlvbKlt4HfCSfmhqBKcCgUtwAnozYGwztkPQAwn6l+VuB5P5plOykOvzr0+y
8nGp8UvQNplxvQqountlIWVjFnGEpM079/i2xXX5xIACwtpVEHBBhgZpvnG8G2vmvcLYaivZ5uCU
Nd2YdT9aKfjBNtrQSpDkmLC7il8ILpymRYgvZFGfiLAAxP8jezI0n0oQNmXeOJFibTHVGlcUX4YA
SCX0a7LzKRRxziKswfq/jJ1jYqNI9rn5dJw4VJjG7/AA7X3F26uaCFfGTQf3T9F2HhotKKX7uga4
E0ieQ2Af3zaK3El963JKBxdL6kOnhCuuZ3XoStiyBlFjCKnvbfd9CUdXvsQ9tCDzvXX6TQ9WTH6u
FjuEl95ScQk8Trphh+RHu441dhfdXqE3PuNnbbMmJkMcikii+qdLNSDzXKQp2YhBxR74QS5BjmUR
aEYKY5rqGXhOEyjQOUBLP57Io6dBeujy3AiEY8n4aj9KtVmhWooKn0W9OsjKfxB8pxFb9tAc1jkg
A78dc7vDneefhMVtXCGPG/fVxVu0nFj4/wup/1XUdG0ZKZdNkA8x6sJ5uBC9PeVKwu+EY7Mg/CwP
KP3AMnzRCDfldWCDCbBBcaj85vWP2lyiYTHdKVamqDxd9/DddI/VmHvFfyk6orq6w1ohT/E3katb
/+fHp8JMeQuI6HUEIdU95gIO6y0LADqw7YahfH4nQ3/eYdnCGlqPzpmx/v+cmz5x9jKBK5NoOSP/
z8YG9Tzm0XxFb+xK6owb+AXQsHSOq9h8WTqjI2WvpTiTKPu7HXnEn45X979V2FZf5Ef0+9bmM+C0
erQF9tj0IMOC7VCdHqR18NeL+w1zE5zMAFRldQSWL7aAunkwCxl7nCHI/1koPavVQF8GGk0/V8bP
pxb+WOOsb12r1b5lA72sBTOBKLrQEIzdqzIrtWSGUXzPyJML4Acu6wKZTjq4kQUS4ZOWYWZL7ugZ
So90aAtpFATnCnjsOsy+JPTJLT+SDiwnYjni9U5XbIQLMLu6LWYEtMjn/UBVHRO+v/muvmjMAdoC
XH73KgnRuusMBoNLDApspuKwckfPRKgWalrRXsv5CV+TTFcr07hE8JKNnti+vPXoTPzd+yP2iCJT
QYA2R4ejSGV8c3ntsMmnZPMn7XxRRGWuTfrtt7trIhv4mpWIztyt1YUiYbCsHj1r3KkoHho95Dwy
KjxrTuTmpFoFUfg+pDVicamIdL+rA2WtwNQE3nuowDdlS3sF+cWqe1MEy6geX6DauGja0kI4rWR0
llh13EVJmBL3eZs/DeNhKczYLci05bd5tfuEuuJsNY1DDmkoZ09gpmBDBw8uEC1KT2pReK96y2Rj
T3YTWLxhvk7d4OxEqC5TKmWUPvT7KaIgeOR1AVyDznjZc4zJ1nZOuIC4rZ+EwsMK1+RLMCwXwpMS
elAIc8dOYpanep8lWDUrJZrvbqWAVeGH3OypoepVp2tAgTT37p1HVxnlOMj8yanU8V5i7xenaVwT
gV1vUbJy5pj+SGGP946y7kGWjnOYNpws+UoJ/uIXK3a50unlgx12QNzIkAkqqrnZSz0Vx6A5Dvn+
haJuoBZ/mRoGOZPsO7eBW9gT4FqMU0Q/GIC2CKO71X8jeOz6z3Bq5HATwtI4XqVnkJIgOVUZAEz+
TDpNHQnv551NxdVVgBPCcVyMFYhSnQVX7bNPOtrUNWJVXGwNc6kIE754isYmrErSl7VIIAlgYoDG
fHm5irfJEhbN040EKO4TIIsaE7ehp8vX2fg1KlBQW+6sh+g4PLzfktRWuJ3J0GKseyMYS/KFrabc
fWnWAsBwZZUsNaIk/umMwe/mXNwmd3hVrGTAFLMgH4sfK9VAvU/PLZrODyAq1zga5aABcQl7R8Ya
HEYVeUVx2LhcQGMppcEq+P6sVAAyX/e3QKgeBXk4Kv81KzcF8XbCC+MveJdyAPsPsEX8jWhnG8JB
8iRZqIK18aHAG9I6SvDiiCtSYtCK2rordYCZ04CAdKhG1m5+puL8QkJTc7XTuMDdhfw1sCPmErIY
lQGEheFzI0BhnYmT8UTvsLjk6iyJjdeVKtD1ESe+5wrfjRHq9Z54596eX9cQv110mlbxThhwmMHF
t+AvMksc9rO4PytNZ5TTmA67DNZeRpDTg01WYX7tzXbPzugtx2i8gKXoNsO3FzSxRr+pL9ODZjGl
1YaY2jl9P4mS/DZDYZzwikBahqSubtzP9nXEXh05D49LlcaaU4IMl9ZmBG6xxnn6jWQ+lR9bHSFd
uQdePX4ORJgYqZlrarhPbxO3JkjiDo0x+fHVMjm4ibl3/ocPZiD1hqm2lDGsXd+Ee7iy6bZI4tHz
40N95L+bgFnfUBXi0UtmYZtuuy9B9fLvMBzH5Tpgs6xJ38uXuLWbSSiE6wvmL+xSnuSnYvFU74f0
TNlh5qWum+6MMSatKRQslBV7YWaqBTvBxXrO2YKAdYs9+sDB6q7+6E14yNyYcQBEFa3So0lewFQH
omL3ee4zA5iDztUL1yAVHZyg/mWEJ5VYGnOiqdzj7LDZXuWNj/9b4kgxebKYGNEq56rMO87UWsth
/T81OFHyjpTmZThu/Q0ZiWMD4VkCQ32OTy3CCFNANbxpv7ak6kD4/eW5IeiZyyzjImJd+79/P8T4
FWhCUlTTEZKr5OrY3AWJPKK70bK+CE3q8/uXvckm1ytDhDEbIR9ysui/7vLkwHhH43AyYh1uccoa
rJkoa10IgZGAdNTEvytGi8LOe2MW1kXaxYh6YlLZKnBH8E70Bkf08IDxHp8t6YFxVgVxmyfJuEp4
ALWF5sEwP70K97+eMcyl1XgayuaieN5TMNYsB21aMxzCI+vcLvFmfysGQ89tnpJYu9E8LzWRIqwg
u4eO3ByjQPA7J0hF/ZMEzwGIX57XrmE4HH54Bqyb2i6heetAnT3nhEyEoOR7qf5SlJZ52yPGdNWH
S1P5F5d++5MwMtoewcZHKJu8BiBWpNz/tEvFQxCyUN3WjNOeBbChFN8L+jh/qxlch0Vvw+K2RiLu
SsQGkZCPRKU7SfIJofD67/FDvWlhKLsoOoBXNQgDncd48TC6Frx9NaI27p3P0vSP+KBfOwMzoiHF
uv3SYCFfq9bHTez/qX1pantCvFFY+iUB5JK+Xk+ew0y92jwtqnc/dmoolNL8N+h7is57nagm3MNW
FApaZMppr+swwKRRX8dnx0TaXfOsADQdGWPdLDg5mjO5gDQ9TLCxcLEwtfX92ayXTE7kZLynBCHV
OQqG6l+hDxbgosmcegQs9LS43J198g5CkWwVx4TQpk0rHrUPk4HF/LoG1LJSxY/jWzcV2Bmg7fci
VNmCauHE84nPiz1O60t4U942IZxKoErnscJhCfK+32kYDbXO1zwm5j4ct8sIBaMH6eYgrYQLivPU
mM6gxd4W8rAsMbF3fx7oHkE0jmJVF0u+7NG2jNPO7w6EGvIlBeh/B9Oh+589VypRiHXmPj/Lo9UL
p4eg6g9UlRYdvokwhxlCAFP3EnIhMLPFfEiq+5AklyThpdF6ETmUlKMH2gBsDO9IDBpViCMp2hDg
eJLh1VMXi4h+6qn8te07FwZtoDCN6sTXcxDK6qvFvtbiKcd5eeNVSw1GE2udihsm6kC/yqAK28H2
PY7nHt3UiXlzg8lo+207Jfn2TIlDHZ034rE9n6aGTqWNxlv14iKWpTQh51nfcaIq/MvKc/xtvG36
Zo9UEGzYVWiR01bn9kmxkkJNeA1XdEBonbnamPsyzGPs14hf5KsyQstw0WND9l5eEhk4j74xLQaH
8uW4tfwuifyODqq9QprGrIZHq8TI/FuR5y3CTvmsRmtoR0Jo3E7onV9CYQ2blBUHIHq6CftJdXd1
Hd+gMQOeQd+d8qk64OFPMSGo2gqI/uqwSNcZQL7sQRgivQR+b76/t48UqrWBaMC737gBrLJikfxQ
J6mzH/INZdcLGGCI4pBwAdiFdAkX8GSdRJMOh30UzIlcKYwgdMj7Fwiqy5RS7cf5/WH4TzrUt97q
HrZMAo+MVjKSOXnNGCjPth2bBwl1vctLkOXCwUoUPt2U3hPjhh1DBfy7ygUJh6S/06F+rVGsZEnc
ED5x+JBuO29sbZotXUXO7dIPZkOz++IoGlQ2oL8I9WHezUBgjXOGDJn3BcFAFqkF4GsZIBnRV4wd
TtiyEHVl8v2Bce7U4h1Wr70OZP+IWwD5QQ0OOG1/e4C1zvX1ZTI5OczAlc+ECIFrs840Elq+dPeE
BmOi0kQ7USGnyzltORV6snu6v7Fdw9/8rR4d8sE2UoLDSS/TLC/3gT8oh4wa3yWfydJEx90a+eZQ
qyfEs+Q7M8oBStaQrowgAHvc8mvtcranLuCwI5+oB8fejhMvOLIHFpGhfG4A6y7cfodYAfoMFsVh
LHtyu2ymZJsYsQ2GWF8kPzVla+BemNmoPGy2/pPowVEPteOUflYM7rpCcpdcapMNpPLLcc1CX8mv
WOTaPh+TWwzWoMmc2aapgy/LZcJmpjImFDBTVohRvFIRTls9rQv5HOb67ttts6YDTkkNN5eAyT0X
0KIjhc2cv2TCvnXZ309LT+RH4KWbzZHUksJSMotda/V21IubSGlV1gb9ZRD3eGCM6g/ilsEz6hf+
eouPDlzwpAlGCuaE8ZXcT/e2EkoGfc9mK/cU3n3E0lFC3HZuahw8I7Ev/cxn5hRbsQtv8QId9dmW
/GbZsO0LliWcHpmNyCSxFJ/er/IWEyhxi8jsAJsAwaKpIjlLdLvVK6wkoKj4LSUgX8vas8yaut8U
gxod9dmahXjS6Dwrd+vxLRBcTomBvKu78iIglT8hd+F8gmSiaxIV01UvLFeucslUkpqSGaHWrI5K
uK0bmCB9Ygviak0AFajW+XzVPHdmxKFVkvjhBliBNTETMnQRxuHQUDf7UBftW7K2SVRswF3C5Yf5
5444pKQm8Vkmg50+d8hfKk0T5uSb0cvweF5g6Lys6LFzfaUwdomJ8Neett3DaVNWwN66lvzYucf+
ZrSZD2vAVB8482lVrlC0SLYTafQZ961TBy/rY6gtnxtnR5ij7OjVBAfRraWH3Nm4xK+2HJfYbKDA
Rp47JWkYznXpg39BtT5/xovpLWzHSI1rG6/0XP8e750wh/h2nlGC35+cjVjMU39kg4WOKDk/ESL2
wdh6Fk3Wub6bgaUl1OkV58/vGkzNK5UV6mF0AoY1ZtMuUJGltbt2ZbRri6nMEDhTrBPfew68XLwq
otkeSTBpyGkgvr8l3VvDnavt4MCn/BE2bAlzuiJZB5MQr3GNUU4RUcjvO7whxVmiTcsYSLM6h35c
sXmfxvCONk2NCvDs7gqPy6AttTQCzpcNNhxZ4Yu9WbFUOQEpxdoA91xaVUUPyXUBPoMGwXNtiCx3
2q+SfL5Uq1lSmTT9w6tpBeBtChUeG/ZiSmL4OI2/yEGITJqlgvZXdLtu7b/baZMTCPhjVXc5lNT3
3z2cnGEgKIXu911yu8IclmtCc3DqiVzx9dAC7ygPN3Y34jpyoRGFfDhaT+hlxhKMGb2lVtq61jZm
wqqcPMY+Nb6n0jzI0pYgFJP+nozT4IaFutDgpdXbR4u4OBzMw/NdkL0YwQjl2xbLFae5pwYstWby
cRDNjAbulC6tIraXUwv4cCf8BpxNfIAotX7cNZBJhnyZFnhK5IXjIqbCdeH1JjEi0SXaHQP+emim
SffALV/GYlLv1bA6HU9GG3LGge3iwZ9Hs/FbdqiwoRBgNK2lMQwXxIbrhEVXI4yqaSanKzgpVxcK
GZJA9WGIysPafBtC3usF9/Cmu1WMh84dvgzXOEt/ylQXvVfErMFHATKFJCjdzxmgRhe4Qykt+QBP
Y+vST5fhF7wrz89ycvHLYVpwaOmTBL5Fm+F0euYl2wOg5t4DP8cth0GBNVW5eAComrmnPlGHCA5L
DJAHcgPYi8sZ1hpkq9XLG5SZ4A7SFBEHdBDZaMITMyr1BI+JjbaO6E/72/A6CXn3AihQQoaLx4tg
rTXJ62ej/8x7K8Hsv4eOqDjhnGpRQZzdaNQhYvN291AoptXuiUI1KJwhGUtEHvuCk/y11cgdNPEl
t8JtEDKYUDXlcCXQzCUwdnZaNdqBEbtfTm9vvEEoy+5mt/08tLVTSk91kO3A6hj5eXUqnmDoH4in
PRTC/AcevmtoCt4nxVonRntWs3+KO7GsoiOB1Zmf4Uq3rKwzrVB65R9h+ChAkCVR+10WkAsGMuPu
1vmxUPqkDdMZCAM+xbwf/f5xBZkQUwAEwv2u9BfMJFbTc7BP49dZYrASLI2ytvcnENYsvPghb9QQ
0cqk9scf5yaOK4QNJf6+4dA+cSS9/YlRT6C9D+Y7K/xHv49rFZKfz0iascZ+bZIaCgJtYebHQgvE
W7d+Vc6XezSNYkr7QJdUSsF0UXUXT5R603Y1Zys56dlT1afYhwzruWz5YAXQcHfRHwOiX4gYW49w
9hgm30r7o09F3FlXYgD4ZD9asRUON8rl48429kRG07QD1P+nPupXPxH8KMKhD7UDx44g4gURXI99
CaQPiaos4XwC1eFB9c26IJ03kOoqiJHvXgUYzHGt5GPAsj1azR54abDFoBGiJ5vsdSdh7uLyCfFt
g1Rh2pBg648opMhJaJ3mXxWxvCqotR1IpdrvzQxaTrNNsH8ca6DserDDGg9l32eDAjGAKzYKCwso
KiuG+rO1lNNJOg8dEqoAEZCjtuiDnL6qW3n5Lzy7lOk0L5krNHF8XTcdmdlLe8WHGF3yzIqiun+p
9d3CvhJwX2i66Hhu2+D+6eJhlxfA/eRoVmg3Y0LjiJZbl6PQq9DuNwCzsrDrBy0tbB7JzB31K1Wg
VVNES1CogTvJ+7ljy+ypga83XsVadsjeiQRWjO/5KT5fDJxbTa6YP8HpGv4gq3VM09WrdIi8EUXs
QJfJdUAt+Oj9ecMxoLbt0co1zf2PSMrtBY8Ra7uO14Gy/qAF/EmBHk6XS6NXXuJZwvzeJNRzqjZw
eWvvyyNwRpnveCdy7psS4sWrVz1cu2xxg6OnOLA7kChkKEyWl8g3pbhRbXklb1pE26a5D1CLxrTY
qhiMjI8yJPTUjJYwAVR2HEVrkjUJPZMCvTt2kOGHZtMSEtI7WYK2s+UeocNSC7bJa0HKx7oUJNGt
iP1Ug/v5mZLS0Ykf0BgJaH4Gre0+MV4+tdCidXtgflYv4vNLO6NgCnBSQLk1haNCwdP6RiSziKDw
50VOHg2W/JVNR99yD868XQzCofIGquNglIsUuFiAIGZXEDqHf2iY5QaFeIN1AIG3aVLUR7Bk6v3s
IStA/JRMF9XF2yr4tZt04AeL7gW2XIIGLp5uuoTH04nUjHnknuldk7L3IIl6I7KEFN0EahJLsX2B
k46jnFl8S3jZcqJgIQmRDJxJXFLmb1mUXlumpC2w4MYLtBeN5Db2LDhbCYuR4M4kcPZuDWcFF0RQ
wNf83h4J4ZPlIWkocTx5NrY9f4xLtv6K+3L8UfUpp9VOSNwhHs4TNPkJqOs/pNAYWZh7IO6JFaGn
TwhaRfu4vSXjpzPZhiMN/3W+x/XP9XhP+gOOVormctWLSDOUYTBe8IPVfIv6wPcb3OxOSzd9VvSs
Yx8cxv98IqqNUfoHBU3AWpltk0a72mUcnu3IU19aDeY+lD4597yoCkhYewgTEmXj/ZVPGj6jTbvX
ZIfLgWM11ZTOoQ5V7SiIqFOLVNZjVtt/xe0PfwNuH+9RDlvVv1EptVDf2AbeVHoQC1QvZVNCILHo
olWN9KHr8jmSKTYdKG40GNnZ16g32HG+HzXIXMXBmL/p0tdAtKOFjlNfDH3XBIp6Pygn74prYCJV
qi2by6ti2EyQs/jtse4lVZMWWIVVpNxwJilT9QX9iv3EbkTuO5l2vMFo663aPa3DwlUzn9zRi4eJ
5bNKJpS+z/W99oVx7OwrjX58YFlaYHxCD10LQ6ZQIhqsYfDnsLu699k6I3AiDXdNmHhaAjnPQg0d
5t0p6HfJyZax/Iz/xXBlbhNylMAOSxhWhkl3CQbZoNskCOiQSHNuLhNJ200iQJY3dlVcT8955jNX
oaaWTIAlZqvJYCHAsP4TzB/72jyAXd3nhciU0a9h+Tf4w6n9Ge64PYx6IDdBUu6qGrzQ4np429hh
IoBX27E4zKDk/eL0+/p6z96kK6JuXCVIQIjfke+dufi4oXXZn2KhW7gavGCZDJEx3g8ywVcnHjH0
D5mZETOWJi8ybDfdKIUvXg0R6W+O1jRxeAX2NIxQKWvvD6Kd8KuBlir36ou/IxqQYE8Sw+HssTMf
7piQjP67uDpPDBc+W+miS559HuYhzZqeJajN4EU+Gjpy4OerXllp3CHA8zu6ZktJYfzKt+v0pCjd
ZG34w/3qjjxtyu49yg2W8SQxhyqDJhzzvSoQD/kFpqAMKHSVZaO54bi//9nZ6XhA0T4TRJ2OtCyL
KYADNt4O7Wv31EIqrgd/J+QocEADjTIK9B9qxwFJsK7JRXX0yCVjmVqRYXjYDP+RpGBLOKxJAhIn
spNxpiCQnKyELax+z+wz4q+Hhv2aVRrum6sUk6Lu/jV+ZgsqkBRpMwwha/RWl2MQ+nd1YPnlTOzm
4leiliogLCQEWsqYmFBMWcSypzkBs5BtUmMYZ47ved9jviruT8jcuw1LuESaQM0EJNHxXeeNWbTT
tnVdIxtOhSkpYG2GCCj1B/TCbAvlTer+dCYoCabR2Vflm0SBuYP8FMwpBp7M7A0FG2akaYCtFCWK
75DtRXfctK1a4UmHv41Prviwn4mQ9VC0KA9IgKLQgSRkiz7NmOblKAxZEIYu+t/cfFOMGRK7NgZy
NFglFF0FAB6P3fcUW4+I1eorykcTkV19Hoh1l6o5tbHrcFOvA9quxy2tyZD9sOs3Pt6bu4sPn5Oq
Yma/xucjPeDfihreW1bzU3QqVmBRTIA5HE4LneOACLRbr0422jWwuAK0ZRJR67eIVeGeSu+PnCZX
Uz53O+lYvtCwcJMx8GqBGnMV2VfVjmkmRVuhT+y8TaJYJqgzQ4I/ngbLZm88Ej5yaqCzbKn0CAJK
GjPRczXxpTkt1Fvs4G6yIwc6z1yw1aIiw1ofAsVrGk+dqzxohWCzQ5ITCWpdKfnyqsNNqEE/wEaw
LJFolNbTiMaRFx23MJlSBWZC8RLKwes4yZvTz3MZyn681Yuxud+H9+7WKrKv4/084Vk3tF3H6BN0
bQ5DA5u3kFXq/tGAe0XHJpSjVxuh6wBUQyfvthJYTNuKRHWBrAe3NnQ/bJcwr6OPSI2zsk8peDAM
zXMJkLV3dAG7KXAPRcLdshTUUAvej5cH5RvNRCAAGlk72f7V2BfQmiO3K2O3qARiQW4Ir0PPRBWn
/Wdb1djwy2jMV79ssP/lldx51CiGmfJE4ER0/13x66DJlX/aad5sYt8pG+tLEtQwTtUHwl2aJhbZ
QOEjlHFYrDlkZWlR8B3CY2QT2X8+f9DbIivK3WTB4+TCJH7pK0F1FLpI526a1bu90sEYXA0ngai5
t+G7Bg74scVeoFy+6vW0/REAWkdHYA/3uiXSlMyQUpCIYSMwgVODU30KU1f3tyC5iQ2QnKyXSLaR
RmHEk6NvoMigk3Q8tf9YbRKMQM8xiDoDnc31csaPSIWWnRZwiqa762Ma78q/XFWrnu+24z0Ven6Z
W7XWWbEOD5KX/sBpLN9cW0LSOISvry9qH2AVWhllj7LHMmKc98/1dQNJIxotyvPim+05VnWtDJur
d9ZOWrgP7ZBUzglN5Q3KPMvjtfeqIMajq9K7YnbYdMEudbbEUDEh0/i0ng47clpSmlQd6nRw5btH
ki5kaZ8DLfyLJjgy2bjxVh3Djv15Rp47W6WEaiFc20HjzYuVuH3LN/xhX2vXkcVOL/dFdXM8thaZ
PZFs5pma3YhyNkgWwhAxzh5UTZnVytU0Tzjkicy+CA7F6w92sMcIoZmdUcyZnvOAAq2jJX4UleIa
Zn1KnWDUBXRqAqil0pcqSNS6Y3M1pnTVe62y/Q743hwGqvd1smOPmySNdhNpz8PgkqfeSZvNsG+A
4Uz01he3/OHLI9Rtrths1DdzNlNfRe8cowZQ7BdyjFAVGvKMB9kj1PhTqq5dRxugnBDpPczhA8nL
anqkjYdcOY+kvKwfPlIgZO5BTt3UqVjt4OGlKGeMQTMm3pRE5w6jDoxLlJN8i6nWztPbgPcMeiQ8
AWqt8i2BQqRmaejHQaxfhJinE2nHXshCHy5GVHzgLwNmlsFbtF7llFLCybrDjHAYaCkYQ0K45KAw
n/mgBkkZgzIuFIO+AVH3HU1LYG62HFv+zaFUZYE3uL0zAVINTZ/M81Hvvte3JCto3Wu5UWLkLxUq
vtr1hPOyUpSRigry8bWwVJ+pyQyoV1b6F53XF7crzy2c2+/5CtLjxmt5dDuSLVqC6r1kAzB4EgUn
S73Bq02bM+D7wIrRw8GMI368hN4yxKf7CRFdhGMewK1NGX9TC00zZlga3p6WLB0CIbysqyPHiip3
/6lna+NTD8X5jEdHCcuYoLAhpRQJXD9A8tzQoRkNTeZanMtu0Wu/MFbUhUYHxJnQ0eim3fd89H42
0SQOlmWY1pdhBQEfcyb8hXRqLYf6X9GyHEoXRaIFF9rwR14CiEFTVQDuVaveSbXTdaxELDUqo3tK
mmUo+Ik4o+atBNk5Rycf0Ns1HqkoBUlUJdlKKf86jlQb0vHRjWYuXIcoleF4kd+ZVNbKGFDhr90v
dleJ/Cbj/d9QPmRWtd/kA36SWK1nBIPPjfpot5ksXH569pqtw09yEhG1xpUOL28AZAjCSDFLLmA6
FJ3aEEWSnxQiAdu/w5Lv8aQrfZgyzaKsDviXXy54gChs0M1c7JIiWgUoXijfZ2GKnxkVnYZ2JmNT
fvTYubSho+QlMNNPi4teQ8E4y8R87dVWCkz6Hqv4rbKw9eX+7Ykt2zI5L8w8YXfWqG4B8xr6+d40
MxTADlypD6ApPRdt/JLmA0LoGFVVoQ5oq46ZaY61NELm1R7JpJ4TbcqT2Fpx7/cpv9EKvQDsI0Xr
25L1NM4uABQT3+vqV9U+iK/4xFmlY4CulniG0wdHkxRWOhzj6fTYg4RUJppfSkKkqeAPyA0fIxcb
+TyTTstdyMAOvc+ADihdoxPl2GbfmMmnBdASGIYUVgJQGnxKt2v/B3Wu1B73xAriI/BSYn2rLXiZ
T32SeCphPAeq4AhvFMwXzaM8Lr2nc4c2Q7xj8xmpY1Tm/36TOS0cfvnPKrT/LuISi6xFJMDm+flh
GBHHM+CCwvddb4rP31qvPEsPMcRpJnwDYol8ccwlM+lfT4t340611404jkA1XRsOBW6Rz7oNu9df
iUpD9RLnFRIN5tjzoY6iB1vHsT0jC8w4aVDudpH+UxB4yfYnh5wlyNhlPPoCU9PeV08EQDjCZ1Oq
EJVoDk2YxqDosxHkrX4yZ07+PGgAtvapItUA1qcQ+w7tpJzSaA5ptwkiolfLKmIKjroXXKFhIStn
NV6lFSUd7YwRhTAxEd8McsXLoOYvkWyAZz8dkxM60wW3oAGQUidO5cxnVxQhckPGJJiFB1QPlyRF
c4ByPy6BzXlfiUbtFgSzIpCfiw73k5s6y6Iklvo5mjqIfubihaWmxVvsmvU2DfgOKrzX+AcO9g2e
fVEtPnGrrhGb1hCbxq4ccOogHbIlp8sHLJyaCQ0Uvt483aHkqSv6YpbT7UkzaYoOugKy+py6GCW4
b7sJ8ZE6s5nJEn174se+4sA8o/+U3LfRQRceFWC0V9rGWMAf4UHj3vr+6JKX/pcTBZWXWc/1QkY3
BeliOGt7PqMfbTwKGublQSxv9wTHPCNHd7QKsk4w1tMPQkvyQ+7umm0xvVwKJ1IADak+9iH079f8
UvG/bYASRB4xPexlmm1cWl/kJvTfwOSrGL5MdVJRqNWkTFYrs9lskTmlk4slKWG60m65Hd5gQ/pD
mHpkshM0XaJgAMZJJv7WLZXt8vRGf6T1zpaiFrCAeOUcgQY7v8rxNnRzroTAekC1fgOvUU/DnoBD
vdhJffqi/Ny1+vcXf8t6KXrK53VcHufmPdU5A73i9l2Fb2JGawfeYoLFCTRqQkMiZFIGNnCgQBkv
zx6wCg0hExNz0oko4ieFhpIegBO0ptRpI47LKMTLXckDIpWCm5E8j1GOW8P6sZNmCGpG3f17AX7B
jZU4j4SQxI70sweq6J14KBTr0bhSBCF8R9mzFcjFjfUZg4Ct/j212sElvtAUptlpDnAVpCgoAlEs
uCUyLoa5P7KSb+lt2I9Sgjz1m2b+h+Y/GGZdATX30pk1tb7aJgpH/1Bv1iBFA+HdqzC0NYhIDjph
WmH240VzgutZWxpP05juj8K0b/4DO29iA/gkIpVu59/ZgKO90ERr9iFR0h2rxHn9BMUtK0PR1oJ7
Rma9g0ZQFoh/XfqBsxuqcFOS3XVpfAnm0kOXbUBkdfHc4V7q61Gjo66+dyhQ50Dvuq9hVBf5JbuU
6HAnzt/StJo2RzH6Y8sziueDtiFZKSw9RhqvI9hzXRwDYZNZ15EJUeuRT1V9As3VzGD46Q5xFGwU
RxpDdIxRQDQHZeq/4kzRAVQrvltYOSw4TcncKMVO3bcClmVVXmq/Lkbg4YTHwO/03baNmldl3vAp
q1m3OVhXZ5/y0NqXYzZBpRl9v2O1EbAxbw+ltvwD5elpQ6as04nDyUeo/8jYYsp1sP/+uD8JLNne
vnzc7vtYjn7uv1sENyfhfK83mC4CXqkdoezhHQFVleF5ndDVsoXQ0WI5ItNINb3SsorvvAb01W3Y
EHEbwHmMdT1/hBAFKgjJMVjRx+VpNUGsIkxxuuFxQGVO68uBogdmkYiMsfGOw6t4U9JubKqK8CqL
fRsZEEZ7o9W2pHneyDiO6+0ocP/yDAo79JEfuY+omr3AeOvyU8nydondLXn2ZGJCfdW7F9wrIa04
YX+jF9/tgl0ON9oB05QpR+BURgYsn8e8oEI/aV//eoQNR8f7eR4KBnQ+tUO+mkXRVX1zqKGi8gc0
BsfjGdWefj80LMxydMYSHNjK9uR/V7gfV6F0jORnRKW0gx+JAFbHAWAQhcWoe8STVRwBLSV6g2A2
hmfD77AvOnA6IUNoTuPBREpZDAf3BMgPfkSMB3axljS4hp1jPg+TUY8qrBsDKYzUMeRIoe57gj5y
az6bfVExV5ZNi3wbL/2LFm+AMLe0znrNlMt4EpENI12mzu1utmydEYNnVkmBi3Pv4dMBTDsSQB+f
AwFV0VLWXkRS5geWLpb3/DgaxHkCftRkdiYiS3Q1ZBnriV5OWoTluxM3bMnLmCV4Q1AdKf2VEDlp
cg7RA2B85vebLt9LuTWeyYCpbaDQsKrWOFxn4SvGDsC+ZBeALb7qpykGFBoSVx2MEHuuJD4EgcLU
tlQWFEOL9mYkALUgFk9bQ6vHA0ylhnPZfVOjjHjJRYsqOtp/DmEAA5+okLDbfg3ru2qxB2BaX92V
zooJASK/wwdCNu3rqxDybqsJxgqkcjqsqaLKiDD+UPnAZjPkgPlGl9WxiONqnWRgHsHDRilYp1fa
d0T0oe/m+kAkwQxyrzwh2gy7lRnd28d/ahoIyiqaxB069C/5SwUeosBfKuonlk80K1gUdLYGQlp5
n0ycnkafDVmChUHNtGFNtCCPaLCHw9k3LcSScdQiEf2Khua/40YNnWfXkX0Q1PQPNMCRz/EfnIwl
jzI0LCYHDiOBZi+YxzQjZYwEHJ4nLDMKjDoWf1WW7nXr3jizSy565HXA901wtNdJd0GkvxLRSpxh
UFmoM9zubvVWmHaeJyryFJFZKbzMAUYK5hpZBjUp0hyVyFNUXuurL6fhx8SkkfSfA18y/V40e3a+
WtxmHgW8X/8zy1SkJRur0iOL/0w3r9eCHckzztA/TbzQExuwc4JUoSw3XVGF1w8Wf+fp2CnQRGDL
Y4xnIo5LNES5MXUBiFO+Hgx5hu6JRmnni+vADZlju1vlmoP/YwVXIZXKmyxP9VE5HZDzEqu2VyL5
x/Hzdd8V1hrL1yuM/1hcDomqZyYtoZ0cM6UHrdxIkYbfW2Rm8NWzz7dVfTS3JVOQMpi5OhcR1cIr
PStic/Mx4kaIyBf5KQUOirxa+c0ok36Qc2BjDXFhiO5AvSECinJPTeTWJhcLkrWpn17Zf2t7O1sZ
M+n2JxruuqmQpw1leQTTxWc2zwxXnFG6FcLjqNXPtct6+3vTuD5fnAxidbYlEymboX00fIMtmhAf
CvhKI3/8NOuqo0zMACbe8UY2kWKpgvfRN2jdZBm1pIYwoen9D1MqrLLkOyw7ZVBrF917K25UhZuQ
4GAnST1Et8NvYGkVa+zTSi3p3H5RWeFPz6HuhbtHX1nLsYedPW6Ol88ZS1lnVwShuiUYPa45NQlK
tBWaDv9tQc/keIJC2gQTXcXpiVnGYrPDksCpZAT7cjHcNiWO1iHLivLZ3PlbRuYwS0pHsM4Fv18L
1Mq/kbWQuJX+cIx1mdyZ+aVOdywkv6lQNhor6XgbccHZHwiJPCDc2jZk3QWsH/pSlFeQMdvXQdSq
APAXy8S6l1j+J73qGpwBfm0yiTeaopebg9wuW0NfgxptdfTTysv7ajRk2mc4PfvY+LJLP8HzPwTN
lvuXq/rCFrrd8KplQ6MBgVGQ4kfWqT4F4GCb/q3Ype1eY0uIUh0fDPyz1+o/khCCzttgZiK4e465
mUI5jtKkGFCQy8dzGNaG2quRPkWPwTGHO3BYGZo7XYg/CQUAuwKTMRkCO70Js48fql43sx30Ax67
lxW0TRtnQsWRaKNtok/RX3l5yQBG/OJJkZQOcx65a7Q76zlPPRyjqmJzTz6z78imSQPaJUS+Va56
S051Qi2vXQzWGnhUCkg3QKusRD2rL14yRkN91t9b+9Zqc4sTGRYsTSJCTKCFl58A2h+7xxwxpil9
NIJj6kqFk0hLWzp7ARKUa0YCm9P5v+X8AJ9cOKYJDXTpM5OZXnfrVzYY/rzchemOMuezRFns+A5i
bpJkpEO/HhUwJ3iY8+KbjEu7n3+3avyR1EcFe62A47Gv/5XIdBrmziP86ja/+B2hFI1sfTqE/aGs
UGg7jSL/UmKeM21iy1H5eRfL4DaiIddUC2IPvDMScHIq5LGe5H93VGUvq2QwtGbnqGT4rLmQFSsF
xP9bF1u8gD7rcaPZzBG5e40vbMvMUCh6jnnSg60LxJKH9F2YEFZWp1924uEjfJiiRqz/hTz40q+y
xZ6rMD9VfTZTF1EXio7FaGwcjMdFn3sDAQtC3YiDKRmjzdo0GxExhiS4f/cSLXk32p8icBNczW7c
nlyhkJSHXXdxM6J/ArjmdYTty+2KdbNG6pWwE1anHdmtySTyWxBuKIz5/t1u19MZriDI4xAE9xtF
rBHmacYQA6n1Br0Hgi1yjrEy6wp00YG5IN0i5xG48MjkAdmmg1bR33SloieIYAnDQ5cwqWY5bDMp
Fm1iz5Vle2YxZmWPc40Hm2vEozG6v6e/6/sZHc+Psksvx20zGoCH4E6cdOXTg38NnCWyJH6MRTDm
1BJapnQ/onWfN1TiyYtJ6Y1OtD2O6UP8g+6go9QwYRgYKQjKPLsVi/V9FN1LJ24Eso9RnoKgQCCK
sAydl1kMcQ/6lh8rEbhBkP+7TWFvvDRcX1cMOGbo5jW8w/aWWKoz1vTKuVHpB6crPCnvgFuStE/+
I+5ANh/yNFixViBtmcxojzQx2MtVz+JRtCtcohhCutA97XJdgGtmA/qDAt0zQHCGSH2Bw2SMVbUX
AAj0bCCx7khNJ0rLSFdAOexoT7AHzM0NBxmJHVHs+mwePGPdH+YWk7Eeswp9Vd9mdgJJ70JnVgp9
kHSoNK6ROdKvKGQOw2N/kYUnFTlxGlys4puzwMaqLR4WExUoslqizJUw0qL3cTHYoFz8uQJQguhf
chYVimbJRr0U1lhJG7EE8l1S+N5Ab/UjNXRXjE8tl79Tj0BOfuxBl+CsHPE6SSdnsxEmmQXC50AN
usxXCylX/4y987TRM5Vat5oquqPr8HCWcnxgNsiKaih6Uvqd3B5w1gAtmbhJMxZvlc3adZFHBjLZ
XVNjk5Rp0wboXlcIBvWjytSK2wXR28J/oPclMYVbKpHgEA3RlfwyWNXbzWWIfv5j7bCaCaaPprlK
BQxPKBmR2J9cmP2HBs+4X8eVhIgACPF9OjNzxAz+lpVKgayR0C+7anyKXzU5c6yU4RieWd/JbmIl
FZRgAieFTr0jW2Xs+qgsvh4T6hTWwxDHTv4rcc5W8Jzcun0xf+OAxhCl3Wps6gn5NYb2gMghDt1L
dvLpqvppc2vgOTEEczv/ChPJ7AtK1edIuiWjQzSG9/xgjGslhv65LpznrU/5/pi5uUbosn03/QaO
lCkIvr5x7sAMHyWzfFF+MzwczZMCvCwRvclpW8xXtw5khuXgVkQx+mLUsNy2s3VUToU+4dkoeeMs
jhqv4LsShB126a7aATxr9YW0Mut/HLuYEgB4bvghFOV+BQcn3ebmCKYrJXbDs/ak1eOOmqvG1In5
cEvlhzKvFahWhqK/VeyWbL1OhivgM0qJI/M0xqQ/MdfzTNgjnqPCFyDoMoXslEGR4zuePi/7dYoB
xFwQFz5Rumm1T2j0ssb5vGfIAOGpOkVwERKPNAhn51vnO093+Ac0InTpbOZTc2dhWXRdCa2dkdmo
qtjhT26uQeHeB9m+tQ/o0KtBrVhvhWLaEd+dt818XwWaIEMiK1CtHpMnhug5YfxnUsgpaNuOWWxo
/+Tcny3hmFHMvLo1ierYicOHnmmP1BESpPfP0JibYfZxcenxuRORwckI47hJOqhzI0x0fQn+wk2H
mta2CrvGaQGGnkMhfFttz2hKuo+fkoEVh5/8u3RZBEPgF9pONYCXG+nBbvTgQqVoGCyI4jaC4Zej
ctGkKKk/WOaLXi/J1rLF9WBq+ovr+e34uF3gSs2A7expQ3gLujKuuAsTEnw9aVElQ84zw0MWMiBX
wt8kNuq4VQK873UpOHhdzFelh2joEPHwHCtX14fYqt08B0Qpbi90EiPURYS9d8aDOq+GW1YP2N5I
K9akau3LPrmOXTkOxQLIBgOF6wMbwMOn3K9qduDvSXAp84mrUaxJedD+896Ab4IsDTj6vD4WtGAp
phTYYCvv289bVtOY3v5SP8reOc8hoItgPwVHWBkyDqVfZlS13TFh33pOsiOC31ZGyiuBgO2/G50w
MrPluaIK6mtE3KdKYWPf/KuhXNzHj9LT0zUAIqI8Fm5h8cnTBxBLVbbTUQgZCXIPf07mS8nWq3FX
vMQFTS0NDW1uImiPP8uM2ZdzZ/cqXv6yC8oFvEiAAyDrIQ4GWWuDN51g9pGTuUTh7/jmA+AJH3hG
7MkbQvz/ZAa4AMj/aQI0GqFoO5789J5rzwGpWQXKSwVlq0wEnJH2FR+dkeCG+HWvSl7AN/DhRGIa
r8slpK1MlUuivM+W7RkITgCAu7AFpbjWHr8KGaHgXrNWKbQ3q74DcSO7MfoEAKaa1c93Vk9VZK84
DAfkcOLxNGxpADg0Y5SdB0zT47w1sDCV4Vr+5POGju0fia3ZnG+X+p16dh3AiQcGIm3ewWEtl/KD
AeutA/J9MTRyr1XXH5zLs78k2FfR/KdUtHYtfYRwOZKm0yQjpw8CqJk0PwmALi/VlUYGje1d5LVp
WAU+yDz0oy1zX7Cj7jUXLNuckhf9DZfUwYiRq2M9BIbPA3pJSf9J5tkADUZ5KoLzCFFY+M0bSq0d
ZidS7FNUShbnCpMLIzAHLJeTumFNHVlAx8IW6ZQe2Kg6mA1JWqa3HNc+FsDI5cgSk3Fhq+t+lF5v
UajTtL4G1/nLwX3ELkZkXrtmCcRAGgdpB1ASsrgdPl6SVxt3V2xFQV8lDI+7i1XnUFSYVmTIosCL
A4RLSQAhe1tROxEiRjNo0LqDQQ1w1xuVoaNXUirfJX7F0uiqkEsNuNQI/P2VjbJGdQYulDUiZpE8
6lEi3nunhthOfyEFLcV4HcBHMtD4MZ/6Muyvhn5uU/eXLaWYJAU1oc1wU2lmnQleaCJls5MkyrsJ
WznrZDJJHkYP9zpBVlajZc4FIsSrswzK2+mAa/DUACcP8DVnKX4X2ip3OWSd2GrBCECYm5dgh80r
MRuRCNgH4SzJv0BA1r8/Ich8lIaJDq3ZO5cqiDi8IuSYPJcgHKVKA4f2lehxm8IUJnzmvF+v2sCw
eFb0af0h+f6T3zX99xsMfNFs+zEpMtP/kRzKvV0bfQir67J0HVM0bwVb04UeOwqf2gUOoOd4QEbX
JZyu1C/Z44b/E7RireAIL9BLuzEKHmQenwqs8rZcA6J2i0I6oI+8rlgc8mWyu6APLOh0Mgj2M62m
YerhP0tiv8rHoTGNX1tylS03eTiVE52M41a9/J6e3jsGY7nf2GtDEbk0wsAMaNL564Ktb8YY/AGs
IBl4qhy4mfnHxtlBahDAFq61vwLKNnIWANoctMSctbAe3xQznKi2PfIitEBzWPqVW/Tq9mMnQQgy
/pgKq/N2/gNiQ47ETHLD0CdKH5kErFRxJ6sKHTmtipybun/liFmHvXziHfopUzOFbZpT0sdZqbaJ
Nq2e9s3Nm/PqIjY/2brRLF6GPw8T3Nq/nk/CtEREyzqIcwOhBIp9lJxsnDe6hjABlPrnxw3PG7p0
DC7Xx4SftbHwSPWzUvVQ4HWdBGd7Mwmbjae+cPixMexblD8P0jn8D9nir5LGUVAWUAvG8c+eRGOd
5CvV4T+lZnXl85OXfxzdSv/xzAWgDnTeQAz7W3DJeJC1kwpam2wkx/YVZZRwWSOxmbgqyF6ZZ+Ii
qlgwpRF0CHuEm4jcBKBv6QY9lNvJTPvvNg3uzwJHCbrMEVzeuJlROh05lv8KtNVMhh1r3vhYQgEn
omwswSrtrvB5+tM/CvvqEz8e5oe5yLF7/uzVmZchqquFwS+7WAkUDjeMJrx/YVatiIarsLLmGNZp
7vhauOMCdfIvkqmZ0rxbz0aQinjy5KZRbmJsyB0uv2vNLPrIOssKaAqGkxEnHHJYa0ytHgZWB7XJ
7XoLPcHyA1FHX0CJAemN+evQr3s5somZY0laQLFo1hEA21nru5su04ipF9SSXYnAUoA+oC06XaU5
jqqbFD2EcQYf6wv4IfKmzXMbwa8EEe1ec1TcPnjTX3qnB5YTA1CHJMyVpw5BuBR1Rj34dnE28Q8V
gNI7sD6lB2HCwG9T54QDWyq5cGCNK0gH3ZfLMgkFKInc/d+YePX61CxT/FPVn5XRLmoYYB5YkuRa
EcuDnU1QhtEPEfXJ5xOtZo021DCL4pMx4KtxfmYtjDIN0wkf+GZ7LUxYHoT6jl1vnDjnrX1coTcs
LVjphcq7m8C4YJFaUI9k0X+3r7TV5TxBbbJ+c1N5fBW8hJTBmNL3JrIpxZt7pgJvrUh5HOfDe0BU
wjRE1VB6vAKKL5BxYdWjYWBqo91AZs2ZMx4Gv5kBkqJHIOp2Nggl90LVoRVLeUh/8baVJ/Q8P4IP
3AfLMT56hn7GNs5f8Ivgc3jUF75nGq6GvIMRHXAypjLadKwO5CtaR1JhNM/e23IAD155jH1E7Al5
Sxo8Ijzaovz6UR4QsUAamx7IFVBoBp7ODfNNGrX/H8uGwM+QHNWGZgDcGQe2vbR6YgCmWExQhJdF
OC1+EVibW0fCwDQRD0fkKlEOPwDr6aLG2mqXfN8/utWp6LNcPTagQZT+1zmeqZ975jQUeA6zTpTb
kdhmIfmwNSy0Fl6H+wd32gh1z6+L4yNFadRgVF+M51sf/tLKwFFXO5wLCBmMlMyDJP4zD3KpEz0a
dVtqGRDhc88Th3Q7XdsVaufL0XTHJNfrd/pXYn5KgZEOgA2Z3rf2BzYCY/Yf0qXJYVLB/xwFwr0C
bOXtdLY9cswnhc0TQLHCi4GNKY/n5VfCX5o2iEQFnWDIFzNrnVV4l7E/TurswNzRYKibItNk0+pB
l3ccLy5SLyqJFhh5ThbU3Voezwh3azw9YDVWXk5e+ZesoHgOcG+yi2OqqXHYr6QgSIc3vE/nKixT
NZ7tNz/WvWbZ/3tdbUIQK5taJk8j+5Nt48pdQijbcryWVyy4vNgcimLjN29mZuKvixc/9mfMcEoD
4R1Uja+X713mkJ+6yE9OatNgxTGaMxwSP33i+l30unTBijxGJi294XmnPs9YOTZTpvNvMju+b45/
XanLp6kFnR56/+f7+LcsZ7fYZyCSzKoY4/b0g+xY+xEt4jp41AAvjWyUhejkuYz7sJxNmkFUAgJM
qITrCXeTajZPDc6kJuOEnnzCEV3xtGoFeu5dDSAF+tTofJc49RkyI5AGrBFb83ajcICQnoXYUtcH
GMCN4mDQYWaqe1tkbcAWIi4Mc979X4Gm6XbUy5Ngtyw7v3awAE/HVeoV/22QY9bA8n9wAWjR0X9C
1uHQAa7HL0DRE4P6BdEtn0bs4AR/iRaFk9fRU9RwZIh4c0yKr29aPAjJ7Nvkufa9wqIHlwObX7wf
j40Wbe3PYE895UWA55polUHxBCmZTilE1uQH5ZrR4m9oTKBlP81PhSZgq8Lc+282YsY0Sej+5FKg
d4KdSvdHf2xY/wccVtc99r/ZOQKFcqVP1xyov3/TEVX7iC3MVv/Xy+1D/dSrrxPMVrxNQ1M9tvKK
8EYHWY/gZ7hmOdAF+W38Q+YTwHumMNrofS0uKHRlS7o6UTWg1nTu46s32SJe4l1jTWNpUYpNh9te
jkwbOOU8Koktv0FbYEE09g5WjSAI2ZWG82Llwr125kCxPO7q4J1K+06WYu5MSGjsmRRowrYpWiUg
8cTx2dDGPU5ISQbB5vHaKDD92wS4B73BjGlX0Ekm+Ib3MCjAdq5JTgMdSN1f5nzgSo87hmZ/lKbb
Rlkj1y7OvW2J5vPaaXIVU1cUhiq+gYQjKxbPtDyFceHWEf/e+NtlsDhyP/ofGxdS8/issqI5Ww+w
8EvJcYkq15eAYjwT4dbFDvOdvvYP+jD9N4ZTanbLsvw0MVjDcNxO18aErtNGhFQSuZfysnsn0jsL
YwEdGuy7q3R+QKuHk6uK9sayb3ON6cLQeW5n0fkN2RtJeyItE6/GBqxZoqtQkeptPIDNvMoL4+NG
vY1s1fEwjad48G20HdLKYyJmaIFEQ2I2Uxyb5+XSfNxjqR6DrqoVbSUnNEW2lLtU80+qd5+wphfY
AVUTSeXfH64erJxCUBeTwnEfY0rgn2HmbTdIfAEssGJR1cWeMjyt/u/j0q702zuSmblItAjHaxgJ
JVOWTKUy35liZHaD0knnpu1jnAztmLQlTYlAofkDos8SVSYikn+fCogGcU3CH1RnOL+Cr3F4KNwF
CMPWvJaKSwIPIG+hp54hP+UMsF/ll15ksRc8lPCRG777yL8QcTUlB4FQklUrdhZEiCp1Q7YfgBFS
csgtuqvhaB/+2QL/UrDB3U35J5y05AZgteOh1k1zvz94ubmgnSWUYpsC2dQ6RckoSBLcTYI04uRs
zmgZevWwcja4AkTztmz9Q3w7Ay2Jfdc/jTFHvI8B6MyC135+q7VwnPLTNlVKwKw7St23ZfeJnIA7
MM+zKeIO+i9Wyrb0CJTbg+SiAj7a3dfnqutjZWjGa59GyLFM6o8JsTQg6IfApP95YNoHZu/SO/0R
Q+HyyZYMVGF/ptRK64vXwp+87iPw2duzPIoeudeCXo4rg4ODQwFDomSdnDrPMLxT4OAr4QXL+lLC
z8NeJVzCjUa6EyfXmb2JR9P+OidguFYOhvSEFftiNL8m5hLzBIZWz2ngQ9GOcZAURPGXFA2HltVb
wiXRhpas8zOYE6xnd6jLAKD1HpIahU6It5F6Tb8HjsOUuKeUnODaAsY/TpcYnwBhJb6A2XpjUQEY
xCMQB3lYVKyH2B2XPtuH4yZaDSna2G1r06Sm4cunOOi9oYvcFL1GNtvSFciteU5NLvTl1LACnMr5
0xw8DVQJKdxdtLufHMGDrSrvBYY9thhwTxDZV1KIxmprEJvZRQ6nxtdC41uASefli7eUnrZAiZON
wOnBIIQ8psKjn5ZFXFhzKWAgpLBv7JW6FMjHN5wec8AxVO2NrcAwQz0gJdmCfqvJbY5VLEKeR+7F
3H6w1Q47aQ8rBYHM+QjBukAxzb5opOiL5d8iO3dAIuz1DgD8cvIThP+ZjaSpFcjAo1pbYdbEA1v/
7ahspoDC0Smw6J4zi+6+AmBobSAWlpBdC4L1731moGgSg/c7l9v7PmmeYtTOhuJjH9vxMIzg4LK9
zlDV47KPRGaF93BsrWTpx6+4VttjF0JYvVYTJNDB9E4YdMxTOiaiZHVDr1T5cJGGx6LGAX3Ye+8H
x+XttNb7dbzDIo3gIKJwykOKIvpypVB9tZoaYjylYzllD/1UxcrEtHyHvu/Eds8pSDsuIUEYM2Oz
gB0eQD90aYgb0u1nannvPvsCJtceL9vMWF6LPPDPK2mhuhaRNWeNXEVBkpekpFwnC02h2qZ31n97
M9frMzarYgH0X231SVD7N2JnK3sIHarX8y9p7E5+a8djZhA7I4hktxsaZcYIWOzEHG6lOVwn+JIq
qjSUrvkccX9OUkthAHLdRMo5FrLQCDVsD4/S29/LnVRsbrbN2bJGeAzmoB+LIYCwetrBvMG93R4v
DBjqhLpKY9JpzoBZ+CPrw/0HFF6mN0A1S4J87OoOS698asxOyC4SlAJDH3qD5whu3x0RJUcRrroQ
N0EdMd89yAOXyz1q+3amrafAdYKub5KqaUx8GIK+6k5Nqy1py5ctFiAXNnskXCbl4JvCmNklhKHz
ZCmVAo3T/j5a8lO70rrpwbwr/6D7kPBo3+1B5jeIuJf4nQxv5gKvEb85Mabe5H7vrDA2oL5ZrboL
2yE2avPBq5igePQV54aV2xjM4/KqhE2AEfo9PhS013xCeC2qZSovDdjzw8woYuLdKHgEXTU8jBsZ
7e5AN/i9Pl7Bj1Muwh48IYT/XPpA+7OlaE6V98MQ0IACgfYLpegqJeuAa9o1Rpqi8ASy2ubYrahW
CeBkIBdYUGxfPfNvewMh4k/alSg5TCBIc8vSmqx87TpuvCAM3NVKyNMqlUElCewDl+3HJeoLinpW
ZUHmuCViXbgvreh4Eu5QD+ptJenoD9Tf2psWkO5qBcTIX1dEe8J7NGOU7aWge3ORur1eewUUO/kC
q8y2bhRoejnE3mb/w/W42/Y31CpKEt1+fg4Re70iHNKsmJ0pie0oWrhhixsSH6v+s7Wi0uhXbWvv
4hNV0Z3pJ/gVGqb/k/LNxCOOOP+HeIw12zKuRW6Iig+zWEf9bST107XqrEU2XON01hyMmFf6r6jz
YWyDAKTz41TZtdixIPrPtJ/u+SxvJ18p+pKfHdZRfMKIfh5keAPSrnzatCDhQwEvDReyMhBpcaiW
FWEpzb2O6sZxKu5aUKw4rjBeN32Dn3jlNS0AcNafW6oeimYU0oY+TvMyaQlbr2Y7aVorHqHuLcoz
ogW8UzhAfF09uLAo8XKTlLJb2Q/6oidIIYrdNRh65/oNnYeiURPl1ApJr8yt/aSoHlrDAh88O2qb
IsFMtOvMMwNAo78/P6evCqx5X+oZTWL+5ShCX3S8GSYMVJa9BZ4WS3eEuJ1lALv2JfBWVZOXtkwZ
nMaBssZlsEZrtoyqyR9GKXbPL95gqGOWVbuzxSpCRNt9zxU823bbz7ClA9zM6C4kLiOpB8+RWSS3
UpG/8KS+UpKx3AOj4ny3hZYvltp6R6If7mN8EWIGFZCZbRjmM26eLigvUCSLhpm0K82MZOZbEqw1
KNwHdafH9DA7fhXUN0YxzMCn/q+Zqtt1sOvtpYgY0pZV0FltTTn9TAVg3auSUV4m+DH7cfibSxhH
HfxT/uGXBDb/fWmCTTODNzs+mwt0Ycz7MdWGOmDWhtIZWN8Ndr3QeiyY9BPpi9PjQ/AHRzpUy47W
tRLDXiTE3dNs1dU6Aqc1jk6Nzk04b7E22l+7BNqiBoTjsB4ibFMlvdXgemj8rPFUfZOJNB9cNnEb
CTVvkwBxH1DeiCjwP/+WvRbg9dYl4dyyqkhXefmd45AetJrj9fm3Qi8zcDPDZeDjyf2gBKqL+Eqj
58ACLIZE+xTfp5jAeyQTvja8tXKoh1Ggo0LUypd8yEuSsHsfpe6uLRt3iH5XwhChJP0KHxWBCiqu
OySz/v24Y3eN8VozztgzQKveOuC2l4KQzTMElsBPpl3fJMmX2Tt0yTOLKp77yYtpB9+ohMVoSJ1s
b+M+MlRUZtfT9DBzcGe5HRecbRpyDe2Gx0UEBjFddDpIcHNAr/lj42bgUeggHs17SauoiQtVBQRs
2BM68C0U2mMK4gK+xWN+L+sGh9RXVyZReFruh38xtzb0W6xDA1lOY31xd9VXzU579UXiOp6xQwj8
NwIe6p3jHST7xUZG+M8p4ygMZ55Cg4FAPdffgVzh+8jXF5OEG+68S+Rh4mHea0y5fp+JxJwL8G2Z
0FFWs/qAvONJ/P6SXmzl36J7SHgetAp4FJKy4cBnOBDiHA3lHpMH8NUFEyu7k4ABz23+vvJicxwP
YvkzWhNfE/xLecQRYgVaC77igp95SD4NkMqBO7N2v6+5+X/fIr0M90ilZhzeDYsaS0wYzIwWIe+i
mqpXQNXl93sIxXbWQ60vJSHXfKumdDT7yEoPAlVSPFopCeDg4Kcjq65KLP8l0HzLpWYwwJoajL8J
59T9/bE+TvJ5DBG5Z+LrDU2wCozY/byTVAvt276weQ451Qgy0xZgbBYx42M2Ax8rBejkiUy2/zXh
XsrQKucggILMq8Piwkul2d1GZA2DPy6M62LufUCuD0Y4ueKCdh972EBHyaY5bZYut72wv/mIfbJy
Iq5es8CZ3DoUlEURV8Awcxib3gcIKOAmwyFqHrq7IbKVc9a/16/rFr/1qTRKW/LW0zll/Ebh6G6n
067sL2/h5VPm6j9EVCf6vHEYsVOM7UPwMd/aiJ86pLAQlsmEOYDXJWsO1vDDcnmgGfQs1yerKexe
nbaL17Twhm51aQYQTrATCUaqxe9duehOLDffifR3yFSAEJAhFGclbrsdOljxy/4VN8x+rfX60ry8
4JKQ9QOi2UYg3rxGkJjQBm5ZZ0nAv7t8Qvg25yw9M4b6ZLq7TPbwaWS78fQZINBlW7WAjIR4x7Ub
sA/hK3YtHxqTgnY+AY49eqW/eE6Ha8kgqEtaaeAkMesl3lQLJBgoOqy8PIMkpheia1bGGMdqaAmm
E5HLhMp9YbOX+B/tM5UaiyHEi1On70weLyJMyqAzWyzgfyeBmxZwJnOWa3i+QywZxcHyUMXm6z1I
E6Hh5mSKWHY7HGFOyn1a88Q3w6g9dC5MTrzfyXXL2+6ICptmGPM1KfI2kihex6O7QOm2WbpIH3Kg
G+qlOvey5tdHTGmm/O5s5/Xfp3vVxz+udVSMcLbjmAUWBXCv2ZpBfH38+kieMDRO/H7SDTolVI/+
DsF6DASD5+Wy+QyIO8PkW5fVKnmXg35nXbjT3Q9ODZllAo5HA9CJB3yrXqRWUmWWoA4qkekelM4v
trTH3s94KrUDJu5JA1rhIKoGWsS1NeZIG6vuLQzLdlwOA+uwxMtWA9p2Ygf5rq/KYDXUNZhLl0iZ
CmkvCL05/fAf0Cc3oFWOCdlGN6PlzgRF+wgvJx3Iu9060kWytjBNKsVZnOqbhqlGVa15G1HxRc+U
ne8EW6K8EcoSG5HQPTlsUxbLPZaR0Fpsr3M4UBR2+ACU/6vwK75z3eR06JtahY1DKITgpONfpmjQ
58hTwCuD/7bK6Otmzn/f3g779bCTOmeRXSJizMrZZnfYIHI0w71F//KwXIsRcxZ0qxOLB1t3IyCD
QdTarZHK43JTOc3Er+yFIi3wFcejsH/+K9ucwqFwcz7Wjmy+tlWyfA5HwOG02lwgYL9l2Cy87JS/
tZo6h5jLh3rS0PzPVl1xxVK44Ck8kRIIsRNYRaunZ8qWipd2UCfxQ2qEhLHHRN/itowrKetg4yVC
hTdQ6nbiUpJNydbyCjmSXL39jq2TLP39zlKpSGqzoXdgm17+Z/RH63S6BAg35WGtYastC0iW4+cf
2mA17ClFOwC04+bRJsT4yexOzvA7DuJvqeYVMq6eHyFecYFQZylk8iaM6RaJT4CTD0XvwK1Ovx6p
pX5Z+Yy+gUI/RwQaFwJXVf7B/aDtYm/pRa/bymgXIZfpXxV5YZG3W1jcUiDHA6IHMGbAzkXqle+e
4aAv3rzGJTWfjdTSkbyLpLvUM8ISEYsUaUj0xPLyBpKl/YAhHuiRWqqZ3Ke7hTckQXSwWgKb4/yo
BZHnoynz/7Y6LnOfo8x6/jxV5eDVHlSp/KsR1JMO3uIhGO8qwJNmyBfPxCjKkA1XtWm9Hf8nDWf4
6G1W0cIWav95xKrKdA0JuY346p4i7ixXRpcsFWRDGuv8q+vtY2mTJV/Zh/sWK2/v6UnVEMWAx9F3
4OtUmMcaH4SVlQSas76EXFP+loXHzKBwvUcIe65gkYIH27n8l5A2D6QJ0968aLIvq4oYekY2gBgX
ZL4O4cdn6iD3Dn/XtVUID8XGuhDcnFKry8r/+c32FPp1j9CVBzA4Yax+ezBZuw9l6NxAZw7GmiIR
nIRjCClmcLQ6wKMvug34mH7cpemmzcem4sud+tnjzqizYlDXhBgb4OEkxPBkIBpCoTKfEDv7OOV6
mOOxtL7++pnWfVyzarrVIUdYVYF8OrCyfXEC1DTbJ+akGfFeFqvW0Lonp/yqKxXwvaUKZAuh2gD+
N2K1YOj4B5soZrCbuT5PJW064zzYj3O5HWpd9gEU2eAx+ZAOV+NBmWzJ5Qn+4Yjh6d0efqfLGSTJ
bL9Fe/qUwyGo6RKqnhvNbKkSGiRzV1fiQ5u8n7Zx6/O+TuWs6nRax1oW8O36nJhLHRMmic5f5bWZ
0J+M8EXYD/py7sJ7a5JQ3NpTsTn37EvYkNXzKPb0HIP7Rjh+pDu7nSwISu4EjHBG6b0Qp44EVh2o
M7yijLStg9utiBNzplukIM65VJ5TDTwn9I9NK76p0Y6/aAmlCda+4ZsdBGG6Dnkx7ie0Ar66nUOs
kFEJIciRNdywPnNWh8JsKTMuXNGwKN4t27nbNVlDYRthA2n+SHKhohJk2AqIi2sbuZq+jztasxnc
dfZJHgU5RFBAuiHOJiMetZ9QQIzrVcKW3xoGcz0IBBYTwE7PKul3rnTB7JnE0kK49oOR0zCWQxDA
4L6pnKN0QAEiDS+s2apCJWRXWEVpUqrfr7PXXqlluHNg/EZjcljdGzur025/kUA96wLf3BjD/Ika
drWo6lBchJrZrT3+Bh3T0W3I5XCFFAIoL4vHr05EtVp6i0IkDL/Z2SCx0Rv//oUkfsNNhN137H0y
jbqGVIvkZxDNld3nB7LuMvigDUOku0Mc/V+SWiy3H3lfwGrBmJL4rsHGkNzlyZmrmQ==
`protect end_protected
