`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
LlPohJeWtELffanTkYuIMJWTMc0k8muhVXamIlAQraw7qfV2e1JlMuvjKKRyulkxqT3oMnJU+Bgm
D7Hk6dOUyg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ganGGzXxfBNbjBEV4j+MkyOm4NGufMSfpA5HydzYXGIhJZQkn63X09pL3vc9IPftjsKEqOjxUFqT
JfTAYIJbk9ub/9zz8maIeA0ZjMIFi1IxG4U+i5MxNd9eDPdGUgOLPeXrUcTS1A0Odn0981gqCUyC
pacfOyMjV7YxMfxoqyc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LHzGoULztAD3QebNfEn7qaKC5YzOdB+jrZQFfXU6orb92WACedqNAZXJuJi6VI8OeiPVXK+2xmRs
QxsisLSJp3ufnMqSondtVGmTez2ll6usiN/uai2IHkJpd6J41f9eT+Xdv4aQ+JOZgKxYaPEoDT6p
Yx/HXqa0uWo6uSv/wjYkyti1TzHz7O/AaignghgF7keT37APuiOVxIS0nNQgB374dtfia8CygBWY
OgUJRWUgoqhJ3D3jfGmls4H28guvVPhGarbMthzBixTVZQr8BRkz/bvBfn6109lIyYejKLPC0bne
yCbONSjkO5tv8bWUneO4adTebDZ4tkqWPmGgrw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3de9kypHUxxJrPSWTmVdpBZf83ojoD5she9KGy8pq1jfuDunf+0HNmZajGvaGKTJG+KtdlAlytCh
EmBZrMBYWJV8iFKPW7MRX8J1Cf/LxebRiahLL9xBizLro1JwvgS9z+2HEFRhQr9io/GGlYFQOO7b
zx73j9Qjl8pvrV2q7os=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yq69wphK2gcaPWNc+rTv2q441AIQCNGsOoUj5ExB2neOJAJ4mErWpKR82OyaZ3R0DR30En9EL2jt
hbODYTmPoNcVaBI8GnNOO3pGzycixTHa2dWVf2Crbpss4j+bYz/4+fP4gNsOIN7bxfsxb69lamcB
UY4574z+kE8LtB+RurkYjiBEozAX3TTWdnEgnaIry/F4EfYvqtQNu7dCQUAsyQCv7U/FaxfqUwdX
NCpV9w6Yp929O1Pq4Etumknq3Usi91aMrZFOV4xiWRiiU/onMSvPIPf8hHV7vKXFAwY1kuaOSNMi
VeoJSWiujlp+Pl0gXDBJjnrhzSJzqgjHWnhWKA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4928)
`protect data_block
6swAmC3uQKZDC/s8kR9GQLiSBiXevrt2MDZkPTUgZS2SEydDIIPOrymRREpH/+J8sWMmQBExbQkx
mN7i3v7lRZTXsCoxV06fxLLiGgXTEgzahF+ItzS59zVKfDClOhseu7XPZzE28c4Ic50FgFu83QQO
Ne1vOMJntTDeVyp3ABSiuL6tk8rRA8KVJrOzp2WDeed6B0dl2YO6FWfQDpo74wfbfep9ksdJHlow
m4yITUdQXD9Ey15e4jvqWO1G02Kc1tpWC6BbuzdHcskypjul8WckGt41ut4aS4Mi3J9iuvYi/xR0
vNUlgvHhT/gXnsOkKTiQ0eZDsKEWYaTbHppCwJfcXj7whPW8U43qeKLr4TGY3DaQeCyU2LEXDAdi
GNexo170C5vREtMmvDxsz3NaFuGqz1uxsDAo6xu3ZuF9JXBeM6ciTQvPPVByRAhfKZorBtqBhOWn
wuMTgs+sT5t2wwQBiwQfghj/A1s7QBZwLlQfS9fiHabw43Mdka3mEFREo7xkqw+R1jYtV5TmJMdQ
tRtQEQVfbCp6nI+hKioe2oK32crxwv0DC2z3T7ZrF3E2bBb89dGz/nt28IUi7nnJBnSPFk0Z/9LJ
Xc3glS1/efxa63TM1B0ifFsDiKPHx4obBurlCCixDEs1HMRo6GPdtXNctuzASZLOKBYWyqq3X7bP
Iv4ECwhuFHxU9JX1ZC04wKGYotVpIVzZ/TthQ/yiyGM75qhyRb24F/D6ugwYMz7F2emU0KkQ7195
yqGN3AlLicwTen3Vf/kjzcI3uJ7mjNxiQtMkrW1GY7pb3Nf6xdoQw0MwDptZv8yL3LgjLKFdHrNn
KjhHovNddXbSVilNLbrndHd29eOW1DlLp9T1VFGIlFhNDd7A0TGrzgOXOVaEeDUhukWwqO0nvbf7
choRPu6ZqBCe8KQ/q8RiFOh/p0q6IENiZz3/y4/SWEk6bxv42z8lm1X3uEczMHuC40jKyOCQm7Hm
rZJnObQXvb2xiqd7QRs2WNFW47pIHcJYAQEnw6wjKJcORoqlVHqrcXHNnmt9cpOtHjxvLPlxo8he
r2H4f/i8FB3mRRNtLpKXK8nLo9The5KYY8qd1hsHLHymxRtl+OPZ2ji0jP9BHJZDYiEHXajvCG8Z
diLks1fdk0Z/FUtzQASe5vC2+dYEiLgO4BydEsWLgJJjGRYbxdSnmtep+EsGb6lJph7usaGMQcNK
lqOEB+PKZTJrrdksDK1O+BgHxH/FLpbzMxKbhm0C7/XV0xa1VNGGGOvFdZpWadr7m+25u6bifBYI
6l/OdpXTMCldNMiBYxfQnlKQlYVc1fgDixFwj5wp0mdFnLf28jburYmvuniy+r6fGjfwL9w8wvaB
UKcaWg8eIIT0JDHCCrXFEnoHFwhTT7DRLL4drP9ABX/dADauVc/lgZmT3wlGZA2R0DrE4mXw7lgc
kYwvaYGnxAZmQ++kJbTFtaAaqXEn68L5Wg9ZlMrO+VJC/ngJ65oifBafajCsKCwlK3IsPlmdCQpC
Vu/IYnbMuOtOjjf6oY91uOeE5Ej5wLAtVYEVdOgAwE/4IxRSd5jtS4iwnlLeL8LBPuo8WsFIhGal
7XsdNBr4kA/KYJJH0z1xZfQ+hRJ4xu+Zoyp/bk8wpt8wvHzQDD3mn7eEl/JhFjuABL/K2oTmrs35
tQWxQUpDjf6le/MoFfWyR7YVc0mCqoQb2sV5VMT2HiSUAhxp47jXTd53IljM6d76UCOGSpPfTeGX
w1gnDaoDHjJuaFVGaifs9lr9S2+ZG6ll6sEsZ39VlU/LirfG8vXInGsARRLspGOSL6oqiY9lpLzP
px2de6EH0jqq3FUpMBH3pyf9UaAw1yLd4ISEtnjhtArklMDpK94euZKqWOzbxVnPpwI4I/I2jk8B
mJk88E0wDTIfVUNEAGbjJhWKS4ME0IrOvJa9Umnv2/Ics7mxFjycxOKarkJMVIVkRVqVgCyT2SrR
gO/6twcMdl52lranqahrqTLxexoi7aFN6jzov0ose9lXctYnzFFK3VdypCAI66rsp6r7KxsodqPR
iWPA0jfadKGKf5j+5PBafQwp3vKCAPVPsJHFD+7bwTZYCVxfCKlrUxiMbmiczN+FWYtZdaHNiuPk
wcb/UtGLd8VtyRUYAP+M8ZUHwtz/pEDeL+AkCmTbnyuHGL4+EmrHsAEO4VLSAHDGPHC7qvyRueAJ
CbelO4k3umwjygWks+kAowVs6lVORHZ3xkad7ymR2iXuPJLN7J9FIeduuhgaGmJ3h1QdIH8zFEBb
tRuGmQt3DfuoFmRW16F6Q7gb/Ow4e4xXC5HBtpaevLUZpEGvZH98DPq5KRCPgWI3yixlpPh8DoVS
s6Yl56E9ty8zJJrHuNBH16QKrCfRW44jl2FP2PQ7qSbDu1tx+l0cUKO5ihgSvGva7g260pFkpHTH
c3T9Sw+g15nrwnxtOKgHmsX0BlHMynr815F8oLbGglP93PjdlYHW0q4URZVsm0KqreJAoXya7/TM
iKSGhzJcCSXOoKcQAg2ghNZuT9rKlqH3kCbudjILtIhTX7JEAYvtuUnTfepg7+N5S3TDQidBheD2
pYJz+2CWC9BEDFrTsql6BmiPrUVS9UWreli9EUFl5a19v0Bfp1YBIC8nu4xQfY3iaYsEYa485DTw
tZhkBNPb3zDfqL4wBy2Ckvg4ZktGULaEbdgAV3oQfu4MdnJ9VPu/qSq4DrNA9atm/Qz/nInl69wR
G6mIOj7j8YFJCHkLim5eMAN3HbedfiA6JC9/xV41XFlxdafAGBcJm6e2tYqQ090RKsO6Uq6qmezB
hzo//HeKoYVcl1FPOq525mcrgEhsgSQBd7hFXmXuGCh01oP8sg1N/cd+c6ljeNMLQP0Dg6z+X/An
T/uCqCfxaQd3MTT86xY/0V2+vepgro8+i0MvSnw7leVbrUwNWBZiYbRzJR/qHfCHRwOFnZH4ZMeG
z5q1yXUkAY9cGc7sW1NlCWFfW2hFfwaI6aJQ1lnrrB1sdP6WL0WV+BIG010MgK2yLMwEvXUGE5X4
zgcNvEf9N/lFKNy5+S1lQHraHxUQQj4eDlQ8kLnEIOpQw4rSI/CGdELLGy0QDKDmHeHubY/V2xAZ
9ebShtI+vEUcSeZmyaCWsc22TOQ2K6SqsunOeLzDeoKbh2L9SAI9P5cjyP0r/fjEmnpYMmpEawcy
A/3OJFsmSyuH0C5dg1cwMLtmOa2P7Bo0j5nk9Es13p0YGFv3P10LvKwa+fcohc7TzzoUafO0DXnj
kY6ahWqZPDVAT5XS3LOV7XYeVN7yISMQZtgMP9oKp9rPjg/ocA+s9yDxmt4DrLhu2ydaFNCmWIvo
k2K1RB0wcns1kk/bzNJeZYHuULObFeV9yXzSbabJ0Aai5n64bPZ736vpBVFfImTOO2t0PlCMN6dS
spedMb8fOi3gNLvuOYSxhYZWK8IWH6eUD3sRBvJq3InKOU3rJ2N9CZXj8Kw6knb735TofDNN8vh8
g7NC3Sc1V0gON5cXKccE1yJn/f3f2CJubrgyr91S5wiyL+DUgyQ+YWOTFx+wY8sVb4IE10Vxo4wS
uxs9UavcnsJUq2ltm6PkcRqA3pEtm1+nfvdezOJKP0g0+aznBFayiqNqujXJTQOFdZsXVX9UBAiW
jS1DsHBJ4eQANuXb8RTQNOMlXipic0FEKGJdPNFpcbzuoOYVki+ZSh+D9PfQgq8DTr3+l2aAQJz+
3NhudfcfdSlYjiGNklEDprnR7UPchhTFLUqppEQV3JWM/Gc4DOnI090qO2NHAw+9MEtXkQh8OhjD
L8kLTmBnkJnQGRK8DSSo2MExaefqjrX2knE3tGnPmej8aaRZiAQw8GkNoEIFx6ArCrgKFyYWSo4n
KqZMuwVht+hKlVdCCR53kMIDWxhFfiy1yqp3GbUJ5ru0hWhtehe6xiwTPT/s94Hxdgxk+pXFyZEZ
BxSQSAofPIcSc853pVOreX+FgH8jnwLZr1RJczuG23QdeejGKYAtdA+g4N7e5QvIcdR32eBXmJUB
1D2KYZwyZNFdq/84fPAxzcs/+SiyDFrUpotCQdmjG2opTqsaf5yi+fneuWClmi0v8Bk9Mq5p7cp+
zLR1wSy7MwU7vhTLll3DcjLByKxOzG/HdHqfGWOnBRHwnQIF8TnrZxbhN+eejzaA/oGpN1O96Hvq
WxGdxDgkqDNo0soVOadnjXZzR/zvNY2uwKN2TbWXPMqZtWJBCg6OHzBo1y/1MErg7gtj0uMwerNF
o8gktn0YPe3+SCk1jtraivjDQXQKmvLhbjlvENifZ/0iOh3jwjwBOnEKh0xDc3DkXywyKAKHnG5N
LbKq5BIckuxVPxASWBAI4CTK7h1VSK4DNKqyL70b+n5u/EdU3/TfilC9P1AN1+204GeJhxiorTxX
kDrCDG2ni/QBOukVXSRmhJh4IyOr3oqImUXTRx9ZgLoHbmlaLX/+8qe56eunjrjqX+gAmArorkh3
rszQfoLxqK/uPWsYvyRrcxsoPJaTrv3sG5Vt7Wua2fytbpp+PVm748AeJTgLKaOtRAEboH8tC9Ml
vSJvynNKII68iaVPlZPbXAel83iwd2jfp5qkKaGg6LPoEfiqHF7RCA5mMNG38/ckUvTwmHNV5Mfo
WWCeNWfotGgUmGpjMTKZ75Fxp8bUSfBWwQcKmPh0sfHmfHrlnxUtL9ho/pqZ9lQG+k4TwXlZ848I
1GLi8rlHG2Di0t6/jU2zxCpby/Ebp5b7lBz64pozF8N96gW58t+jZVNtKUs6VUutlp6+BhW3UXbf
hojMFJL1+NUOLfbw/aymJZMaa8pQq2sA9MNQh28x1Q/FB1PCOqnz/y9itPbyIDXJYipK5ja8kKiA
LHv+jTXRidEtnc2Yv7vpKwJKDnvmw3H+hqIrphH4dMLwlm/1J6+9cb//Jvn3cokVqbgN6htgTX2f
8lT6KCG9nLZkApFNDtVJeii2Mt2ld4wP6GxBYQMYPBHnSe89PIEpzmzgLXrNvwRNNwPJ0WLQfR+V
vDIvHs6d8O5XqK77QHyOG9CMDWRoJY4DpPT4HUR14Azoj7xs6BiqOMrEBW3N5oGSeB7rV704dbrt
jAO3/6GVdzPQYtgrrbfEW4edihbHyw+CcicPlNJY6W/e4IoWMgSFBnd+XKp0lpZlenuumhrBErHB
hAQx2seoMcEDxmHgV0aIsUR2IxfftWRA5FIYz+PteF4fZU17wEpL5CRMyHcTqb+k6pKQNZsJ4Te3
uNLdUKpVtE6VBCMQqW/Z4GzP/16Pn0qVL4TK8ebAWX8IOWQUs2lp4xF/UPJX3I3mlKveb2rEmX4F
u0NlwZS2p8LzEYBNJzoFBbvtf1U++desdFgFJVk+0VU0posg/GANGxUIx/TGEBPt27xajHiwS94B
+S3K18jmjeLCyqhI9eOOQbUNkKTPOV26FXsL/oEvPgfwo3/2z39Cs7wv7hUIw0CB4exJY0O2JnpI
KdP1QtEtsZfe8AXlDMZkJFLHWCSHrhCQfweEMCs0nJ7QEbQ1XYRXWSOYibq/g5nMSmyjlnAobYuJ
2vln/WlUzgqGxOLZ1yz8eUtDq25HikeiGaq3xy2myoy2eRrzFg83CQcJBHhHTFzOTvjhNxPqQfgJ
XXqwaWOSGa9zfFajcoK8lF6NtRGT/LdhXKUJwNuTcu/iEF2kn7Gbo/6a10yqN2owxuACY0grxST9
EEPCfUAnxmvi+V5YXgs3jP7h06aJsrfON4lzKcaNjnvuUcVKPQF+WStq/2ZSr5g9SsHTPTZElbER
9P77albAbAxej4J8Wnw3Nz99LrPgRAXpmyTPoZxFeeZu4soF6deJ+lmWkoKesxcwF5Q9VgxrTJf5
+dzOi7+vLPCQcYphl31BCKqPekUFZNuu+BmpwTjkLgdNnmzjtsDRQN9NjtR+n/DPg6L0evVr/tiw
z6Vdpm9UGmxmEThUN3fceI1662sE3jtw8ta1GhxBk0udkNwpphlpsyZFakDRP1sM53KJcZ5gE1eD
rTBzUn4ZoEGdwYvYTbWGxgkLjkT2sxlaKssQg610PyZXTr/gI3JP67Ia3jmBrjXVt1CZXqqLZYn9
hbd6XIhs4rfI14ql/XH7xkwAyFYEEECfkUXTga48kx20rQw8cdMArjCGantNzGcXF7mBvCDSOyd8
zAs2hzFkE23KuUtltVttQTIwAGE4sb6TWjG9DsX4jeRnkxz9ikI/kU5OyX+2ZbaH0V5Xf4Up36az
s69Xegu/8vaMwCNDIAJGgHxx3ZtOiYXfDimHrPWqMaUr06DbKlbhbap0HdWd3oYbTj70sMQYWUaq
P7UH+YhEHhRFySdqJfeLgvviurAwOpPSKgl5KSLX9Z6pbj7rfQZ7jN/9KFQwyR3YJb188UHlkmFD
qkRP/skuT7V4YZXNNvCy899hGQA9aYA9Q6hoNOhlDu+26jBZBYQ9K10QsmFZvtY1CfaxZwSC2y77
yOSmi7i0QUj3gqSGY78ABM+J2xHvbbgIvstbNGo7SG4m6fIagU25jo/MJotpeDTZDGs8C+ih8X6u
KvQhHnkEdeBfy40yhuvTYGob4gXFzKQrvNc=
`protect end_protected
