`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oB0oVBcm3y8N2ifTZHOuxAaOLBaEaiYCB0P6zw6m8rACAxJLcWaNISMi43hgtxUSnkGDJxzgOl7s
BbAoyvBM2g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gvtqmTc+lqax4nLkc7TGIYq++AY27cp9q0Wg9h99nHyDbNdVbkLmU/64t/5tCPY8RN3QU+YW1x6C
+d26KQWmThI7e0lS+BJosV2dmbofUPO5ccoxsAJcdOfBiDecb21R7O2BHOFA5SbqjbbA8okBxqR5
e8721eiDMRcQTBWFXJY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cTs/PopHi+O+Ki3ijrqiWDAcWHoQA3ralIk/zghT+/cPVRh2YbOOisWtLHdzkFZ1Dl4kI+DRvgLW
SR5ZfJQuRs4Kq5rnCtpEj5YPkZWAWolcOR8yjUQy1y82Sbw3rIsnOMWJkzNNvcFxUpx1tXwfhK7I
K2rFetgg4hbnAx/qIF6G+0LoCEDKf+ga1YI/Gxw4hgccU1nP3hTJOuPwt900f9fb1ARVrKM4D+1E
cXt+RbmrmVPs/KkpoI2IYvKEH4z+zZGyo8xhhGyBelKUcYSGdVsYlLG44bPKyxj7fFqP8kIGjk6v
odDnmelYNQpktuvHMmAGWqDh1dS18EHmvuJlEw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QUwgcIuaQjTY7c1nsOyUWft6joXG2sEbC0Z2S9GtMId3TpoD4ItKSBO36e2K2ENvn09DVtuxPLtk
kem2tJgNLgRx1CGsu2GoUP7OaZyX6O6zU9XYSM2/mi6bg4eZlbD3YauPtjF3dPZq194bwwaulQTs
BUycThjzzuxoOlTsn3Y=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fNLiY6bOmkiEZhGN5tuxQwOd0+D6JzsjA2hVFYfAxCQPtsDGZIPeCBXhJsN2UkIq+xZZzdNylxYN
5RlI9KXlAQLOyDThUY1VTmo4Kjfw/qanAKpWVf4oEi5llenItPpaG+c/gnmMyZ4jQsaA46APgN9O
ykBY4ONKEdBl82kF8woPu756wCyg4DTOFYc/DaYUvaONYjBGzvUtmDarKCQtUTgXMWT5tNisw93v
yo8xZQ3lwRC71uzHRlETZgrurQW+J+S6A6TJUACKKysIdJ4pZfJK8ZQGVKdZlCTiMZLstObqb6/J
Vhjxh9MliXvDIHax37sYQgHZ3adX1z6m5JMsLQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5472)
`protect data_block
k5MF8z2QInftZgsmJ4dNgxi0lcAQFUZOLWxItIRW+J1UPXLjFLliv7mB0W3dtnWip3AcPitA14Pa
6C9+KH3tauBgAPJ2M8qy1Yd29WiQrpT8kpWwtsSZ+SnmawVUdyYowYZZWFx6fN4qsD33T7qAJ2Zm
PxuRIZMQ06oXaQgGjPQkCDG4SNd6NW7pwhIxI/JpB+TLDkN4e12+6EsVFwQBHnduAUEQSwnPOqHh
vNup4vWEgx7YiMt+wlpIiMXfIMg6Ge7loa9I9ZkfcXHIN/SjQEu4LgqtQggZYzHNObEfdATZsFZu
LuEsvBvakdmXeda8la9UzLslzHmrd8GvpegfCVCoDHjecnalKOaDyFXXlc3RvzlAKGCpqQNDN3S+
sGR9I6UT/zOIOC9BEBvaLw12UcgKLqLOj3lhNKVZ7Mxa40ACRr8AxCFxeO3m53xYUhEvxSdZiYu8
h+5d5H1PFoRBBU1tGoyp0p8mcqKQPEzbBze53gSApkFWUxCjb6hxF02Jn6SQhHez2ZS0awyIhgAC
W1hPYW13uSK8NgK78A/Etv1NURoxxWeO9wd0sXCYGKYIrC/xypzeDRKTBfpp6iqaIOlMPzyn06yX
h4/6SXpTIYtKAZ4pAR8PBuWsbWnBj78kmBV7P4dv68Pfw56F7/7kZl1t+VGQx6m5I7ZFO4FerNwA
irk8KlSWemo6+Y3YSTr4cVOArV1RFteR73hqFsSpdqPyndP34yJuT6PdIW5lI2Z4IB7eJZDreNnJ
1cOovmMOZuyHREVlFUKgMmQqxPpGDC8nzM/yAvDff0TZwv4ZdB75JXMdMmdPBtSXPBg95bRj/mrV
fveN7UpLulYJn2hTAGzf5shf3+EJM6NNlr8LdbtiIEobetVseF8A868YWOYfbNgKq1mshon9+pzY
h4XuirlEZZ7PCVGYl67alLucvL54xctuCpm9pENVnDB7UmJqyJwJaNgeIsbpCq/OSqj+eGAhPmUG
pRKqYOE/s/IlLNCWfcJCyuQBnksmZ5pALmGZ+CWjhnTC8vt0vSnVQFjNK2hzy1OevOaJXFCOcCvY
RsaRjRKMRoCRVAqY2d5uPR/6//mCWBgsiQXUNjKUH1sXqiCEGIqFENjUNOiXPn4vuRxhu5qzbBxV
D6LqpcTdx5OhVtxhuNMXf2u5bFyCZ0Oh6KN6m9nRBJJZC9UUraOis4Z7ncfxcw2qXV6eLDEeoe4b
MEEOCn/ns2uAUtpzDKl4cN0X+7zFiDOz01CLubuBBj/JlmoJ9Rm3+rng4tFZN5yLYpHVsnmWUFYD
KIOZPXm2/4ITvvH9vkFhMRweCqvfEoXFciJaWu39Wv5DYqQ4Q3gvHMusM6iMNuKW9uByNO74j1gq
+jvcqUxulmC014uv0Y66OHbw2z/++K7IrV3ikXBqslx8j47nrCG9FvpICB5a4ZZ9ppmSVNZjjAfL
qoZF8W5uwsYdDIOWrKXug1CHh+IzS6Rdyt1xW7Ygn3stITrFkwKLfedSJ3GYBp1U2IunSAUmFtP/
FQITzCz+n2JdarLE0KwFueD7TtYXSKiAjHFzHx0CZ7FNUBHYDJ8iciT3q0lLRPm5jfiQj4h872Ra
A5B1riP66w4Zt81YOob2um+7jWPWDArHdtjiFYYNHniwsngV3ymggnpegyXsjIEPyVGDAcOAbpzb
QIYAJWKbCc+z0kpf4Vf1KumtIcnKsR9PRB3D1E0MoYENSz1pVB46wSq3iWdAHWfBS2Q+z9L5yc7g
9Gagj5K/kgR7inGiwp+94kkN8lNR5zVK1JC9XcA9J4l/oRCy6rw6wi79DgXseiiVaJPp9hjKejcP
+5LnqdzDosSHXVKEoZWZCoIyQrrmDLJqgLEJXp4zpHRK9TnNG+MMjEVGiqmqT0cXcunLT62wyQqS
TSxcjcNjWUxGMN6R87+LkaBXA8nVueRob1iE5dNEPLgkt7Izr77d8XpimbgGq2/IOLAcSA8sYdqd
WJW6+CpJlTZZl+1uen9H0dkxGdr4LsQXaILBpLdi4q9LKkesvNB7JONrlADVZ89pM1iiClcbykH8
g8igfx/HysWrDHqd4jF0EhliqOYETR8KIDKpSZWplVChdfLUjHJthWG2AOpSRXRdtwtHXijs/uf9
JAX/6eBEwGBYYxPoAArXYiuJrhLTzhuQBq29Py2+ZIfbUxwTi524cIhiSC0+aPmF7PQTynG9jVq8
rQwjNy2XPnpsvaPK58h/V3FabPVDRJbfoX9OPCfR7hLN1wGDvan/BDwvAvhUhGtg2xYRqWZAe360
ALAXJgMMsFCzz1sNsryZE/AZge+pEfuRM8y2DNScl7yhaulIjLPsFQRFDI9KVafh2IqHbYjrVtjV
QLPRFdq4T+FN640T9WNZ8wRma/nG0dNfhbR80vEtdMP5VL/gd57KUnsThW+ZgYOicQVsJEB7neLz
SOPnvvfvONvw0J+Y8O7j2jh3hGsZ2jNgq0uCJK99U2sgLPMoHGU+7RpbRNP33i6Twf440T6ynOMT
1HYD6o37UL2RcGomMjPM/apKCh7Ejfm6Er2Yovaea5ZrvnlJNDixWvih+bX39QWHefmB84wl0NSn
L3er97hroGupidgAkFp7gbvUiTLEDl5WrJhaLVi5n3OEuEKniH5G0BsCB6f54VB2LqxVWDV5Tztt
p3bGKMeuiMj+kn+sAJEm7BU9IoB9pLJ5G5rj/HxfhY8f2/uwqR3+Lfwaq+lM0CG8PDz1ouJgs48W
fjuuH7lrj7T9F0zCbt4bGAoOYJ31dt4l5MUwS3XgzkrhHHBWbSs+ztyUS+ZBqsinqy0Uwak49Sp6
CtTGG0L9qLN8EsRpXjjNLQLjAMQeeVt0azWOXzIjNZq3wxC8qNhF0aeLb+qri1+gGp7qsk7sHXlk
0iPebR9+GfwEsvsmnQWNnV7glfFu432vkFjc4Ui7mURVz+HgXvL6AkAdO6wZicsiYwxE3ezbdgpl
9Aro00kIwibU2CvRFkqUPaU6bxMxWaxZwaOuTUBxh7Ytv+N6SAhwqcc1+jjg8gP4SuZbytRklvY9
AUDlXhhBXpKc+OGV9PG0Z2vjs2jiDM5LKqETMEKr/3+Y6aLC3P8bq2QM8Ot6FhAwKN3MT0JgPvHx
eUNhqdmaJtdD7HwgofvqAFjWSQ7EGosTL4+4o4rkGFbaETtm2H4JzF2/S1ir+QJsKmursRh0bxGl
QtIiM1TdefdsoVylBLUHhpdd/NZhTYonysZxKN9sllUv2fFXCIDZP6bXFmIDfHe6T4/vfLpoSra4
URIn2dQdGO2r8Zs61GkNn2OzbCDPUv5Gon+oYoBuGuwMjdwYQz0MleJnITAAOTX9fAq8f72Hhas4
esPlCoWXGvwFOcrWGtuY35spS8+WckE8YYl1XaEjreAG4WdNlmeKuK1VziZRSyguxRNZiQUOdvAR
21ssZjl/uuzxE1HEcjKly6boOq6RRsx4f+VvnTPlzmYL5rvvPQhHyXbmVrGiBWkCD2hnX8hfZDe3
e/dFQW8nbLWUAfhpOVtUW7XWpfNA33kQFFTkoSemEvW5LY5fRnEq6vs5FqfSSlKpv+7DQPqssB8H
uvGKzDAg3d7kqD5jAwU4Yxizjv7HDJM0kURtzz7dzVQx6GUspE0SUsITI7QYhDor/HjL7D3to1mW
/nf8Z0qR/sGVe+K+mtqdIJ/CrHLw4EJX29PNBRkt6SzAMU529otxZE/Zp4dj8oXgMfjgvHC/yd2w
aYT2ojDQGRmJ8m4X02MeihMQ4XC9qNHKiBOj+esJtpJx/L9cpn66hWlJgJQ0Kneo87sguWEs1OqM
lpXZJeZt0GDNFtlBa6ihT3tk7Y/hyZhoz716TI3strY/nLGuRaOhzF6jO6BsYjEb99hh+MjRR1rU
kup84MwZK1OxXxxoqxvRKj9dl+1+9/L4MVa+ijRn283hTSx/AMKGzTdS5nkRejxoAkouNoAWsTvY
Yb6m+UczshzlwBMx+XJxBPuPAvBOGRTRHuuNhxGtO5XexPE0Df3CJTdbMNupmYG95siRtZ+AJgyg
ib5/Rcr5PJqfylcGcOp2jnTtaEs1PTrP+iHvn5TUItk7tn2JDE1APGbdsMFXrQcoPL1Kry3OSMZe
CCUftpcHJEaADHtEjEfXh+oL4b4nLtg0P2paOyGRdPsyJMhkPJrv5PUwvBJfPyeHy1yffu7/3vEz
beZRwgOqtB0VqMtqYbBuNXbooKQWmZt8tpWx7BC/cpQa/Ps9t8lHVy7+BpQKQ4FJN/P+d2bcvQ0e
XZ6SMYldDur4SyKI3c0SwoICy4kqXGGpFu06oDmNf/u4D7mjl0zRM+wCNgz1iKwkZ1tDmwxqgbtC
AxLZ1sF5QYhN5L5Qhvkouh/1ZpA7kwPWqdQsmEjlsnGPhgQZujMca5aFZ4ArEFlFQkRxl86xu9pw
mkYQ8akzHmf8DdHvUIL9X4LWaAgLtlu+jDnIZ/zspI2gSDwUPmBlvzNo8fYpBuEEXDIUmN6CjvQ8
CHWIfkASPadZV2rCERkViXuEeRhfQQyvtahutQW74HfC4yDqodkbEPtXhzT5KWwxul+CjCpes6HW
RMLb1bxUqVUOymp63cGSy0ZSZF43gIH3xWcVIZhamTShpGvYCUuZpUwa+5X+B24nAkYy23VwSmB9
DLl6+PYReRfGVkKcmwaShn6phu2NC5WFReJcwur66zXxqdPOuqwmsV79AFTMI43vEi8010eJ7DjK
I1IfQ5OVBmtQCBERsCDXixCbFHMdom0a09GyOn9O684MZYoJjOzbPNGQwMH0VnkNtVhrZRxXwtnA
tZAqItZiWWUwCATrLs75Bg94qDbbesjKUgfP86BqMJxGnsOcsWMhy7zd7f/JQKk9rYN78WWBofxl
KXaktvOBwIos4aBGxFZnCarCACx82DMlwAmdd5NCBdEOE028QE/B0Sd21X33E+2dTW4RdA3tEjaj
AbRW0ceZODxpaQGPqTxFq1RqHOG8ZA6fHDbwY/fbJCIeIiBsMpOCqrvwOJygFJ+sz2rjrj4y9puf
aN2VNq0yLplDzriPtnoJXR41538TiWMFtHhs6ZfA6nfTurhoS8NnIea6b/DYJGfC+gfmQ7wmJOhc
nCDJ35tG3JwdCty5DkMG4hZI136n6FQOPgE7syYo9wpKmxRNJPrxqXDWFOoFqnUds/wBm+S5LOiW
2GIybqhvg9b6y96/ro07rqKUtYfIyls+c9bQ+g1QZ2ZGeHM0lwe2ZAZ02yw7BwxzRQOBFLbBF+j/
LuEIcIaHyhFhgfjoLkjlEs+ssIj/ror4A6fL395ZyAHp4JdaEPVAF5qpUvsabyC9ePE05vSYr6En
HmCrIo1VeTwPOwBvRRCvfxJivZwzrc9KOAvmZ/Lpwwtmqe6Xre1pxDG24COTm75IlhfVRb8DFxES
yk/dnOWKQWWU/DrTZ4bapy5l0TCLhmclzeibs7rc/P7YZRrlhosKbAq9N6h/rCT5vh+B3dh1vBbm
Sz3mQjQAghl4bE3zlc6xkjnUnBpUa/MVlCr/dZCThW3DCwYCgwV77rSGDNzmoZgEegtyT76DQnQf
/Ci0UeFvQKzj1Yx4QwE4oz8H55lpMiC+RTL7bKaD9SNkoP9kCPF2XKqPlDe2IJi6V0ozFNSqMcDT
mXmXB2H6OXHp8fBQN49v1V8dfRdk6oUkqDxw3f0N8p6IHMxpkPo1wZ1PHLWCLPNxvBm2GFt5ZHO7
T2vGKXcuBvJymYTK2IitWG2TABVp+CxSzZ95zhxDAkraQTlKkV0eA7jye2HHI1Jc0p9py3aLFIUw
dcS42xv026RrRQqHT9IPzO6owtS+HMGjfnlPuwuH1UWLFOP5jt1ugtBeoRGyGOS7ksS4/H4ewLZm
AN1A6F6oTW46+I/aQB8Zy8QtpK6mwv0/NvpB3GdzLBPrwgv9dCxcMmUF50xtDOdoWa4oYONkDzB7
YTOkD5yDsFHLsCkNGNxp8XG31BWxYvUWNHlmqaHTs27zLpxkVUO3vC4J2mJvX+3RghZM1l4iXsZ0
SqxGFCRa6n77B3UTgo2271HiiedHGIIsv1hhL3ZkIXxILTessekpGSIKcRe9/ySXdg5W9mWNsURM
MevPUdPsEwWBVu3yOAOqzO0G41ny3jFoLA2sT+JTTQoJuYgCYxElpv2+qJ+96ZWXx2IgCjVBGFTq
tqLunSIDvRFGZUvQY8yYPDDZsvDxaRhYYz9p/MgvEDth4h0PukrE0YVmcdWhQ6PhhlFwogD9f4BP
w1kpNlYWL20eZP14Klk9+3hDtXdX15nUTNW4iZHUufpqaiSnHlE9A6elt2/Pev9deKPZgTkJ6apR
Z1imRDoV/PhSq1Rd/bth7+6ysuid35l7EbWSdS0I1nKx+kxkPtQNl4OlPnIgw/SUKAb6O4JNhKMS
/V+nGvHWiqvpFzIlE4uo7SOYDJOvMJZqi3azh3pNJ97Yj78wZXL7qK7brNEmAjEx8ix3BehgtJh0
BngmfbeMNE5lSQyeeOAQu9VIU+XObBizCFx5PI19U0kRZVBKyzEJ+kTFASZEREF0XET5ezhr0UR/
r5J5oRiXy6q+T9F9F1tcufClkKAvO8O8EWZnsrGu4ZxtBLM2QdaW3+KllpJytVseUlhmmoFV7vh3
Ey+c4SmKn5MWljv91pMmPCUQFL2O5oR8yibLnBGhJEKie9LWtZsBte1TScvfSeABM7sola7omAHr
E9/sAfZ5voOWR2yT2pW1DLOIShNO+osgPAiZUOdCvraJufcdrV2LhBVaDFh99eFmmHL9lWI2rTDq
SmM3d9x86Ig3eXfvRSSdvlYp6Dk7liiFsbKk9F6z+tDkS2mxCIIrqdPNEtxqOVf3D9DhuEyNJI7F
VqThbg6GR0qmyyi9ZCTrJa8XHS0+ZlzDMMYMF/Ln3eW+hwP5zsxqOJRmDqfoXo9TuYxY37mwOVmD
Ha+i3p9UbI30+3a6uFQWobgY+qG2S+WreodOXyy3n6wi+m1+U+rMIoXGs5s2quWHPzC1qAxUBe0+
o3BJrG6aJFp6ZPx281TO2j3a6cQ7TCvkuHmrWISGXGyfSqftzvxRTI1mPVB0XjSEOZQsJ1ytIwN3
WXMMFUa5YEVlf1Kt8tBfKpqJvd51DEl27QBx5t3gJgQS9ALQmKGui+zpo9mJkeTuFlNQI66RhFV8
zjXVy+EE5PxIfFn/D2EHFfZXKN4DMdcHQeVUFBBYjNgf3cRqAzn6a9lTShVD0Y2wiuVeGX3a80sa
2ZPdLh9P7aWBDZ27Uh5rsFkCXLXGxzr5I+RU1h2Zi2FXIgev51day6bke4VFSPeX6eHog0z8qD4G
`protect end_protected
