`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
LJ8TTUmiOBnKqyjvrjQO4RRPbzkvS2M9GeuAkFspashmpAtxGwvgrO1aZTMrvnml3Hg7OONiTVBr
qBqgMPuSTA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VS+pTzC4UrAbiDaGN6TEnTI17CGxNxdh6qlckpQEE8NqARqTjDo1WCH5g6HIDryQp/sT1QkHbEn6
5mj9nTazAOK7GgnmgKocjkq8lF0q32xjZwMF0FLH7v5RX1izdrkxncZFwfnXQvZAHzDe8asem9fC
2G0Zjx01twK+Pi/IekY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SQXZM2ilYxsSFPzaDoBK12ps0PBV+OqjEIj8T2bROjRHckGx1sdY5BBdQoM6FGXkTBb3VXLM/7Yo
JZaDTDTmfRd+x4h12ruRQsDqB2ulKpaFqoa97qu/ld3hGnIwgeeZ0R6S2OLOj152soXnNwsQdevm
Wxsz3wZK337efNENnk5ABNR2hgwBzz2qSVqzhg6sUNty7s3Rhf5M+EL/N9w40otKJozm/JyNrJF8
Kyur9NcX25CpunsOMejAAKPkrZ1lYNZe+go11eoquQI/M6iLpB3amhmOXJNmM8ewj5Y4UieXwcdg
pqxH5VZfRn08STQbyduPpdDXAG9V2T/svxmerQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aG+9niuynvThoQAhMHE7UzEvUEAA/MUx/es4zLnv40C7VlW4fx/FaKfL2HyFn7ORf2S0BnWz5wHE
Xc45RdsSPt6xbOsYsu/T61cPgD+5IXKUrsm7FaSIMVY6lUV76x53GgqDecC6rlguLG9BPcijVifz
Q7UBbqQBsNNqkgczY7I=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
imUtdIAmfnpIid2IqETw9v0Xocy2YhdJnVPcIcedZj3U1vhXP4rjiTKZZtifPJ3Dqz9c0x20pFJx
sn8We1SepWbU2SJ5M0V8uh3K/bNecTNmWNDSVRa19NyJDqP7+UNXsB4+xt1TExJaYIXmfS6TweF5
V8mkuvfCxOd6zYP2bQcfb/OgR01T1q+ayI8lHuk8RRf9xy4jZP36tTsShOjKL70Mx2S7SpPHgFch
uuVxgmk7smHXOV+DCarfYQ7XykyIfCk9NHKwpIfO/ww4iBGer75F/SBwJJkRGwJCmrhV51z3g/rn
QSIh6UAMsRbFiGReFJfAj4rqxVeFiIoJNu6PyQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16896)
`protect data_block
Kaq6GhHnMONcEc+/ktCxtEzSj9AqfWuE8z3DsTOjlnK9ANdoDhraOBx0S1HniOtwgp94EtT8l0Ju
8A503VibFK3aQC8hGrRfGZycE/Zl72sN/eRBtNUsDGfm/Ri5NQf4HlEOfP4cZhu7GlmwKA6CELjR
0nieZut3lpwpNWTRugLo1IH99LmxLBEdsMCgfoJl1GQmS0mVQCT7w/jV9x2bD8PHs1xLLCXyERtJ
5UWoY3wbviK3zSVQcfXiOljLdeNUqvhQJifuCVI3RNwzGFmuHNMNltsruo4lqGgFsOHysYNNQP0O
7lsMmShW3LopIFi5cfhj5SERXv7lYDlSCSpCC70n0SMlanYJ03S2leGGC7ne5MyKpxKyWE48/ONh
FZjQSZQX1ed/nmfkSlam3OcYSviQo3FIDUSNQNu/1wvVHbnW4akKM3b1n+TwAcMoSG4v8JZs87B1
PihyDgZR5rDw9Z/VlUbUqqAsJN/i5bRQDNKPHCa0NLKjh6DgilWslu1qYPMm1ek37Q/O2uG/BAe5
3ns9YbvqM+DEjQK/kXxrzvBnA1BX2FDZwIwGoyGeudbP6HMv971eNNM3iFGypRuYEAM3Ap5VvNzn
Or8VhxWTzhAy8uM8i01EGujz9F6TOxM0PCX7hAPz3Qc9YzPZ1NDKClgQ9/275pYfgJHW1/YFsVVs
Oq4L0S4Xs/TmxXmZvCoJgLv1SeuqvEM7D/shwDwQnBAqv3akmj9Al37gK8jBAwb+uKAV2c8EyCFz
Oe1lvZr6MSHLNV3tdDocY88yvFnxKOb4Dhms6B+lLP5tWFR7zECv2wCp8XtF80ijC0wdjA1/f2IU
fTADjxPI8/OLUGio3tDpvEyUbvgw4IqqwyFkYSDWBYsK7JQuNHfMlrwh6ftZCVS8QMdeZWzgqknJ
/o46cqwweMnMywga06SExNKijIoHVCV7mYgWAPmbh1wHvG22kfa5qLJ5OFl7aVuga5Z/OHPmB6P1
BH910fj2JKtB1FmGNGzckglzq1Z9kNo02cBmbS9vo9VywoIjKHA3nWacK4zsjNV9QniE+eCWoecW
VnhBI4nESJoOIJlA08zxtPYsiNSlutmf4b/vWdFaSvLgbR27u+3zg+9A9vrYAE2HEZ6bm9ysUCnE
tC7rLxuMV9HZWB0o6knKPWPiLDcJaeTl8u3vm8gxwf0+pEvU4mF8UbBDbN6K3luGEAJErUomDq9p
6o7bPIBTOGfKMtBAYC7SwncpT0FQVGBvULi9MlvykFMRChnTO25NYthyDQ8424sdL3Eelr99ri0Q
MR7QdXlHlTOdkxIIdMcKUtqRMpikN6HUv6zr1B/N5CK3Zk272qD77VE4fqJ/Uz9JMABRfIVjKDVR
f9EeYvPfXrij5NHZlgux/xKhVBKJgRN5uGr2RmvQOeu6Wle603clGq/mBjopGGFLJWDbX9r2UOds
N2wh1por5rIqKhN0aSmKtb7CuiOqKA7B/ZNZ/CRgcQg2ZoUhHSPuxUCxb57iXRHojh992elELDEJ
SALuGE66GL9/UCNWzK2w+egFXpwZmpptr8fhjMFTz8w5UP8apMhPR5mnCeY4WJyttivQWgZ4fbMc
fcvnlP8oeBQjhsZqjrLAlJ02OUu8RPufyfF4JgMCjg0v4QcmHpOzPxqrVTTANTsqagK24w7P7Wnq
gDDo558bwgqhb4HgXlFGSOl4c2mwb2Q7vD340VYsqub3TsfeDlVTOb+3zaEJoVc3GVmuy2Cfit6e
grqE9wiSxe6ZkntDW/+I2J6eVcSR5XirF2EB2iK1i+4BSQPzgCWPm/z+WG7BzakHqYoANE7AwCbU
JDGrv/iZZbpxi1vwaQeVeV2QMTOPY/geDWURqYVM0EN6JGfihE4li+J9GRTo+Gm4mbt6UHC/A6Nh
EAE1O4DheiCUsllyvRXaFOgpsfw4iuXUNWn8ARfnzjwd+W5B8M5pCtmhpeT7M+ng3rpUSeQRdjnU
YP3qhXS5LSFFLAWbozB/57ap9hXbbb7k5OflMPkNm8scIJvHHuv1OGXtN8ANBovPTphhE7vA+fOI
FJxt2DAf4dM44Fx6P0/BHpkMbAVlYyKWJB2VVOxzqpbLtUT5hqhulR6t162Wvuz7m1+70GimR3gx
RXDEupQJCriYb5dqh8UTe3LT30J7LvFavhXV6Igu8VCeblXVmctVH2c9OtZfec0OQCc+6wG50LtR
YdCdXFZ1Hkk/AytcjIE5hFX6qVQcFaFVICJ5+bgdJVdBJSWj8TXp5nfVeFlktM5xezMs2rqmZtrM
92vw5xSOwEKhAeQdXVrsk7TClye7TLgxK5Y/UHBM7cO7W5FojOO8gMC4tF1y8NZPgKPYkgRs9nrm
2GLF35m95u0bXncq9Tdj0JW5c+YJzFm3JeAENaqTUoduuXQyXkBc+GWnaBp/zq+rrVgm9GWuTWvs
+7kPFjDcF5kCnwz2I4v9lxfjlzhgagTY5ilqUabF82+myJesaOq0sNzqpgTrHvCwpigWUVmt7gFD
SDsZ1VhbweGlfhcR+JZ04Rv6JuGnijL0+RsG8Uim4pILmStFzPSDhKiGxAL81YEQKqo1c2UaolJb
kswqKg3dxbi/HAM0nK98KnEzlgEEXwMr+jB/ycX73F/tY9XPpXnNL06CGJbVXP23FjFDKQ5AsSfC
STFIfNqBzNQpCkEi6FXtYGDp+AGXG0mnS0zCFPOHjFrvrk47WvAhAKZo4NxG3Y6hnzjUKBNcixkp
MNUU1XR1aKeRBR1CSfg6Nf9jAPnqJmveixNvS43bytaw9KqKcHksjjWMxVfiQAByq+CipJ3svHMh
HvSCma6tCD//+6wzkxQk9gJtyj6hF4Y0WjN+ZlS5+i1IB6lOfjamA63OdcHrzGo6Gw/pAzw9g7fp
GGG7mhTpUuResKMJQSiqueJt6oBfnFGz9cULEbH2DBhX7dHvaB6oPS3HSzeco9SRrXQXLpLKir7t
0y0Wf6izQ8oMBxsK7j1gxrRPaX2OXpLfGr5dCMIWTSrZvzscy3tkWhQUF1OOqnyBByjD3p0TR+f0
JdI+yzzTzzwCaIlwwwDIPne+SNLT4vQQ/QrdlcTS9GSWjP3N9Vx5YVrnalpUrHMuZIQCWpPi0wj4
bNhAYSo1WNzFhbus9g4MVciWEtCagI8iekNfhFP9ICOy+eypQK0bqKzPkMbX60mIYwQODOiKme3F
BRfay8qZmxNlNaSqihRR9mP9tSou06FOxozKMwNTzJ4ZQvbhikuHVx5VlBePYJPQvJS5/uccHPrP
6tTKXkIjRQZM1jZoBnhLTIpEqp5IW8+De0361vbYdR1bsNV2NMu+qQvBWiDrPKTOiJdmyeB1uoTr
6UVuzBsWrvx1bQkkQ2FOo29vvHC3P5wvroVdoGbwojIAB7rocb2uZTw3JybNVS4xg4TgBfXIQSLz
uF5noYIQfWmEFZiRboCfDq52Djm+hQiyXnV4TQ0N9Fo+9+ftx5swimg0jJbVj6PIFzrb4qgBPs+o
jPqPVdNrgzWmOL6w1ur0HgZTFKAjEWQi4dwiS2FpApXrTPSJ8dK4pBISbj3ymW20yMrM7TCtxIgQ
hG83w7gy/nmiACfFH3eCo5jVAgIKFPXAgh6Tt+XQdUhKHuFTA0QNl4npK1Pka9NSslMBOspOty91
6+74c1YtAkYXdaWW4mQPUl9FyM5Wps5vC62LREUv5U5DN3/C9At3JCSa0yh63OJLo1t6IHb+EsPG
UW7g35bVlNfneNeP0Wj2+twE7Fo+TsI6yaQrWE5Ua7WcAg/sFheC/qMGkEB26bdnFDKrMF+25G6j
pv6xsZWz5D+JHFhYAUzwIRk6Tjo+F5W21IX+P2YMAXuFmRVf+UcI9Uxl66Y2xBwQEXID5vFbTwc+
KfyLg8DJz0GRFOrJp+4AMCw6+/YyNroFg1lBwOij4LdeJjn8bLxG2ppl4C0U3vcY9DmjB0jPAKyU
nyUmlhLKZCvrB2wUYrSa6Fk/6aJdE5OkDnfvAjp+jPNMr65mAbdISnXMh/oWmxpDRJtknYmK9jHT
AI0xZHoixHw2gdpfLwTehdS60G945oNr/g3g/CMpSuLHoE6XE3gjsWTzyblrLQOg8u8mhbNVvDKj
lX3tVTPKkWpQTjodt2hZA+ZdLoTp9KojGq7xhedVjD70z8geZbgP+35sEUbo9UbF6L6url9KFWXx
OH/m2PoJ2ADwX4AnizYOLJxsKDznXL8WK9A9srnRemChbn5gfIv7B7ypbNKP7lYW1Hljlhf44xq+
i0DvJRbqBRzUnuvYnBatJ7gbWkqS6Vei/SVkiJY3ZzPzrXstqstnaHdY1q4ZF02KzZGhLDi9ibW9
WrrhEZnZHrsybL0+LGzhdvzvKBp+ABCziDioluJuZlD7RsfWY5attF1fBacMIP4yv8zF9oSxT/cm
SNtfQeH3pJTJ6Up2zwCP+kgQCvVG2Y5vb5w6GYjuFB1S6DOtYZeawhE0KARtzgPNsajGCkcPmddF
zBAL+xmTOuNXUeb5vj71u/GkjmRZPPWdw+HG9P0GuqPRkOneSpbnXJclnxwRd+JO5rXIW3O8ibQ3
kN7ORyzwWjDTeaW1qybqFteObTlrJVvLatyA5tPZ26ZaSziyZnEEZde/r+epwjKvJ9asv6RUEE4u
fR3kfAyYo+JVfSl9vX70d+Pp4slZz2Rl93Qs5gl1CeHdHfC82ftGmeDA5SFHps/hThoKZ55i0Qpn
xOH78kCfOgIvuBCH1Go+RRerxEZcewJwXm0ZQtZvOcyAgglUOMu+kVuJ3xxGPUflQHLnHQQBPdZ7
5T7abfy/8cl1r3DW1Ou5/p6BML3R1Hm2gUE6byOEqGC/p7ELhm2HlXjwZo+x8Ipz4cxCCN7BMRHi
02iF0kQDdCgBjKqh+0W0fmkTImXcjKj6BjB6hzk7BP6xDNi3VzFQ/MCitryIZ3hMJ4Vdhq4HiM7h
IjSRp5AlYuMIMcO6MKaJUvzGqDfx0L8ElBB7mxruyc3oV5//IDJSVy+7RYlZYWx1KJ8DuPxjbw6d
ROAsEMYnDVzafGXM26ihDloejfpFnmIwNFWHQKLnwdtyndpDtWBxggjqh+3q1D9SsxFONOC3HjqN
Us+EQO16jQgKNQTcqKNyRllY4j8PAJz8JINhJHSXUFuL/wci4ma+FBZXcjttChK+GvFcFy1siknZ
cVQ8MSo9Z3ovN81PC12fGvox9kEvslX4SbtbZATQjEz3hlz59dEjUFeWtf39mOE7cKqtra20/6of
Zm1Hgu1EnRmEIhU5oaLVjx7O/FFUydIg7jL/LiCAN8WmhW1DCv+SQ0vz73x3JDgtacDOFpq2xhwt
XAvwSSzEilnJi8i6nfkSenUH6ianW/JVt0XwXbtdYIaddRi2gWCmNJp7p/MDisafzbjQ5ficRWo0
/aLC/Rx9lkKEtRPpcWe0ULyTaltb6qphd3Ka/FW+amGjwCgtpUjp7pKFzRAeu424AUQuEAl2JJbs
Xw4HwqTD5wANeLllDcebhGWNVqXInnRBewJ4dbv+pnn3No2X9ew5qQd312/r/a6DJQyrPK3Kcabe
tBuXlDihToe+OdLjTRT+fEvzRcSeuCm1EsvtcRNXoN/taJ7ZrjyjYLwCf0T1W3kPV/inuiFFviyT
lT9BZeT7E/jNDQXcSB6A2DuvF9V6Pkh7o7lMcavSF3dPenZcV4UiJbdRlJbJwzERjtSZy4hbgEvR
Bu7cKvHiTB+83qLIMd5gqux9sZkD55ymq69dmpVoADR8Jh/Ff6pf7xkuUoYPl/ZSe6rfO4X3Nwx6
LjN9enuaV4tibDxff3IF0YArueHusjN3DRjwZ/xoKREX/2AtG3bTKWWD/nO9oadG1zNdpXQiC/6T
LW6XTi8DUbDtq5yXSPB0KK6a79i6rMAy46GL8D+dbkNO6/yeuMJIl9S1793oA3VBsEq2VVH3ebj4
9uCkmC+NbXqiED0XOgWegNBUKWT5TXPI2Kn94OoGs1ic23A/rmBkPoFIIEr+DwNydyu+h5C5ejRd
lZBXESSTLDFhjjqSwkPCAUi5+JAB8dc+S0s2lAIS17iv+u4rH9H8+H7koErgXylZVbcux0cENHfy
ts8LpmHu4NmtTsR+jE6L3cPm6dVfKzdTNaK/XKI7w1JCoRj2u2drWxCi9MpaU20+J6vYO/+dvtXK
tlo+1NeUWkQHsbqn3AcOn36RlkbROhVdSq7t10F5TdCujfBUkk0A9ipnr4JpIAxHlJttE3FslJhH
blr+EaB0lzMnu6DZx88YHHzLiFk5fOb1xLDk0E1F972ydv8JsDCEhCaJXQ9fWF0bb3Y7QVf+ZSUf
d3/IyWzxJivNWlCxnFCR82fljXEuJq9t3foYLPGTk/sXwij46A9jak8TM3A1tJ1nvBIA1fLfZiP4
40bo0u3zsPzOgNh8q+X1ysKmAQkiwz/Hh9BadAVnTCD8imiLyEMpEnvFsHQ6wka3pKS4enhdcwz+
cbwRFyT2qu2EV6GxD5AjnmJcUoWr0Krgvu1XnnlpL8LtD7UL4cBj/6ukkYxOA2fnP9Aelpwpope8
y1DABl8jgJltpEesU17B1mBn3fyR+Gj7xE871fOvEvgaHaka2rpRRA6Rz8gRcy7QdVhEgUbLPdC4
0jMXOJt9HTpBXKwR+I9aYGt2/dbD8dTFzn3ZDPMBq9qKt2RDTY3kKti+KZ8iOQJJSTdDrT/wP0Vz
8Spnr2e3Bci6/tl0cVkx3hPVvteETNZAcqprC+PZlWL1pnQ8ek/yV1gTyS76+SFq7qwukrzWmkil
n/a81p9C5t+U0i9lBUif/dlNBh9o7BSpTrj/D2COHCnkCeDwIOQkbcgLqhuKbQqkXINSEUh5Omvw
ywGYApTQ9bUIf6nUnFaZ316bJ1ViGMqyxGlvHNPXy6/vj4IfWSkP6dlT+8ciOTc3t4wEnl/p9MzH
5AzFRJi3zsTgg1jxAq78ad97igrJ58ihv5yz1uhbL1ppjzrYAFdtFLwE9OKZOSIa9NyeFISuQUYM
v+XRRzfkgWvTWCLwb9PYFt773au7wLCo4gA/k8GafUe37ToRUkjLv14hBDv68IcFd1ta5jHVRdkL
b5vP5Vd/6vGWyH/zUPXYlH+0MGmrc4Oy4UxTA89C0rskpCj1flFHi7Yp2NcmacmGK7PnJjfgloHU
GLNomWUXKdsdYRrFLlhkeoUe1O//147bIomuO7oto7TvOZVeWVIS7wzjRLNylr8uxvNlee37+b0m
X52C9eyw/Gx4Efg/S7Z3pPT1W6SE4tAMKK+xTUBWZOwmBjaYrQxckXrXW9spzzrjs7KsDPtZHfou
yHzu1OAhRT9Sb9qp4b7e2t7a+mPyovxUSfc4H7uA+L4Jgw0VrFBcxe7m2V3rPQaZq1wBUBLoADam
LAG+dycJRn83ZdEseaxKYS04QoUzIV4B+yxP5y25QSex/yD1xNTnuPcoRXZeaJospg4kaFVctzvd
/M2t1AiCmEuhPnc1ho8I/F8l7FRBRNh5OhVRRZfBOx0jJt/JSm+3sXc9Eih7QAch6N48XqO03E05
zbli21GUVhT//CDhTRwOlFKmn82eRApP4TWlSuKva86rXkbO36IQHLDrsHTMRXHjnPIk7una7T2b
SJNzJEtr03pMCyUGngSVKPJ1qdKj7b+Ert3dGv1/eSLLGP2ewK6CEdy8e9UfNxLkLbtcDZ7htcEW
cYk0pfoffPzyZBrzjAmzPUgQPDT8gr6kwJtN7Ar06X+KFCN3w704s1MtWHA+wnij8DAXZLjUUQJz
hTTdJaKwwLB3ln/k6qvrzGZq9PcGaFLx7S2rQQxgwsEZf9B1CIefdAUBvyotLhK5B6MMqa5tCAWI
KZgbmqJi4I3Pb060nE8nXZ6ln4SN/ohO+7ZOtztJ4ttf7pdKwv4VDmayPXjj2C1gGhnYuqQaqWO8
krwI5phU172yPp06T00lFwhmpxRdKot0S8m6GcNJyItCv5vXBbVXR5e74H+yacDpfuMVmNcHWVwT
iOVdNkj5IY/8+msUu9Zq07/uAxpSeS8irVLwKQrwRpIhfjMp4+/0x3/ghR72GapCVF/zQ7mL3o87
HQ0Mi4VU8JlYy/pdLqo4Td57QUwFBM2ghuwHZceb8zSyUB3V4VTAKZM9TaORA01j9J3XIWvwtJP7
HegvPGqEKoO+TQJY4HyI201TTdHi0rfBsKqfhfsa27Jmp0VIansD2z19mq5Opepu9gF/1ggRw1do
+F0OMPlHhE515IPjnS/TzKGa0+eL7No0jhYqX9Qdq4k+smhTGwM617lD0kiyK0InVLXUAxuI1vVh
XsqYHYozVH6V0+VjCv/Bu8QhKubp5xeICq/BPdYbB1xgtI0PX4Utfq3vRmvAb7OssL7R3SUJhtuc
F9WPthDEIAzmQ+X4JuBiM+NIedJJHks6wMq6W3fSc/qEfmPZiY82XzHaEkRAptGRonTUB6jxZXes
prAgnn3lIQkhjsEXAjis2InkjA/hfnGHgrQIFcOR5X7JG2tuRyrE7xIp6JYLnEzi49S7oJQ3s9lP
2iWUB1ijeGsWAvhPwXJ57lbbI/1y2K0MC1Bxs034/lBQdcmD8Qyv9EvHhQ2l3549/0K6cuKYBzLn
oaJLSxISfOtXnUsHTUNw3lqR+I3qlqtjP01totiqYFv6uqlt/SU8VwPDNU11Mr8DxCCD2AhsZ+D5
s4kvD1HrU4mV9OuSFs60D8D6sjsGuVLDyEIGwV3Hbv1y+NiJ1IIVSPwUvimi6S6oHcauPuS1la2y
vJmMUBkPoZ39jq5lCI6OXjU1pJl4tYyVhAmc0Fk3t9K/UKeuvlOkSAIe/2YrtyBIPxWPnHTbBHrW
4rcceco+zp+XpNQqfS8NAclXw/s9EdkIXV2ds2Fi9uWQUji79Iinx8Qkin5jkI/lXqsmmjcPO1Mc
t0doW2GovA7d6+oE3MVKYu3AkjpOcMPihtVNb2bXxdWIOaEwv6SoHFrB6UYSs2xTKqgwXhoVSMt1
ibOw97pR+vanhTP3YfX4+yu0XME7BQmIwJ8lF8HmI+2FIjy2pizVLbteOg4DQOGjCjCaUwgxf6sZ
cx9wiOhNAgOA2WMQoHKizqntsZ5CZiTHAEH4EAtqBRmNsTK6VHKN7wOTsw8vJXvSDuVTCnZTkDof
XPJ984ZfIgSdlRVrBbkoD3ztrq+9IH5S+AEO9CKxYiYPhRpBZ/zpLvmdfQH5dUX01xt3yEdGVjPL
4wJgaXQQqqpjV4JD1a2o7BxEOOi97hLe6bnjHP7fm46+UU++L12004M9f7BiZBoQ4VGeIOBqyr6E
9P2PV4f+ocU6prxvxUXcJP6FBpwYemQ7ME9k9gux4jHBSBFf20Cm9cYg88eaPtZA57svFwLtNSEE
Ogy8JQQQxXso0jMk+mDr4aRk4sKS/HXEfw34Mdwljur2DPJJ08KEKsOffz0W/ym3gWJMPRP3l4dO
L8sCuyz95fMebt2VXDRdxkXVY98+k0Z2rALxs94x8CYJWynwrRh0K0Jny+/VxZvHxoLhT8YBX1Me
q3XEAQ3bUoDSMDg9vIS4tzHlOBOI9OhdhvwL5YstE18jhcnSzt6qvNRdCEzoySs52WlfNDRQzWWq
NE4MuOFTKHpA8ClEenfq/XqC1aDMuYdSu6yDBtf9z1wS7lhCbvw58uvNZjbApJwLC7GFw8AHAcrE
hO5Ak5qrzra3UAGZ0IJF8XpwM+QjyHRczocSPXRNS3ky6Fx86Pz3WzFlera8/coMpsQLWnijtL4+
G7pPQC58jHe7UPpYzYhvs4KnYJU/z9Mo1Vt93HKiMxoolznL/I+BW9FTXxSTnGQNyEn0dq2IDYOB
bf7FFry5qAd4vfvirV/p+Faaj+kE8Q8DAQzzhv2EVbZxNhxqthW/J2y4AuPwle97VtLtUle+8sY2
UY3hmN0AUJjFiybZtv939GkCvX7U3uM1fErEBG1z8/MzjfR1BBM3u0PY08nnwQpQ1RFRt6KevI+a
YuAzmvNp0OhDOgp9wqQqsxZedlOyZiQRvV+40Cu4bAEnFVQ/wseemncOjUBFL1yKo5oQTaD6vLCX
SSaLY3F5GX1LJxXR1svCyLdqdJPeneXxOF+Bz6fZJgi9eMjwtX5HBRFz9cgnOnBdJQaNc4pb7es4
9qV/VI4X2dkaQW2JUn0+NcOYGn94e+auQcXWV3ao7mKmWmRE6znfYPVgLk4ndoOLavjPUDUpUWcl
hELNHqqtFYBZtLGJyqEniBKTI8qqVHswloGXB+ohVAf+5sKCpoAMJAPLeqwuTqdIRA+BaL95DUeA
3BHKwhWwy7y0CRrpgMmFermRz7OYeiEhPWSihaNP3IdtpuFoXhfPGMWLs3g58RbZsD7EK1ba4rKv
o+riLfyI8kQ5x1pv822Q2ck2wpFx0r9T6KfJA8Z4j3BwLLYfDa60XNq21UOTNh7vo6AwKC+tlPnJ
JJ/yEC3vEsOzkYRBtdcmfECtHjrgvMwMfhBqGASWNLQ/juLb6phwJeM6moWQi4Iw/C5TXSnhF4Da
KmXWHRGhJjavsbUAToIU0k1IvJAv89++VyGRd5kF1KVHCa8dHitXa1B7ilzLli1ChrdbewKTSIWT
WBmI66QI1M9xPGUfPEU/pYCUPF4rLU6NcMynCho3LTtw21/B0ztps9FqZDDotYtzKCtxGz1AL0YG
Kgvjq6ojhuUXcAtrKzka+wEHgrMLijmq9mGlPBmyIrDOjRVUzIQlXJP/tUHLeuxDtYxHcWg8HNOS
dY0lyf9xW9EFrSKsLZgs6GfVHNzBR+U10Oxoc51B5twOM5095a4KabXjlkqqT4twqYDEBh/tSkVf
n9D/ZJDM3lhmj5w8CZjItwvOQNtHn8eYOhheWmeUCB2rt8V/vwBj+wyrUlXsRrjd13VGE8liGo1L
ij0c5A/AEG7dGZFWYohkX//NOnuDQHDWstNet1GG/Ky7FmWWzOMl3cqosjRkWF23HCEcP/P4AZQ+
1MiBx8/jK5r+rDiB8yWoZ1TUtvV7fkhqeYLrTeDU0gOR2IA/78SCkYpkaVvHS4r3hkdmloDW20vE
Ii4HQaaso8iPPUs80+88HAEd0pyHnb5+5oT+RtMG6dTxkqpgxWUp1CGOp/6mloqr/qCqxhNnOQ2h
2uvgjmUXOgoNPBbInGZzJbyMjYy9ic4ZKdoapTTXKlcQI7ltKDebQAxZGIE3cusplWZB1evYvKPJ
CVhz4yDbL7rc+CuJlbl3qEO7vBS8tNQs1cFGPbEFV1Wi65cZ+CHVzt1IRI81BwlS7DhuyqMtFK2K
dRjA1xBg3ngz+av/YV1O1WPdXtR3tzgG9WJ7szNOPWaKNpC1nVnEEjVAEwWL14mQ5KONJENbdgAl
992ZqjFWY7yJ2xyIbsYU2Ta3oRNNIjf+RUhO8x7Z2d9w83UeZ4OJbyk+HcYrZDLsSneuZ1A396xn
IGgPrXmQ1/FP1pBxh+QEmUdnyF7ThFl/zScDOWujGBGKUSzQ1nxr7BTysqiqDaCVGS8bTJwEYvHH
UApTOk6eJ8CYCZ/7n/HRPpGT0abtfQ6rPGq8wKrsrTxYNBdVK6qfV+gqH0gW+n7zEjHjtnltZtul
kroscqyqhOPaTpSyarTPAjo5tX99rZ9Da+tFVmwGfLg8/dOBjRNfj8xo5qehQOia/QRXB5pVdHsW
fPWMp/NXC+6PheMjLX8A5yho5UK/B5X1QvbJVNAM+40OHYLAN8BD6lFWKmPYcGfYHdfAaWadmyOD
qQa/tsfi6qgRJdc0VxI9cmrXkSQwzy0Lw+0YNldqADz9IOpSBHsqwcelh+0ws5jhe/flvxCKBtOY
vZsJ6Vt8c+Duu3BTJejd74uQAKHO9X/k3sXxCgT7q2/0rslwGg1CIK9M+tcq92bFkJ6HtRFHGdRO
84V/KNM4z8JGcFC6gsok9xLhPrIQaJqYTGS4LabTPUnG/0ECBAX003+tIxehUvd44NoYD7WJowIb
Lvb3bp3I7nwdNiB44OpoR8rkjgYre9qdPVzt85fnpOdfo1wHKuS19DGVNfCb6QOiUEdNGyoEyERY
+2p+42StTtW16AyPhQv57pcvFR97rLB/B0YuNW4KeGqYmBrYo5OQLMxrdlbjaObK03Oogeq4yyT3
csszXFJBQ261M1/ctx6pQyylND71+rr+yn0ODYhAmp3gziCBtvcpOFbjYtqBP7vmlvmJ67+we0Iu
ZuwYtVtk69+feBbicp62x17CdxIE1G4vu93RMHR2eF7pS5V4P0fgSWgg+I3ZqiLloC8zY8DaX8Kv
PApar0vZzLoULkjgn7e4y3Rh2GJl5OuL8Tmu78drRg4gpjvNw7lyuyGA0C3LxekX86Bcm/txH0Yt
pzfisYacyUcgy7HRuDyjx5eBZQupbBvK4/jjBX8k3zUsjnDHw6+fsAPZUvofC1PnE9jOQtCRTdVp
5zZjgkJRPX48zN0GKnLJryxKdmaeXZEHyExu7JehdIkkY1UzsXsyK+ZTEZFeLd8FM6SvY27jIrBB
h8T5/d7mjD3QNgwm/v8i0cLPdKH2dZGDtHpy23wF1Sguvnn+bGimnUSMKi+ZgAMfZbQqPnTAXkk8
5mWK83ACpmgfOQr+KqRzxcI9F0OjPD80iU7xW1iP+wrZXNSZgzjJff0AKskY5/oU3h3m7D/hDyFE
QKSjw+O4ODFkXkWIEEb47MaalC1INsssV3NrYdZ0Zojs+FmNnakHjoRltMi8gpmJgMBBDA4AY584
a0Bi9VObaCVXx9AqEy8bzCOLRYTlNZ2Xj+54pK1QrSceD6fsD9oTR+b5GQXHDcw+ZLCKlfz2PcQn
zHA0HrUeUXpM73kO7OMhlXFyljgGr6/QjQnV5YQEy6UAj9PSrF/zzIc+7WQWDg2p0ZShxfQInodJ
0n9BdfoXGGf/rtj/ihfEpzeqD5M72FngnH9WMO93xB4TLnHyVUczDMnJ8AMHO1DjQ/cVLCx4kbZJ
8CJEQkRyeWDigRoVBIv8DAbedf32t6oQmqH0LSlKHIIdTBruDYlO4U4ayATocKHi4LblLtq5+sfD
7rLxp9EM60PKei5bvz/dFuF4dP3ZlrX6wjbQ7qBunhOad7mIbbIeVqRHXyxcd/4AJ+QaSh6Kh5k2
zyYIXkL+KXTzifJ8RuTLYAOsPGBvu60Rxsf7y3Ph0bZ5+OYJ6Ba8KJucyPsmyDhq38ISfcMsETJv
s3ZEnYFsvbDTromw3pGJVBo1d+RSOfDBGHL44lHP81H2k3eT4oUph5CozrOOZEuSrCSgpv1to6vS
gGhCnrlL2zv1KLrzyykVUDlwR+01c4i0b1s7Hg7UxspQtVWCOVVJ6bQNxt4Wlt+wNcQ5dNggswqE
zZ/VNK7ob3AATM4HePqtco2XFZnZJ8UncSeVHaFX2+IoDDwRDvQQKeyS9H7mGf06XdOfqtfCxcx3
yt2fVhOV38izGazk/eeO1pPhrCldSUJrCXno7oIR8vIoabxyTLNFxFk6ZUJ4aWssC6pK5/fAcnhu
sVFXOCea+GhBnteVrQnKZD9Tx0KZJhI+V/8DQ3nH40PMRvLWTGJxWaJXRp0mX724/8ZTkb9YB21k
JJL8dbTMelcuJDLSrQOJAZKs9ByLTjOGQ4wJ9Juws+6B+uVAiUWT/jC4TOqktR5+tU1u9ns7b+xA
X/3GghbnEKZkikAAwzHm9QCuEPc8Rx9tj7xQQrUvvhody5fOvwaHST8wpbmEnUefTNUunWo1UXAq
yjQxWr41XlB8Jf1wZnELzAbFl5uGr//Op2+9GX1w+1kxXskfR0HEtSKhW3cPc2aTMGWqjpfFS85c
yFhDcWIKHlin8rF3gC2VjqcSqNSSLz7YmP9VqNMg+ilSHuxaQyJ3en3IBkec4D4GXbPgc8D5Gs+r
rSTZj+OBt7M+5PeCsVI9ISYlhg+8HXe6G1u6HsKw2l848ChIhxPMi/QmMDacZdqDvIHsAQYiPNB8
mHvmkM1M+6Pn4mfL7eUhl5r/YzvNB49MP8EZzuxIlgffjbaWIamwiF31V3Bv5xlyqJCdfOLgn1qC
+/mpmrzpbOvyhQXWKbPgMs6wRCo+N1hSUt193e9maQpVdXnc2yoAHMnWka0+h20LP3qsVsyuCAoa
yL5ayxYAeCxUU+EhjpBr8VcTO6iTYTeeW5P8Qldmqbxu0zutGMP18u1FwGCwnWJkRE12hJvyBIhx
SBBTJaCdk7X71FGBarIx3JKCsXBJlKh08TB/TwEoohawOMsDc2T4L5kUOIhBkpckxvlQ5wJTHIlq
/JtsQ2pSwT7mUpldY7WE3KgnEFzbTz2ivT85IXR+72fOE9Kg8OMj3HT0RrPupVl5f7SK9eYtueKo
11spyjR0SAGg1iOgpKPDH9aE6Is7j0DQhLfyk/t7+UIb5HhzdzDRxNP94HhYw2Ce8oBm8DYiDGmG
QXumbaRrDH2IXAPov7dMoS0vE4+gR0IYCjdhlpE265us3tCTsWSB3uk3wGTf/iJOaAERn2Y2cHW0
RVc9xCyIdncx9qXVW4ke0fFIbVKRHW9N9M7t2OVdRNKadvgf3Yo7IpY+Qxa8CZedF7ukMHovN4mE
yqUaesB3zysByUEex871hnU0OoDWy2x3FrEFwNAfQrDum6RiIH66Mc8w0TS7qjOckUGjy5P4licT
e2AArxoj2m9kQ1B7CRHgvVwaJ6m9MBA+jOlJ5RfxcPPlvTgYscT2Yuz9SIFtxybkNZwQCV3bnql0
l9T8YRTOwFMp4uFBxsI5GxAzb+bAssjaTYtBruMw6iGFjC10qaqqQC8v5HO4lKeKVeEtvUxaSLZl
dlFggv9rmJurt1rAVpViWJfO8u1tq7TqgmWLX3zOp/Epw9mvWtKKGdnvZoMlsVRpEtVn7cSwCzbB
i/eJTdTBBa6CZD0LXsbitXzKaFhjbsY690tAUt9nHXu34YghtjqDQBsWEOLeg13yRWZY7jiV09VN
ED1BSele7hht2Ldrzgt9MhMhwpp7HzYtb0PTdQ70FCCdcp9GEqe/rruOltuHstluEW80Ai+2tH4E
Yqu1jtPrY9n4YFTRWIH6DELuRwJazwpLmTQV+ttFy0vgb+oP4y8ypyfZTtBLaGK2Ze8EgkfJ56nv
uiwlOraSQBR39uMuvNZ8LUCNlkacz2wb/IgCk2JAJ/VwobBxq8yqHf6T1zKq9MtQrVrXikbOWPNd
xiynWdCwsNzQ79VDUqzaf4ZVmBVM5RCka4qSxTHFe/L9HoSwDlfs6bSf07cNzmfpjG4vZA0rAb8n
rj4OLcK9TH2eq+6FxsN/+e27Cxp7GiDCnZmY6t5d1Vk6woDUT/eOGGUYkXA643BQog/HN8eU77oW
0WqR4ZKe1q4uZT0UTqjMrfatxm7o+Kd+JoW+dsZej3xWo6xtI4nbQRxG0+JNlwo52OHapfxfQOOq
2cmDVHQjoroUwKKkxex1wOqGWo9Fwly99tJFqQ0E7UYtYAp6e2+3w3kKAH1baNjaA9nclZkuDTYl
++i+7N7Im3B19G9t8bQ0kzAbIpJ5AycySsCqYTuQzabfGA1X/ccrSZD0ch5zvM+W8Y4qmP5huKbr
JhsZDTltno7KW9WLg881UbRKOpO/ilaQIXEKg9X702qsDTQmqoQM2WvOj2CmbhypXZhfgVzXWHJ0
OKRkho01nh51fgWbGe1nLTxHhsLXHs/KKw1x0+pRoLiQyBvir1geoXpGV3Kka3feeUzmaqZnlK4k
MZp8KYIraRDN/jCe2u1yPkC96GDxm0FRUUkgXO/eiq/nLBvv0tOtVL+MfUeibG//f9QLRjAtvSCt
pQt1v3VV7kH6EVsvy40kBooCfj82yT/X9/LMvwYjTmV0EpMuM6a2bEtGAJQqYnoiiCjhvfbb+9qL
0cOvfo8KVtc2mEu182P19Qqd3INvZm7fZwuEnqTZGc10IGmg+bBR3QhGqlTBN62qJPJdkGiQ7irk
d0awHpOG9VVXo7BSkEV6KExNmC61Y3Xgyd65Wy5+CJdMTraw7YX/CaYbetcV2N3+2BKwH0+ra0ec
9ShlR1IjI4KicHkCXDUc3sjcKZ26OTd6h7GItqjtC3Vgmgl84AbDxix0GuBYoBmIJa5aA5gQCDnJ
MG0Tv3psTuXUlUbrNqp0cTE17/qW5yCR6wc7Ch+HA5H93SpIyAeaKwUjg0OulWhQ5AFu8FIDTyOr
iXvf/TZ97FlK2dMc/X1kzuIWJvbU6Vg3LuNRImv6QZRp0n30jvy6K9BQNubgxoc37QqM2DAfjyxN
voW899KWcMynuG73zuFtTr1t4Hud9ET/3tX2BMkJDe+C+Z0dunbLt9oF5uEJybRqMI8eFEcbVYho
UAYchxnONkZBJj9ErwiaawD5/WsAEWAX4FRCP+Jqye5zKdV54DKnkIIKr3gVeJCeaPg1jaHlqubx
Hcyh92proxWw9/pANLXGBrQwei1WIK7Nvhl+uIwxEMb33EXJbe6XSzAspLJCHfAD6P+pHI8/7gm3
QwbdklQIP8fuC5oAgSpGBe4uzT89GIDoZttrWb7itcu/gaNnzocZV+3WOsASjfzTOq4vV7PZgHVc
JvS7wlw2Fim5ff/E7/d0YsfReSe2PZuDzj7kotf74l1Poed/mU2wwyIAetN6gPGRetfVw9UOGlxE
e02eFK2IbdsJhD4SA4S6FdWaiyf0vYmXZtRr2kiQcQM5ZOxIOG6D+x0pyh+EaBrahit+pEIsYm6t
HKgXDe+KDn/PrTvFn7Wo9Ma24VEnMoXG7NHTzg42jZIUP15vo4GO77lgxo4+ygUQCMm03iZv6k/Y
Jw2W9pLvuYD9W90XxXfYBvQowjWx2RrIRV9IH1d6V5TsJSt6U4UDGzOXJxyu53iVLyO6rKUVPbDo
4fJyNNbSu8RvBWz2MLkYxa3h7KHqNnaHBpzhB5jZHx7O1enkf1Dd/pMu0u6Ja9hgH4+iYX1zq1Pb
gWSvgwZMv2p9slpiA1wRBlG5IpXVXehh4tBZOoUliSRu2iDHrEOnTLA1a1exG+zWsOnjOIRC+mFz
NCf5gjLuBy6yDxtQUTnsYQfMUGxyABV0cN6P9MjfS4cyX9AxGI9dSMAzya1BrCEeZwlEq/tzLqqJ
QiBC6Rf3ZXDv4KYS0mf1UxfmLRFEHbjW1Mov/1rhK6RwSIBahiJd/MjcszFNBgupjBcNAU4YiDVs
T1Miof3Vr6xMfVSvweV830+1n4bdgZd5uv7shpNbPUgKUP85fI5mCZuDPBzLq8nj6itINSvuzoTJ
Rztzq3pCSlO/d3gU0VG2z+dzuZ7s0WptDWc7qxlR/kvs+BzO871Wrc+rSB5GEEmpYCp85d9Wb/xi
PEYILcTkl1N5unSGnkS1HnaIWeZj4BBaM/8uTFnVtZwgdLobAThWtbran6AnnLzGoCbFVv1712Rv
GT3CKJWL3q4RXE7wo0MCGi6W8qZ3VmX84LRF6R0Hz0otrnkG7OeF/YnN4RQlKI/vdLD526EU1WV+
IOPiCeH0YfNOcAagOZT9t93VK4V/pbfTte7yY3E78BsCe2WE2y/o3eojNGBZfA5VC7xhskohMYXT
No/Uj/RLXN/ie8vUfNPn4gOozGcX1nshYRGbTWCnmWkagF+U+w9mwd+Cg5N1S5XPtoF0Cp+QidN8
6Nu1v4BxIWg+qDHWp5ZAPSwfGHx7ODSqhsP1Mg6QiZYuo2wNt0LebVqEUtBYTEdXHRG7OvmCoWEQ
0llRBkauV233cHWqtAdkSECBdcqUf6wEshfbsvaRhVFtk9iL6uEA+YXIwyqtGhvUEQR7X2Cn+tx6
Th1PMXAb2PNPofGuw0rZMeSoNvQXIxz2aNq7boyZDpGcUD35y4OQJkcoMlDqiZR31JCLWPXUKeY3
Eo6JGIJCOakuAPhCTX9IMI2jbn/rs0MJTcMyTNVgCbkXxA9EUeSDd85U6LObIJLQlR2OgDTKcQqf
Tf5QaAH0nVL8JSw2NUpYtPjpBmkXawicu/SKpIl/ZHI4D7RwLK/jgBIL8p6tK7PwICN/aPp2RX1P
yShziE8vPcuJj02GBvUM7bJ5nMIyQIvk7uE4Kv9UO+Eari3liJ9N/B3gbr9kHbUEN4tALK9rjZwJ
rusljPDWnxyA8yihtt+OIvcLSnwvDndNLGcfbuK11jm/FMHo4ThzHxgrlsdX1+mHIrQ9iCYr/kmr
P/lRfH0RqoSeVjzVCrQTTw2p6qQV/QsQY4cmpCJd+DHJZR2RE5t9mBfnpyyYmuyZZt6hnoB3NHNn
1rbGGvV9Tb7y+uqiFf+mr1IPyndNoAvZKRNWvlT2w2C7ch0UDkzfBHiVNtmtOUo6AoIz5tNjnXvS
PAT+R224Ii5IMvPPIJsVgv41fsScictByjfIPFTWNl8EtEOOuOSPWyrhhOxQJZDWDiFEyNOu0uct
zrYMTpBTyqHNEyGJg/5whi8hULI2aadQb7zxFZiaKT36zIlPjPoMEUZdhNyaQCP8VP36CMvf4B+Q
hK79J69QoVlBSDUJz+PdhlYBoXFN7Rg3TPvEI7JsksZqfpkdybSUwID6+RNBkPgS2YhvmjBOoiQE
tm4yGGGq01PrCserhi28SctjQL5qjqodn+1KtSdUfKgaW3iAT3O/8lsWq/E0ZAXrGwYCoC3xab8Z
x8i4aqaSr1Xr6vwPJ/yNyW5n14TWCMep/4XvO46S8C067ZPO32JWQwzGVSjjp/Gmk7yfy7lIDYQB
bqjhGaeDT0N0SszS+9Q1UKZ+QN6yYac9HqeEXYKBh/TWazxFCBSENbHnnpeWsW7MVWSGy/uUjHgx
EBJ0upH7SyM56ZHqr4zEoSdDZSS1qIM9sWGFaC4tmPd7BdFPJOoeJEbAszhNTxhpESoMRDonbTT+
PeGWW6r0fNtpSI7VWjjqKP10f7k/XQq6aOqT3RcBNQLUDsgeUokcJQwMNIPPIduI3oN7p0OENb9w
4jgLKHYpG52RsCIkG9BxIVcu+Ou0lMbevVX+NMz2rpcvNBNz349fUL5ZcIzlfJAiXaJ8t8eBHSh1
juUUoJLZMb5vTuRIvLQAv0KVjedLoAKvCGMydR8I6D+4mYdXZMfcegjUkQbA/UaOhk+pFmq/c4Ud
yPJnE/VHFK8s6iOVE/NrHbts1xJM66c3TSvSORk9380tWJxnC3dY4BZVQGYOer1AkalfROIJ1XJd
LbE18553bgGTRazhoZjxyVJ8de7gcMAlh7fK9u5mlLju0ZRsKglratdKfxSnbZKHvAQs4uaIuyJ4
786QSr+OflbRUJ0qOgajdYOqjilMm22KSvnf0S7jAc69mfc4DUaP+gOXJY1GH4D8vIZ40cMHYQAG
tYTL2skiuP9urenc+0+Q7Or7rabELvMdiu2sFxSmjazdSBgvVRUsKMIZOSQ6HcB9hJKfBLWt77M3
VIzV3bmM1/CnvWM4pZl0n1M7gPx052mwHZneWHMHq2wpqVL6uYcUoOcPQM3X3Kwh7PsLwXjEGQWz
oeW4pgSqqM5Qi4T+RC+5vd5LF2cHID1PZMrNzuUOBrW//fJixTnj8HWGhcf8JB0tCVAy8UwN0Ozd
sDAxLxzAulwMluqlhhc0+w8MfpBgcsi3fJ47dAg6dv2SwjvXAgH11NbT1IChA2DU5ZawqSfQhDTe
4+zjo0vw2KSflSZ0DGF5DIgzK0OVxPXXDT1JOaItH4kDDFDiYEz8RDMpyE5zSu0yxHTz7kx0tyLv
smkL6/IOccHlCDPPCBXPdiKGxvEzXUUvsbsaq7Ja6ctmsHCwNF+vFq7TjahrNsDkV7+w/YrKhT5u
LrAuZzRJYOLC0h6bf/zRMolH+x0XEQfTJyoN+gGZClLKdmYlkTu9q91staOQkr5xY9QBJNNtEXl0
rvVvhRVcMrnTWYwZz1m2w2gUVZYq7xt8/CmuQy5j3dWDPCAFnvKEHOfN5IDVvNGJJMhUTY4Dy2wp
Cjn/jhK3hAiYFKvJ84kZoloX3t4gW2LTzCZOVHSvbm2AoTtNr2CvH3d3/SRCsHL4e67vsDUkILFI
BS6OQM2QbjQSx9ePySDwYa0qU0uY7yZ4sGJ3Q3ZZ2mxOsO7Q+EtEX/J6axrLsM9GAYw4GKfalTOY
JoRTmwVbG45BrSiOOnt76R1/qtshgb6U2093Rl40JO4AN+HgqE53w78EJlytoU+XWLX49pjz2kmd
ECcRtQ6G1w7lTO7Y8RnElol2T2x41iU2gJAuXUO+O5OY0rKUVBRJvp2IP6n7fO4mg0UBP/fDKa4S
SckdIYCwO1nn6qm+ZNApLTEhROolTdIXmyEsOESwYRGgl4HQvrmPWgGsFoD9uOSx93+VUDq9mmF7
RP9otzyQ5vy04eieAoCheUdaG7RZxpQf59Nu3q9ZYC67IAtbgj1HR3/fqw02gPlWOT13cax7ybhk
FuWh2YH+ENN4/HsM74GOnHpBnwaFKmJI8l3e9IMst0psfx6OYmXTGVfgpIlYAtipAq/FhXHQFBgl
EzBlHOWfY+UB32T0xNScHcELP7xlsMRxjC/qWsfsdnE1hP2KnV0zas2rSkD10R1siuDBmHiPM+9J
xzZ0NMNQNGTy0AXNArhVvDwo8RDFFWRA0rViHk4atael/lp/pWvA24mYY1vNEmvYuxkPrh4Ur1C+
Vo4S4SyPiZKtP1od4fMXv9uD+OL6tsuq8gOHzUzsIN/lDO1dpxFinpxTtIh6ViUeBdw8EKwsfpmP
zlEpaz/TaiUA+F2NMo10BOgdOKrzZ0uM6SxrUiDQGxqTqq4iNU5IMKcsl/En3seoV7+rDTC+gpyq
6XZ9WoEvq3s3ZHDzKle+HrfzNEJFaV+4Y7dhCUbdiTcstQAqhl3e2yC54nZBjLWtJduhMqr8q7ZM
NCewvf5aYGfrHUgr6Kg55/ZBN1oCKj+l57MbW7B9yHNgZMwboCTwtAGxEMERWtuQt75Snovbxwry
xLDXye30EfqTCdgCGQ3JO8LqK3rk6bBHjndC5T18RrfR478pqaOKgO9KYB7nnrx5NE1nR+H7cIFQ
MAStX3lXw4zjsa4u9PFGTom9YkfCtzPm35oNeHb57mj0p3aMU5T+FQX9jxtc90K1xHd4jumHo4qq
XOp32aEqj/AU/V6gMXT4J3okScOSih4wY7vKMYDkxWZc2oQvQTfqsPkLkD8XuzrENOxAjWYU7+O5
RcOIrwXhDVr7rzoyU/Ggd8vKEryCtxsWxRBa4rCD30frS7wh1PNx6zkJ29YAwKocMwH56d0ut+Kl
5tKDOTsMeERC/J2TtmtCB6Z4afqcnOod+jdrnnRHiCIfiQNDof0Ftq0SiHkXRDhvtWkVTK3XVw0u
dHvjnHA496Rd14OX0KAumnFSwKLQinDGospcBdNTnLFfwP+Utom+QUiQ7z2KDek65xsKeQiuVMRq
Sy3avtuB4NVSSOFeDWFTbz6c1ZfIKCVoAaKDLiZS6bKb2R41Im9YQNK19iup/IUeZM4qlzqzulpD
g2ZhgTor4hua/4M2L+Qgt2XatW5UakV9j0EgPmDp3IOtYESTB3cS5gRWSvGIh8T8BLBAGI3VXL78
6QRbHquhshM9NnRrwZ1DztVd6eQRtJN0CvJ5bL4TpLWc0rWOpKUvt19miNu+Oag68y3gTwUgwkw2
cwFtSuHPYkQlXK8aK1+I10aQgdbiF2jw/uFIYeWnkdtAYEU/GWT8dag7DFJ2Rxg6xU8/AKe6u7LU
48liXGdBmurSxhzRQVKQL5YsOM7hBOXFYQh4x3M1QviQLraJlbDxjfsj/+Hl0O7KuiaH4ZJ2/H7b
dssx8SxhqAU42X3F40w/m1UyNTplYGLeQ2ia6cbTKiBvZawNmC7Rua2m9xy3CqDkkGRzh8eodnfn
pTJIW0CTkSArMBEbsHQuPnGDP2bsIHIzFfWO5MfFZJZmVNO+CW+eI9MHmQTN1Qwqsm68lvkDL3DU
oEbC5zW4bj6YKw1BFHFxgBC1d/OjQ0wpPtaQvFwzXXrRKwqzcumN9OdAoCnJ+A2+fSvq6w2M4Thw
l3TvVcJmvg+SKzJbnSGHvb74j0krPThJK6OILWfUXsPNuAzdEUKQhxG3gUF0CN+mZb/wkD+T6ayO
k3V3NrXdeg0IRIBOjYOb3w4rUfmkIVnvnlC507f4XF+9CwMBkXl6SBLuNY1I+Z3Mszf7jbssTss/
6/yUecwCv6aTzn/VSh9pjhZdltKM2ZdmCpzJpgmdQvXMdW9fQfwHIMFUmkaGAw3vKDy+kUEOtCbP
gPA75h2wyP8kReV3s43wnAr8Fsh0VrqrxpAnSSMjzDx8QNcJFnMpfcDmajCqpiaX4YBvKQ3t5nAa
vLHqnywpx9TiKcDkapifE9VzvNE7XuS//T5gF1DIHz56YDu9freCg1Q1pVdF3Ic0oqK4Czrgjq4Y
S/JNc7NREhTbBiQRbJC50rAQN60pEnfb+DCd+V6E53tZtTLfMDNmYf/SDJ/kKuEecBJDjLyaxqAQ
FUeeQeRa4hgAKpaPcpPJJvsBNIJhaK1zEr/01XIrNZIU9+nCPguub5cu7X5rExQYYjCKPZg+j3cb
gQ8IiIxYDduD1R3hZKOKZ0OKt5cV2Rw/lyubCAhpKocSd4axVL4VOmeFQt88CFUtpWl6PqdGX8od
2HrmuK5ioBKtVcT76aUHgfnFlNGwRs0P
`protect end_protected
