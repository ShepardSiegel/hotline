`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
l/jxKdG4lNdaUs34oYw7fy/1c7SMmb29DNnEk9OL33t6XQviGfA8mRxPELlNvOl1xNQ8SqHKRD8w
3tOs4Zny5Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gsccJsgkLH48iAIimOi7DZ4db2Kx2TnH7vVYqgO6ysxS7760vAlM+k2TJj7+AZCRI4aPgWzEbabn
A4DJBAf7497byKRgadX5lxX+fYouxJWi9YYwS+IVXuDSKFNU8/HuwByVneaIRDhH/AJPIYZ+DjyM
Ssg54dR0iBs49RET9vk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ji7l6+rGox1+6UEt+OzEppnvyBwmWaDg6TrfNm8j4G+p0aGzbJys0d+lCO0DH4sp1Y7641cen8rI
EBfKL5dtt30oYCLLC+FswSLYrIkqNjpZteyFynvTwx0H59tEnPixFW5LhmTOf8n3Uv7KB6zAsLNi
0M6pur4GzR+QNkdiu396OwiWt9ovEdKJtZaP1ht01iilGZ6lKumSddgBlUokJBm1JgYNDEmrRCti
0jusS7gLUzXDO/xvPkS24Bw9+EiRztaThk5+AoekWpJLgVfxy31lU92O9i4MgZOBKvJx89BGtYQ8
4+OmIoAoRzk+c9OH2M3CB5Ah7SAunPzhgTTTpw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CLnorwQtoOfX9le5Ffl6XH/baIT7HjNrJL+VILKRlR+90ccZwymGnFn9LdKbob6H3uIzt39orSAe
uvfNdOuUNyZHWHIfQv2eldeWUlOZ1lUhv3qE78cIUfclm+F2hHceDeaFbaN0iOcC0OQLNNjk5qoO
lwmFbn054F242cxYUEI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S/XknA2jg4YGdTBPLocjrsjlZJeyh5BC1gu/y8bbj0+Lj/9WW7w6TEYR/u26BAycbmMnvn4g6Wrs
ahJkCXOcx9bEs0OhysnMZVAz5GOZM1c1BHDDZYUCJ6W6KadB+v99ZT2zDE3zcJ9HRP5QvNKEMMfl
F5bIIRWZE8E6gBib/eEuHe/eZMcndHYjmdl8+pfoolPO7cX9WSlr/PeexaJLx4RnN0hmc2xBydj+
pth4OsR3KEzamTe9CV+yvwrUPnxHC8A4fw5Zd+3fmlXb8+ud8LY2iloM2Y8LdYedYPR8MCkOG7nM
V0hGMEDdodHv8ZYW1Ow90AEtqeP0zUXFf/o5Xg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18240)
`protect data_block
NWs8BnxiszfIH4Nfihb9TzNgcBrgHJOr1Fl1oof94cMyOp3DCS7Uj5Hzy4qTkTjB8xSYBdoKGTdl
vZwTmeUGo60/BZDR1xF5cOr/1q0V/5QDaVpUxRCDoW7VGInu2ZRwQ1o8yh0kAwV4K7sSJLgAIAVN
RPLknBeJEV0QVaI3wga6u+lZNfvp472vFsIG+9fHcVtFutM3l4l2cQfoZLBf3cF/Zis3DFTv2dJR
30C03oxPIXFain8LbQ0Ma1gWwmhlAA1FtHZbKgrlsbuZYI+egKi/DYkPgALho7X/OhbM3ejcNVDD
/FYlRtnlnRaiit0BDhGbX5h9vV9UwrVNnhs3wvD9kp0EQPO8lFq1x461kGsLIOTb2MEyhwnyyCu0
PPBdvgiwaeuNZsD79UxGEj3FFhMQkjaW4AwNaSLgksWNkSd+CFAIiugFTgKLbkGsdNPu8DWwSKt4
UoIeOEHTQwCHQoAl4KO7b9kIOCXFbDZYB9ReIcZkArHAxbgCON5dvml+8oZ55tS4aHaNkHB35Seb
iqC51hI9oYMcPzyropQBHwqSJLADyjlzmRUcqnTj8lzwmyXmemLeooIGP5G0bhbr2OQ9KjTXY2WG
oiDfx6xUsEfnAtc88uho8xESaIvKiguHUirZfx0cLrW4tLxCjNwKHPtCWUWgVMRT/M4d/6LAy/rM
GkUwxeC+uXw5X48/qzWa3Tf7dWEdtS8RFvNi2j2vY+u7sWVejjrBqB5ZyKe65p1NCAebfsFFU9yD
42/SFrcPHi50KO2CpkqX1EVawUUZrittLXqHffsPmEKTJwyN/ok27t4WviZZQvWY5qluwdpHqUPZ
7AXMjswIgS2084GWp+k3llzr3Bxas54laee0ikpVkNoiGKLAtOlhSB/1MTaBq72i85ssGDVbbbu8
EkZfkx2Ds9OVYDWuXsfq7RQ/Zr2SvWsegzL0iezbJQwMw/CO5QXIGFCEcPPLHCOIyvKL1AK7sjZY
Mo8izLyUnC7kulzvit/pGM65ZtPMg3zNb0pxmJfHlc6X0pW/HfjQ1XbqtwdUy3ELCAa9bbBBAWKX
9t5ETgYXwqTcGpO9MySO8e7qBqJKwcaBv6tVAbHTLJaKGIwEyooaFgpmfCHd885aWk8As18DY/L/
HYRzQltB1COlkNPWe50laksA7RNCj5m7a1Efm4ZI22V/LFSHflojftquByqYgWBI2tvYJH4RLW78
aKkEDysv6xYCxnvN5CmP5I0JkO+TFLEVknxA3JSHqVK4UWZT4uFhhMONOz8liIx+SaBiXZiq+FcK
bROK7b+BwD/WgWzMbvw8oPdQUigViRfJGEdayzoUTbYwxcb0h37AdwzLZc1KXpAUrJVJ5vHSO233
lvSqIL4mwx6X4HzxM3bq5hz5vZkNaGZZLkT3GsFa3qdc2wu7XpuPDbVPYzjWSQlYGGujTD8iIkpm
z+XFH5+dgQDtHSIn14lioGzusZRRSK3ZjmD79tpZwB3ZDecD/VVK6vL1456ZKnoyWlxQ+qyf4qb9
WIr7snXaecv71nRuBv9+OMhzSSNNqJFkzh7HAwcYHBz6ulajBHEFObKnaJlF/2TIouc0SDgSANBP
lrWvOaDyb89CkgrG+zCj5UJKtzqituocUnuKUXoeOT/XF/IPrf1clw9xvc5ImjLM3+ME3WO93TxR
keVbSy9vdhKyyXWu8ZZLPqAowm2PmLdj5lKYvig+nz4ZQNtENVGw9VpdYZUYj721sTr+WEwOz+6n
6iCErlhtba0RkL078lpp09QX7Tqmf2jk3UycsuFZdkcIBiUFZfJhSrBZoBHVrlz3lOO+aByliw7V
yThKK4LLOZLKY5MAlu72eqVE5FBbqmJSylCgDawz1GBcJnajp2DOKW10YX/7Qik026LocvJl0VOA
SxnnaV96IPSymaF/lc8mUIri0XB8D/bXQ+jc1R4zUAPq+3+NRNFDu82hft/Z7CMp4jeFVTdurXxN
526Y+QGE+CQnkjrIpAPs35AJyzcY/EnKnREbVzSSs/UbJXJG0TYHVVO6UKR01xQ/6yYeckhkopyL
NbJNGM9dnSN2igsiG557tjrEMmw5TOeODccFeYJf5ioTRAYUpucnqM+fZRbHFlWnc2iT1YkwZQ5v
bZ3Xj3uJM+JPy96KZ4qPJmA11pkUMwDBxFW/4c7MMGqSHqYqvXgLzsAGhdkxfGtbSYaaX2tLAsEe
D9PyKO6fBevRtZVoI0bhIuFsniktdExwNucFq32IhcGoRvKhKvJTOvryzAmxA3N0xFtSPo+mYcfd
vRcb6s9vVbpMqm2sUJQRsMwSxscQTd5IQZpTVG/L+lXxMM2hvQRC2KpmsPo4qzjUUEeXpQeknCil
WRa0y0QyE5blKeuBa3/qcw4QmrZsuJCljWaWqltDIgZSP4woZip2r45rjG83ZpeGec/r4gFWH8TP
M5ADUR/sc1hFzPGQBZfjpfsEkw/q23OFevforbWPhyLQj14BFJ1jcKYvorle+pCExA+0B3jqAFBM
BB/7gm1Bv/d4fUyiso4shRVEh+3xDfR12axu0/1fFPBqcJHo3H3hgryyoGrQp4ZLWCW29fIESvU+
sD7goRzMbs4Uv/rAhdE7rOmitKDUGeg7I1E34MTiK12QQDuRkV+gl6tctK1WqGMVV5s0FfrN/ZPY
NQzIMzDo9q8wg4ud4qCZiSKScdtFBZGEKWujTgqzEdIH2M4TJEvx+SFhUpdnHS6xBHCWt/W8e4Lb
V3mcPG7iZmwKTMzIRDOQbEKz3RZVePaIV7sYVz3lj1fP/AC7ghAiqgW8UlbdzSWRCqYzQlB/sCjW
kFqSpD7iWL/LT3Mnl99O5x1jHaT8sKF4Oa7YXU05X7CMCVQdRWUi6ToBKzNTbdQRklyI1lm/SmhV
7jxGLn81rORh1ZE094QtRoF8FEz6MDuj3n/MTLX0P1naZhL2jKB2RYT7VyQzUuG3aBZonnoWNO25
Ge9DgWVkzp9C6WYW2Ky05WhgaOIgzpQ5z1crixB8MNhlXShSvO2ZI9beNTZVqGVJzow5F2MRuXvL
GJ3z2fHicjxn/rtCuqLOCvFp0YGbqjEnA+WFck/nKu9HNOpIcc11bmvyWuzltHFNYMZHSGWBdAXL
jdHfgdT8HKNawQmEn1rNVxcv/2xmUP4DqZL6A26kbk/mU8W/I6cNZiYVxUDNmoLj3jcCCgrnC53x
lju9i4IuMitnoIdE2WWus4Px2oRd5FCGoWtJpHG/S5/86V2azSZ1WzCfWj8QDMp6vHS4y6mKOVXI
I9UQkt3AuvHQqeavDDT06+zKrUwCDMUNvypHBNRKdbxBJit2pGtEU7rryf3xwk71KyQXuveeoNLB
J+6Vp5vSObrmOwooFivbmPCLlO5Hquq4wvnTrmZy2qw+3yjVdSNjmTFW6vK0MyPV2TrdAIkDvrll
Jvb2ORb8YC94TdZt457qAqKG5hztSG1MFMve4ur7RJi/1UPJbFfJnbHHiea30xEjQqmYKQYNgAbL
MLV+hzacaU7SX2bqGKFUCTgNV+Q8UNM4eOvcDmxCQoKXlcEeVvxe2jugdp6pmgzLi5BEkL0zqKSm
L833V16jhJ5g+iPDHzXdL95rRO8YMJLj+XZsdgT/fFwSOCGQuXSjDteezDp8fxMS8amQ9Y9078YI
qlRATNxUr949NphKdmx6ultt9ivCSvhA46KbzkxIbaQ044TqTZjfOTxPyxwT78FyOQq57bjR5wkh
80g+dBBam8szTq5BOLFeXKiyzsIKdkUdRBiezMGnXmQONI2ijYQOkic4gsMChH5DLDpEf/wanjq0
qieImvm6DMzsK2GDMgCg9rS7FGSxg3NYqAuji4uPXFPMNI9b2m4ykh4CccNjGvSswvPDppb3m9Iq
r59xV8VxJKlGZSlthlYYP91KPX7JDoe7/6Lhm3ltldYf5a7BShjQ1YvZR+Xb0selQIKeQt/AMBfO
x47yupa3jX0U8YEhF6cEVFi71F4zrObnR6Ti0NH/8pbAXzRdiTEB/gNVmqybNNYZK5LYG4Q/Fl09
9/ufJ9OKnMYyVm4ZtV0vrFX2VM36hYWE89pZ7anFc/Me6/U6EwNuNsNoQL5Ena78QqPYnzGjkCwZ
DJflBg+FMdBlw5Y0N85gs2nxs5xqEvLVuO0e6stTSAr9lPnHd+gwJ3Oje9u4w79vc6Ox7pi3hiem
D99eqafC3hOYHSOg5O0fapMA+hLTk7ICxelPnMhrgPxM02eHLjEuKUkAYScJ8qYBNIfyGOIwG2qz
B0i/lxlKTfcB9mTq12w76pCmYc6FMLeytdpfywN+A3ScrCL9TcfF5C1ZW22c12hrT8J7iT9FIPfW
Y8J9iak+eQxeMDZLDEYuqH5bM4sqPU0RQIbBxLVAnmIOJy4f02wc80r6DzW0hN8Xzh2SwC8IlWSF
+2CscrkjCZpk9FpjzuZdt0r63WCH+6bgKxfxMuO5lISeJdKX8QT4RoCanhapmc/CVBpfOtXjNimr
6CKBt605/QrTGc4FAqDuGj/g1GV2Qe+vO26e1Ye5F5t/OoCbNiOL6SjsQwEutG1+fGNOII9V0pxO
vhEeLFmR41Jg8Sl90f1T0agaGD1Q6ZQ4CJeYt7DgB6QOHQpxwyimNq5HE0Q2L35G8sV4pTWYecpc
5I2Ns2BORqZspnuRaGqV9NbZGqMo5rpjorN3VGWGvWU6gXQ7/j7J+xfYjZ8ihRmdTygw9YBTK5wG
vf3JzraP/UzzvLzi0c6etz8B5tFwEHFMyxrtJmz03XxO1uU0YvrepP53SX+bDi1UwuMV1mTcc8T4
5MTcQhmlOCK8p9r7unIS/CYO0BULwb8QIvqtPHmE+h+iqZbclU8Tg/5bUDjysetU9ao1FVnpjJdZ
I7v+cDsI+1Kydjz+XrShMijT9QlqG/C+KlM63XMnNKDxApuZAPj6hV5/dlWWs7DsP+U2h2uzDN3o
k7kNLq/tziAuRdf2XbVPzFlUYNkDpfWXHoC3vOHTeugeE+/SiZqAaIyyrZcqIFDJPvZWMzkWATtw
tUA01w4uLfDevjC+OoImfzPEA8K/217qFPOskJlRdVjnVpSdhzrxR9NjKMAviND1et8oj/p2hC97
bEM97WDrkTVYzyZBrp9EpOWUwd9U0i7Y4pyHVQ/BBQ75PSvq0GOFf5IZsW90u2m6slc9UDUXssmM
RXbIRfe2jK52G8v+Z3uG0dsUhlZB+bZMqDQxa7s09rv3pxPNkAaqpMQ/Xj1NfQKmyiYfg0Vz1J6s
96eXGKJx9cgcizSMTsP94YVrz4WzTjV4KyuKTkAFbsxM6DStCgDspbC6oVBFH/pt2CT1krcQZ0KW
Km6ZCywn0bMir3qeBVJJQK6Q/SW0xg0FLmtule3uLBcYR/rhhibREFihsMIZ9cGUEJThhUpruOIF
9VF0Mb51UMbBpore8K2HsdORNmWLvqEFzJ595zktIApUvYTox1uHD6up9NzwJQXH2GDf1FFMJwJH
YcXVdEvczfueCxR7SHpU4y5cHSQqmuFm5VTI2OsGkxeBIwy6Dd+hmOFmBPw2L3ZrlqS2VcfCfuwp
5z0L9i3jH10pcFSoZJGw7NsKiNImMROFyW90Esfsfam/rVlq6mP3iL5is3LymEFYnv8kVQmKC4bq
M5ShWPL3HmarpIDVAtADkmYMAav7aqtcY5JbkQ6F4qxotPIivnaNpUkmXQXA3kndmtGSBd3rTePl
YYoDZNhh2C0YQaabB4Cb3WHADnJU+ST6k5VRPbrfmQdvnX+tS4mEzITC+pwyNbvYnRjYxqX0JTk9
5iNbFSFatIVQ9nyHBsUXh3C8nFqBsNLZh3tuB9QmP8OpQ24H7Pd4SoLVffe3JzqHMEQa1HvKBxbR
6oGNXt8FJva/Mwr5J5djZfZxpBbS/uNu5Q+8qy/P3upV7qMrNAyAp8a3X5TFYk4tB/pAxbOr3mx8
Bb2ftrhJbK+REKS3D4ZbjjhDgRnes5z/Uya+pmRSOUsJjZ1dHJipatyipO5xFHd4uMehNOHOHQrT
g2tZn2sseZta5bsMDRA4Wi0mtqkve2OEBb5FrGX0wBrnLh6UHvs7LzMUZ9Gg1vLBzTN75bAuj3c6
hzeU6ztHShnXrjRU7eHyqWFrIw0NiHp0YPg/Tqe7UY1KH2slNdwJsfyNT+cTgQYaXbzmdU+I82yG
NND8aMnZJxVn9bnBQe7d3ZJO+ghHX3+TZuip/Mh5gat4kjJt2i0J9TA4IpYqgGFghEEflLIl4sz6
67zn/4RDmbhHtiyMB1xNTcHJYERjYQyeH0hfUPNj8NBRYUPl48oXbvPBVcFonXi1fhqqcho1sxOr
5zUQWXdxLHR1//MP8AFto5UVTgbcDz+cp2gtS8F8leDa1we8KikmJp9nl6uf3RNtxZ1K4HZqWn6M
SzZNXRHP5JMN5uTpORJwUyJhoKXvZfQZ5vFbHKtJkJ6nCdIp62vYsh199Hm58JkOyAthNVJ8pOi3
X03sima/2g2w3bCaFQD6F9uz8LYsT296h7VbDDm9kYU9aiS0ckZlor+Pk0Ig8VYVQKoMyZMq5cVR
9RMPJ++Mc28PJC34n+JR+YtDBvMMzb5DZ+YfxOM7yFN37Fd9P624eJLHvvtWuUmxZXvVRhY575vD
i9EwbCQBPXVZ4mgs3Fo/jZA1NRxt16sK1X3ctsS60r2njIM8wLD1v8cwkQwHyX4ck3j2XjP68iQD
oyJnrIWolujnjmcNmVsR7wtIsYNx7/vmo7HY66YCryZYbCYRRskYQWop/hrBr194NgYihIEHe7J8
NAWucOeP0iQNe5h+1QO4Lc/DvU9pMj/vp/64Ers9ZEeYvq7a/0mBESC0a4pKe8E4DqEE/PoJu1Wc
wdk2sWNmRH7ZAAsR/bRFP2k+7tNF+EY6LM0J8kJqIPHcjyR3vWhuaPODoQSSVCseaMaOdxIZxs8/
mpsEBPZRHfWO7ujfi5WXvdqDvK7DL+j8i07glwPNgvXnnNmwGxHlG0aDEjXc8xCFAbfNS4hjbQsH
7eGh90p0OETXop/EWOFSrNuRWWSMFFHZHvm3utm5eOeU7KnNE0bvQGTmFUsvekF1F4gFTmJVLLH0
1SGTicOtKKLZfYJY67iPZAec+HqThSP4r8VQFAVdQX0ntHJe7FuIPhOIpsW7ASuTuSfyokkvUz08
huOtvtef1VKIFRzQpQaJJOKbroJTAC7GpysQ1Lbla/A96mD3juR09Vo5X/HKk2ZT9TV/hITgPypz
Aab7o4S4Gm/VMowP4DdnRbngEWQCTtAb7u70c4zPJxJG3ZCNMihtrqnY81s8Ch+lqErfC2zvFNXG
H+S0I/TsVvy+bvSIL+wDLtGfmmImLfwpO38C6Oy2xu8yZxpY0ncAhQzz2NSQEnvRTYjGKvQWBzoA
VvEzUJ06ozgJqB9rjFeBm33r4NQ3LBV8veDS8RvaXNbJf731wd6aSX/tFnZ52HOyiMb/Z7J9jrjo
c7T6HjPIq4+uXgZaPSUhRDl6oHew2DN1ZeofNC5Pl+50h5tC5LiciPUpQY82XVsL5kBI50bdJhGa
p+Oezq6zrfCJaX+1EooOOcJQ+tUd+OmjjlD6VuaNqxTOHa9vc8QwhymMxQhBqBp2YBw9z5IJQGFk
TqPlV0n8jaCPUJirMDoizOX/0NNaLYUVzR0CPza+8Oyo18Z/vP8ybvTR6j04j7T/lTTHGoP9j6Km
RAbAUpotOm4Y08slC+phOGOIewSRBMFO+9x9N/TXD3qIxtJtOTGkVtsZkh7MkssVI3iwTNKQCpuq
YzTIAy/FOTnuctSjeuGx+q0FZ7M7YWLGdst/tVUo9SuekU7rDLWcxZQvvM4XZA/tQXMJ9HUUHPxr
8DsMLk6lm5U3iMMaXDIip3Q+SZGPsFSI13cg2RIvA40tYwR1YtMlpkAM2fFi9jeGho5stYUro/1v
U5Eo1Nk2wg60QaN4JsoqJ8SVC68G2ZS33w31pEP5xCI5cCo2kyGORBkbJIu/LT2MqASiVnsxvsOf
8ZGcfbKziMiHj5JHXuqbeCeeAeER7uTakOg+Q9EKW4RanMiCkqnDIyJLsr8XjBpyRH5WlhfFYgPz
CnpkNa4FC2KrdQSwbYyIYDlkC74rTP+oa33jSF/J1nvuyKAzB2kwrXrfWSHibNkU9VN8oJtdtmbf
EyAa4f7lXoJBki0wmxigv24VoeKTLMqlPvsXEu/hFysnHQPiL+h7HZZxxp0WNWJffZyCbPacCYsO
S4mDEfTTYist4TSGQiXK0MrsEDFCpCJx4xo0dJuy+v3fL0rjx7Zh5d8/EHF5ZO04LY1VZb3zS66E
CQuJzHhA7oHUn6NBOoBM0X/Ir8r4VqvO5YKDtykrDSrkxjubth7s0fzOwOCxAHdTfiJX3viJoQeQ
jBwrMzSqC5QDnHTUyPP/e0Wx9vXDcufeOVKp/t70SeJNVQHWYbVgEfWcTKJxGssV22OpbjAQPpRp
cOd4ziZHYdXenAmGKz5BxVbvp6Zt0bPF7XPSM5lHdC9H18ew2bw81R14brciuXkBDmUZGdyhpAxA
rfKiq53RyGvcAfC5EHyeVDRfW9CSGw0eyUhg9WE+/9Poru2smbFAOMMgL52xfhjZmKBk4oKNehC1
5XV3k4Evyyz+I6MVV66WT290wOQxRALEmR51vxq6z6hX0ZVPRwHdoOJ/HZgiU2n4LfZQTkGmsEyW
WQfasAKSQ+1zih/y9UkbdX3PJk8XzWcpFEFCDACK3bBiBtbqvCPvTTXyx8xzUkXcY9jqfkTpO27w
CLtj6iJBaKIi4KUY7CZihZyLgh/3QioLOtS1d+cLmVNBgXpx272CHiqkonWhSLuQ+wANhNuF5g18
iZ1FwpPMIOZ+FnFEaNqNqoJSQvV0Jqsbi/JXGbvn9Fahsij4uav/sGZqCALKo4M5OMOn1RAl35dY
WI2yu+ffhBiA93qZ1e7uYFCUiI0QKnUOzhE/OV40vgyS0BwfciGgKm2duumbz6+FNUO3dwz1DAb/
uJJ+4TTNmNl8UijqbKdZPzQZFQZ87/rmKAR7lJA6AWtDbJPCHy3efv+uuCEuJDzStGLijyp79SQh
6ReGDk502uZUQohuKii7f4QKoy1jCwZKYfVf+38JpqDyj0fwsCe3v+cVryFL62cIFDrqm73dai6I
MrE//BPlalTumnIln48Spxm1mhQfSuflbYMSpHxf++tzxlMpjEGW3UPzTVt61WB98G4rA/hZ1o56
A9V7vSDkc2bQ97aamdPJ1aUnrd7bckAN30aIEfpfvg+LiaA7dsmi1+gJRHwHhkWYuvfKJcfXqy9a
IapuKjzzrEulVdSbusL4LTH5XT0qZm7s7Avasx9OHgL7diPX25FKq8vPtiMEO+lcTfitUNLg9WlZ
/dBBb9H+tqVESUmUO5G5lBiXFsRXgyvowjMWyY9JF3d+92m2/2j6cpfAiQmIXVMzcHKMs+digKq5
hVESANuI4I0tHRT1W3sdmfyYqiT456wHodVmKm02ivJu22U/8r7uckAzTsMvE8llQbcX+Loej30s
haKDgUZY4kchTy0l0SdLPtiNg9j/SsMCijIieJORtg5pQRJGGgW/6JIFtBGO7K2WN12j9++vbHUW
Q8NIyxGRC4/fdi/xx516I+ROv+2ufoPJpqZ65VvSKx9cvQjTm8JmQTMSWEuXJV+46mo5TX7oYF5q
WSZya7xieKxlleBf94wwtWi8L1B0ALyVMkS4KXvmNCLkBHPhQoNNR6EAwbRuEB+sxauBOQzYYT/j
EVEg0xB2ADwJw3tViB33d5571wTJr3hT2Gh9vsaLJRVSVoZ+nyxqfVi9gCUCcXxRNZlh8/Ya17r8
5oYnsIZrpz+Zt6QRJFRxj4cvKSbI8Dw+pKApqxtSgUcLY1qsY5LnvNV7dHh8pZymt1Meib8Kcmb9
WAdOJ3f79hSH3p6H2fIl7Y6gp0McGISe3dbA1KzUswAx4K9Z9WrvGC4Sf6JBldiGBKKgYQOCcSGO
3u5CKkZikrZyhlyUpAWMtjV4IfYV+oURtxe7Eeryu8N4TSmeufo2Bpvaeep7B3fEh5TMhiZhQ2h0
cJLG6eAehkxuwlH59+yGV3IXR0vqUU+cqiGSIcGmprA433mJjzMOjG41eTHpHOunM+FKZRLn9N46
YD7EhPjdIcJmVOZRyLwI8Qm0/L16Rm+iLofIlh7j5LMYzP0gDEiFCtISceP5BMBSCr/Ug/u4UGUh
9SSgnsAFdiNhrbB/BGgOfTWWaSH0n7tRveIEXwFxcnUMJ6+BvOffXFcSCI/qVdFUuu4IOqc0uVlf
bzqa96wEeKPpI9wd0lALQEvdxJT+E4avl9MSuiskbZvsw2YqqX/cG6tPUjorGPZsHK5yNgplyciU
NqjzEzIKiWuFo8/NbmW1ba8pr/LTVKYXksVBcvr+54R1IedGfSYknzbhl/0pzb28LE8CIPKcbW7V
XxfZwRSyHCuIcO0lKdvL4lczx6pUxTOX85NZoZ0a1WK2LuP+ZjR6U393VelTH4asMQFYSn9p4xtJ
kZqczJPaON0fFrsQMT3pmq+/AWL1uFUvhXjholh7465qQH7fAp3INMXZZDggxxQ08dqvNXidsH0j
4GHH6byup9yXokf5OqrcMjIZanGLtEAE7EhLnvnuKHXkVgovmz1NF5jp+cXEGAtA+oN/88mnOgr2
mxOPQHbSpiuNsfwurgbjxfM7ukGXaKEdulskRT7cg/WhR9rXmIzJZpae17qw9AudhnKyJphsYrd3
LmlurQ41ZZ6uqIeUI6BG5qxUeiD2GgYlFm3BDgTO1MdoBs0OlxcQwxnH9A1Jx1YZVbZIzXV0RAen
q9eDpSbEJodcSGR1GlzYVBsb2RgzKrjP2MZ2FBcayJZstM5BWLtjGm+KRGzcHiFG+ySLfHc6+d09
iKQOKHJ0ATSOxkZixA388tb/2y0Pp/d0MGL7nDCAmD8lMLpgN34m/LcVGn5GhPfm2wXK8n5vpaHZ
Oo7+0ZUjOdR6vz/XJTsl0EGxvh2NvWsaosEt/ulYqR8BKcvW2vniphwDTQmtFaUCnj89Ffv/bqjr
lDuxe/RufWYSalqWi9akg7uNm5XZ6FSjbztv0VtDriA7SPtZZFSTcmYZP20GWzSwnN6Ai3p9/Bg/
E18nB+9+I8ePf7ZGesHsWP/TCU6wAwkMrVd9ILkLwXNT+EjgHBbsZr13SX/na5YAmicaGAzAFVto
S+J98pmzL5ETAhbG6yjBN/xqUBTEqQYjhrybYAnn5y3rEv8RXCE1YyV7hCER7QTNgwZeElHZMlI8
4S8KrR31s5B99MO0x2lPcUBpKo5N8JiPler30bd865ryujSAIpgMVYddHYkufRMlUEMuEXnHaFvc
3WW+wHkt/w4+YLneAhWIQhCnZiBcClrkVowb2R3OPSfrgHm+QARzNLOFkSDJQ4IcG7F3Mpu8ncjM
XZt2BeG1urWGo/2TXoBajaavWC7o7jd0/TkhM3su2u2y8Qo79A6glxYoYTVJX9kfq6jYh96/B+JR
ElGwIeGLt9nonWjWye7CxPB0PdSi1tT3c1divn4/EmyVCJ68Qy/3knhVAhhpuqv8tbYxyQrU1wYL
x5rTLaSMjF6DxB+hAaZDm8u/bZNhMZex97KL1cQqU20cK06ZKL3Cp8FHXwu+ZOcY/DnzHEzkgyJv
u4Zna58xp+naNS5v7dtuU1NBgYPALzrrRINKs+igqSKtm0jr6K2oZ6lr7xrEUxa932ctzGGf8BVE
GH9CGuepImogYlzKB91x4ORuHpzpe1DOhuczgFVyA+EC9WyPMOyGOMkw6rh/qjz7PnkRDa+SqkDj
xtNsN9TBmM1qfk/+4leJzVXh9MjBS1Mr5VhmF23el7/EnjbjgyxOd+9lpPmIL/tBSROCMKexGQx6
kp9YdymNe0Ll4yxdC5Qz+nrgVJZnvwRFf+obkhUpeFahS64xXi0sPqQAySwLk7BHe3CTUDNdp+kO
7wDp79Qh7oZEtWtZW90E/bO/osVqaXY1COEZH7WteFQsBDUOk80zLySspqIVyQr+DfUt9F9WzyWE
HuOhshEAp0sEfzXG7aozVCL+w49iI1x8Jer6J/wcYIkt9vD8yb5ChOjUKm3U5ZJ6X00I+rvyTRl4
g/iKj/pgLrpvcIVFtko2n3rNlIv8u+SZg907mAJSnil+Fy0koPHpzvXTiQyXlEdi75CvXsHbHc3V
On8impC4hzfX3YJsJyahG8IMvCX5M5SfET7YWlVAE/Ge/ERexN9sbkcgGBqD4mZP9gp6742HMGE1
0lZFP17c6VRBWlQXR20R9M7Xd/JEkGkZgyDv5cCqgNviH9vjQYclsJ2pGmcMbqWP1Z31kum6zvy0
LKYRzzvPWn7yllCoBl1lQtpOkrmGZhSNafOz+UeWsP0ixDCoy2ofcajKiXoateQaP9Pyw3lSZKM0
BFfsmtB8krOnispKq/16G7zpe25S4LiiPFUPFMHCWWendjl2lenyk2EoT9TOk8pLS6EFpCBFD5JM
QmT6XBhqdy3YrXGb1kgy+OYSBih5GxjA1deBVVczGaMB3Ns5KogNyr5MW6ZqAAU9pd3Qc4cxJlxP
nubRoZ/d8mPMoUCOk6q+87DqW34XU3qxW2oAfdyGUwlx3MvB5u41TVxeBNKTASkvWEgyUDXrrYMP
J2AF5EvmD6jq8L1THYrrcTvBTNHzlUnDR9ONqjATsG12ZZpP+U7xsa2J/fVcOwt4ZC4Jj5EJuDbv
UOYpiouH+dsxKWbrNhE/DljZw6psrrqm3EJfN+N1MAS35TZUBuVGeNYMXxfLeiixKwYzdt4bZvlf
1CkFvILanQXcxmLpGszi8ICrTmx2PjunArh00m83cmb6Bj0BJ8UUxAR4S5rNgl8XYQAXmrrKAXZ8
0PphHdH6CFfy7ICxS3YGtyFBttBfyeZsvtHOKTxRJ5BHgbOSHTcs/eLHw9Ga3Y5XJwFFT5lxG5rA
LjVkuv1G9pqkDKfH5K75lIZwbl6lQeeZqWvq8TCrEgvuabS3Ub3upisZBqrlnvEo9Z/MawulhoI8
Im7W59pvjaTCQ201zj8RWnCscQVuYOXg+2vI9WtWy9+mBiNv1iDntl90e3m+cI4TpEAc4vn/CAnT
3NOttxLajODV5h135Qw84wNenT9RKww/B5BRNTUDfk94f1UChusY/+z3qCjyz4rpMyTRmxfObWyk
Tx8FeHE4afOgyc+8bw8I7BFtOu9ygBqKNygVuhaQhnxbk/mzXPqTMKjsRkRDh4gxBEpXOE6lRn4d
eWHXkxNoPhwiYbBhbmuXAT9WVi8jKkHJkjoVcFUS/hjqKLBB7xO5jc5JP4O8mfAK2LPFHuWB+hZX
O33ZQxu93pHOSbySmrxJ5ywf/AUkieQitZHvDYqC5cxy1np574/zJWOaek8TvELhITSG8cYIjK75
/Vet/RI51d50efIBhfV6nmWzbTdaHfKJJy8e7StipWhTZiMlhp9TjbB75/B8h2KyjVtP4xinwwgT
roMH2n+rEutUvOHZtPyn0FCu8OWv6isiRQs7GsyLn4dtxawUp/e7QvXFV4BQBHcnS6RX8C/Vs1Bw
kyIdVt3MQqShbafM0/eWuyDj3PaZfGaZnAO7TtbjT9RRmyv1lLaqXjPOTw9Xnp6lK3eCRzXB5xse
LZUi0UaU6Md+C7B6HYe7rorPKPgLCtOA7EtNaJO236yMz+F983LDH3L+p1KhxBxhY/wOzpegVsNc
j9lqu8WM2yts0aOni0uyc0yjqnLCW6gnJ8vu8GPR4taiececvj4LiW+EsFIZvy0zRyw0QTi5UuDx
/Kj+Fh5RTTN1Hk23uMExAAasgdZoMXpQDAi+JkOqgJX+J3zX0WN3gzh3CjQ9wEpJXrL7/D5KjtTq
8cPb4mDdNRgjNBNRELtmXhCtQ50yge0q3nPx6DulJulvPp2epPlCSbyvb9vFfWEoyhx8anK+S2gh
vJ8ZgLf/TMNwQwadcw1parqmMCholECxlTMG5OUoJEWM+2f36ylAgdUukxgE5znfju4treUBv34K
Utim+d4+sz5zJqQZutLZ5L73VznXs6bA2nP4jHMrvIxlMdqBZhp0M9vNTiwNnJHvDyS6w8SV4og3
LEMbP7b6hpFFck1Nj9qFFnyeoAMH0t/qljRZrL2etAcqYwSvfOXgWh/OZycCR5bVjkHJ3Rinmx4e
ZjrP3Wg7to3wCInvANrQML38fqRA3vjFF3+Bg4Gla4ni1KJX0aQU+qWUjdeGRfgbrwF3JGllHyQv
c/Ydttk8PlW4KznEtnCwoCEqJjGFqyUYR3QSSC/eBVyc014Ku+G5qlh0nYADi6A3AThvpwOq/bYw
9/6DyAAviWYKG3hS1EwJCLol918u2dam+7/koM5MDXsV1zJtmijAE7tK9fe4rTngLptKaYw1aFBv
Ux0ym/I+yPiILNOhydn7i7I0h5YWc/F/i1f43E7H1ryR0nNhWGaypB8zAVB18fLBKeKwdw1eeAbB
5FgyQyEQ2i0MV3HGiAxX7ojrD/8bg76x6AwfvnUw1Fa75T552qSvLPkPZ+h74TKxGpcOWiKNKUt7
aB7sti3qWsNoMdJbkEAH8jrodW1sWM7LO5sNflHw9UEBaWqeHtp4Uu1NsXLAUJhMVd5lsP9BEmU9
S80zR242YYHYWmKJMb+52NlJRw6Pn+IcRhx2AEVCqYz8+Pvw4j+LnySNDQQ3rsXgOkTmKibMDIbx
ovjrQyRDuyID19BIncHf5pzk8bVOofp2MBVQOra81ppIAaPKG86CKZl97tT3JspXRKjKXT5kOiT1
oHip71XhMAd9y8thsSc6BFVT9eReTfaYbd0cgjT6ke7vooUKRtynmvoCgU/3Nc5hQYMc8cJoEWA/
aqlnqVFV9Ckx+Nn/s+RBD6D4SU+N89Eg7T94AQFOVxd1RriteZqIsoMu0SWUMqOUdwawG+OpFufm
cwZtTMRLZEy0Ibojs79ORuh82ckVI29hyejklweqmIkGnnjTYl7e0+gZlJAhQ4vqWZHpTLHwT9k3
SJK8tDPScvb8bzl+9R+mwK4HEdTdiuqxutNQraC58f2HmatrMQnyndpUDWvR1+7JFv6f24aqLJR7
4cXoT4KXOdphuT1eVCPteOzccfEmfCqSThQeD7y7IJ2oJeJiCKYtgRoLD648wkIoIFcAxFIXZxhx
l2mNQvJbB5xQJXNow0MC7h1qmOpBUZ86stY/0j+dEslOs1QhAxb7bY13j1Mzbs+se40DNqEKflV0
bhnQU8x2i3axXzC7QMdGC4dq3j4lYkkA3xAz6Xn5BS6M6kJrQmDIRtlGfs9UA55Yq+nMKDQv0clQ
2TdeK0yhbe/1A4n1DpT5L+jx28AafBni0u/gn1vReSTSKKGC7eNEaoBs8e5LQVIW/pEFXYo/OxaG
vNrVhLLQaexTOgS/n/Plqr846WT/8/EcbchYplb+igSvCAbTVYbrAfHjITwtt3KXNpSyX8qPxKlP
aa34Nan3sglYY1j/Nnyc+KsjarifpeBkqzHWMSwuYSm0QoeqSXEU+Sc6G34QhFqsb2i+20+gqP/g
PrJapNFT6bEZllxfTVJimKhW3oRZurlE+6dCjAcnxQI4xlpw08BP0/qGSSaLstGWkact+Ym3jNRd
skzh+DEwKTDgcj7p4xMG+i4adAb6DDDvVZse6NajV+11gV6CHmn3xyCczUS7f8fResf2rdCmQgRm
yg3rA35buy1a3OpkPHkqy6XHl4iCTrsS6HLRcsknVWbs/Y9F2Zc5JWd7mhudbSahNw1vaZ1QqB+e
JpfWtIIdsAphkhfZMcluOXCTdo+U6hHF8s8CKTlxHESFWDLWzdbheVGRsYlcNjD7TqNX1F6L5LMh
vRCTfPqi8f59HuuNR0kunsPoUbAC3Vi/rgG0fNOQ8IziCKaDTBYwSm6IOIP467qQaeS89QpTNRLS
B4ml3uLHyRxAsOwFoH8AfKOa5njaBZ0FHJZmk+R5sM5/vUySI8fOvFC1tdrREMLltWhuFZGbX3As
ulbsCr3lbHuPEgl7vweTnJLlchrd+fHqcHtB2Efiywj2jGdpUobN+8mSYtvQflh7Rxo4kr+ciRKa
nSTk/BgDZDgrKKJstT5wFz0L0KriyI+jDjX6FuLZv9/tYdsfd8BgFCQ8elK2mq3sZRHkMbE2NKqT
SRxSpnuyoj+IZC8Wdnoj9KUis1+tBIdnl20mFRnbxqC99qhCGXQm5KYkAYPEXS7AspkPhYwAljus
F4omiAFliAruhhRk9D4aPKrdsEXbMx792iul0xHci4x8pSEh31q24g2xgKu35c3rJ3y3kuDCXF0Q
z6kjHpDrK7iJPMlipySDP2nxByxF8vFlE/P3hav9CfCSVs5spkcoFB7+FObIjbh+xZ50ukBKY1h5
QOf4k8M5wzswvjjJPGpNInBGcE9gZ1F2tArBt+JCE4z8NqITGNvU+IHCJWGSp3g3zW0d4O4zwiQ6
KimR5qQHyyks41kLptu+bVJ4SU/jqunx8JWxbLLPPY0BhI+vKQ++7JyPH8PBnWQS3NhVpqpcbh/j
ddkykyqwBMiwqHQO9YoCTa0BrfS12yofSjhCqXpR6iUfW1p4HzAkRuG/gv+DklPtmMHdPBreuh3u
5xe95Pih2/VON52tTWj45+7yjipYHFF6Vb7410G6WFlsiyFr0uA5Gg/ZiURgGD9SAnE9VsSClOHR
nKCKIRlZeX9UPwWNICDnEVCvs5t6zMzYpjzAtcuJ6DIViVZc3cIsb/X/dfrQo6Lndvdyx2nv4Ijc
9mCzlXRY9mwByFjHE09cDYkaKZDO+o9o/dwTDKNa98EHlRXP7dyuh8PEOE+alWdF1sJPhra1euAe
+M/UCTGy5/L0k1jHF89DM09c1uYFsf/rGPurixfp6OqiRYuoSiN8bv7z2/6ODUdKadFp/bLtcaEh
VyayMI2QZ1Y9WY+9qURwLUB2Pk5FF7xIxImJd9sV4o5D71/pPbZZ1oivc7aBL4uhaldqup/iVSzd
pHh2hsHRGtSdaVCg/KC59qzjI/YgrFoIQEsigtzoyr11bJK0viBhPz2I5A3bPT+DLHZlwtFwsltj
DLamMDstHIsLWTr8HE7JFkB103ihTDQsO0XbSGCr7Y4h9Fkxaq/hkmfyh028rsXWK8qLWwex8T/U
SuFf4utypa5PsjQSPrz6BZY3wQEBXFEPtKMYLhRcWgFz7n+YV91xsK1PjeEtuohyTjGVMlJ3Ama3
d3arEcbFdxn4Y4zRdKLuzbbpwpXbUqNjqdrEYAsBzPDn6uW5I4w88JwPGtAJ/lo8SibRpW1pDz+U
J+Ogw7OOyMnaD2NKyKdgzqYhiXdXPjgneziEyjNSJ8OzjI+df5u519LD3mMHoVOelt5/l3UiLgx9
8jVP95TZDU4GYLgqVt4ZmBp4SHIL7v76yC327rUpXpQ55GWV5tBBasQTl8d4NoYCr2ck/nW7JIeQ
n3est3PAj25HBiixH+20qFacWyolinftGm9es69LsOv8NnITmgwxWJHE5mE2gHzsgupKOxkzVz7W
0oUc7y4lSXfpT7Tp6ku1cWrWJ+jkyvsReZgYj5mRenZ3bsHt2R7Rvm2HQ8LgNIbVbe+NnLzjqw8c
T9tUNcQwFcf123luqq0QdeA8UBx0OJd4woXIKfnEtoDMvhswBOEbf/7Qjl6uLVRNOWPT6J/RF7lz
GepKE7mcx8uo3s+glZiomKf5/nul9fEaoyLqf8rTEsCO1H2aZOFno1atrdQY3PeZ6xq2TS2KkPo8
QZ+87rIaraup43QntFC5wHy38pBP4MtG9wclv8C1soM+kRNLnK35DNVu/lJyQmwfoIJkCWKstVcv
rRwWPl1nxA7Ou2ZcXG7jEhSOFvLvaQPdPnTfy7f44UxwoymoF2y9W5nAengEFIDrUY29iB83sxWR
mTQBEM9MVwlRlbekCeVHuY1e8b5j2ikPauAa5jF+rpagbFwbuU04QX/p/ZjdlvKoFwEBebiGcJJY
Wqf/rriIkXmCmCwFnZIdj5S0GiHFuY85j2mxOhzfYbCyilU14hBA/y44zeTqDwWoTAB58eQHUIPX
iFcrxLaJyVHOxVWfq9Sw3nl5PFG3KYLDm0szosr9C1tnplsjrEu3JPB5a9CSa+zXq5LhOIvmUSWY
xuFEWIHFyxAksiMSofLB2J3fksPcD4g7hIQNTYSAemhaZHPnqPN6QHzJSF1qvz9mULJlVxdBYtAk
XyCa0x3KXYY6zE64ceFpH2yXbV88yeS7NfPLHOHI4sUvypH1omA6E6HpCUR4dRrFrgtULthU4Y5j
99/OiJEYMJpIKYWIkUTjKO4c6bkpdbLurnHnTQFn9xzlX7pZ1nfxJMEmp0CuVxdZQLseOtrdMWzh
vRS0JOGgp9oOVtx7cbWQ5bkz0AfXAFGlEYyxToXr+rd+vp69oQnlaUHASXtZp5HsihzfiUAy5dZs
1Ao64e/waibPaUpbOVSahs24Go+33IIQeWCFcy8kk5Py2onjgVNW57PdKLM7vF4oOoF119Si5Zyt
kjSYY7UWmsMEHk0fRdP6nfbGuptILA74A8lhPtsT5bGG/jm/CTi3YmpzJYufMhC5qewMTHHsVmWl
lrrkC7jSEo6+DvGXUsE3AE69WtSk1LcyPMPtHYAmNwLA8xaoWFhSbmpC1pni2mSFy6mNBCTmC2Mj
j/30H3akDkMEpl6Vc3BERr4M9eHtziRMHuHUYP3Yt/rj6Nfjp0kOMQDf56gxIwRbjegU+9SOgNBT
QOHv+H1PQPz11iLEJniH0XT9aPCVYRUhHA6rlBf2XVt3N3vkb5Z/Q1Aj16WBstbXEuj0477zF8eP
FPuA/B+jtKGW1rtASvI/SI697xSToJcZZAtsB4NdCL84tD8owhR+CzlbB64NA9zfmBPFh0vxrvxh
TW+KLphN4jZfHlfqREehkCRW7CeqhZEtDmEbKdLstXKwNFKmEvMX1HD8K90bUfHRnlmgiDb+s3es
hPPHhcjXzUVWXFyOjeYvy7iP0D/3auYwWAib6mS9NrFkcGGzgoi1/wFe6/IvutDGP2IZicpV/TPS
k0V2eyO7HvLXoe73j/ijVroELqxRcnHxJR62Sj/M/8In/w1MAs3MPJfA2q3PWt1oK34XiUim8O2O
T3qPkhvIpUc/Dpe/sqKGOoKH1KwBkSKUFJ8Ggg9xhL9zSDv0/8h0NZrK3BentcuucuYN3EwDq6rE
T2bZdvWhOTH2dbdzmWM3KsVcqzAMbSQGJtKuA8iP8LPRjxXHzRqxhtgwPpC8qyeAV84xYDY9EJX3
HEB4B6HJ2tYXatKiTzca3/QTtPscImKKnIEyG0zAGR5UlViET/FrPG5PIiMNsTlgTUHa18QFNbsr
ooMucvbfyS3b7WxauFk6bv+3Y4ZzowFSd4bVfJ59XL/whyvKNTK1kVBtZywnkWedW46HWr5j80SD
4U6SkJUXy8Gc3SQGhK5d5cQ4JFLchuk9FUOPcbKWAPvNnsm5IspGS3Qhmoz8f9qQhLjk1qkvrpY9
wLHYMB5vOVvVHH5fdPvLxtCZ0uD3xpzX7Fi49lpQMQR7jW8CYKDnZNkZR5r15Rik5dgMxJPexyy5
lcqRtC7T2ecvbr4avKfYWb0o/wDX00Mimu7twlpnrCpKd9vdo4AcPBtuTLHSZhXs1sjAQUNa/sUJ
uyoqAGRCWQKSRHSDKD9PGr/JMne5VTmKwANsNgRIGs2llXC+LSqOzckrvLL4ao3OnmPCtKS2Yk+M
YgXCrUjDA1MGakyT/9YvvHA/UcillN3ngnW1cJ+x/MfEbNY0GAOiThEYIGT2cuRCf+oncXu/352/
dH5+sDl/jwjEc56Au1KeccfsfCh8XBzW1920SLtqGEipJkNJ11rNHvfunEmL16TIlnEt28IOsgI3
+HSLiTk5rrBIsV9euUhGAlIPyvBXlVD81DcziCq3WjEJZZ2QFVclj9WOFA+UG992lU/oMfnkTi6C
c0ZVZSKYOW6SAe2cb10FGwYJVFws3EnIMH+5bjrBYwwWxbd+NEq7/pDme35k2RR46Ni62norCqCk
FiZSFglld0SZDpoqybf//pFDg2YlZLXlTuPlatGUFGhXsaU8wVGIFZoj3ns6uc3dYN4X/kc9Jd+p
NW/ORi14j/a314fl1+j/gOQIeIv01p2Fun1ypiw7JPCYGGCya4Ktj2ve3QJBGFrIIAK2CJLnOwQF
RcwMFvW7Cvy6PlAmX3vSJR5pXGTx6tPVt5ERxykd4ulQNAZjwqZxkr+b2YQyrzARBcSB/cWmnXLF
Q+Pzr+MmZfRljsJzeyfCdxN/G7F8yeflOdYkFygsCSMS8FYchijntMzL7xPsrFdrq6fce55g1+ll
hW3LwskTDYUMCLZ0Og2RbfvSGDUCQ7PKTmk2uSzUiKM7s8CH5VSfIehu/nRxnGjXlIjTP4fpDLlE
9DoXHCyD5GitmdutOCOAgigsK1xnWqKUbQ8wmzPJ8m3/sAPv5Cuu/z+KSzTdKntuu/K2sqgES8Nn
aXsWe0tj4pK5U59saMYfCi2oId0Y3rmU+P8r1qfKi1sLE09uNg4HPwSkjZ5JfWPB8NRDkbnE2ezI
didGRD8diNfx60aVSALBaQNO5kaLwnDea1BQBUJ7I1p2sPMwP7+GKfFw2Yke1VxnOLZo85YLbyxy
QkwgQ6XqhEDpYtwmgZ2ajsl/IAl7kw6ecBQe4XVMoC5m1WbMooziUjr9oCZ7p3wv6bH510EILgFa
VjhZ4m900wZD5ys4aiQzxR3QmkJEBZYAoC4BG12jUicT+2N9Z0ynAKh1CHvVexKNgbHpTcskhusX
Mk0bsNunTZA0e+GIF/7ahd8MOy5gKBNtEq0s8oGOOyGtD8Lmx8Q2x+8VUzY2k5clpE0yRBH0U6ex
uduxugFeQRN+nhKn/GzOkAKp6vvJWaQZWxkC0U+jUHxYuH/iP7dyTzyaJH8Yi9Np5nu2KQqdWnE8
OIhooFT9/dwk3HdrO6TF6e3DoQQsrcM+8LDaKUFxJSsseT3ZgQ4m9+p7MUuuASXvzel2qzPH+Z8y
cKPMGn0Fo4q4de8nUtWpqxzCeftTmPsqNJWuOZsayNe6D0X6supetdyLR3EXG5L6NrtO1kvDMQ0I
AUR2nMm26BPbTAFt67kyUdHl86tRNLBj9iJhg/gb5E02HQnQp2dDL9nKslhUPxReVKMq6XFDw7hG
F+8WmRrJG0utMB07JOpiDk/2SIYSeD8lKFmzV2DhLh58cQ8Hr6lmkeCEvEhjVwhpj3vxj+MBAmU+
J0klfk35/z/B3KQrTNG0jjX++7pOcMGIdQiyEnYiYdr8IQi/PoDayTymkHyvWx88piTBWsTcx35g
1t03g53o6xK777+82HS2baYugv3gPxJzgYo41Kq0LnMJcl81BTdIamno9TD2KmldwHKmn0W7TcJr
Gas0/IL6omV1rIu1sr3b8la9I8c1WgqBL01SPFCGWkyzP18teK50zGbHmJLhrTce2zxLRgYQ1DQC
HVq8FmlOZOdGs0UfYXxr2KNLrl8OStZaUeGO0bQDQ+3MapzCps5RS6rpAkVVOzEJOzD9+srGlXZ3
v7KzK5Wxf8e/GXXcO/tT4UUmuU/qk1gZWdmUYG7Fh8VVvAwmxtEb2odHuAgJD42isvLiCEf6u5p7
hEhPkl2+Zr7v7WIbhlaUZFbWN86Y5HRij1u542a69pPooeDCkpL8ZQ6UXysPvjfRDH/bSRebGq1W
3F4W0TVQEEc9d/YBZ7X8SdG2TkzeJky1Ju/LQ1TgAyYI5btkLlRowICtaa6/vzWbs7XrehJVp23N
o7RbEyZ2L47NqjKIoddEf6nSqKESx9Pmr5eQLw4t6Xl0pOaxmqHR+FKnQAOhLo9u1df/74pINxMQ
ySyq4dyhjPOIy93DwURVcCNeXRn4vi7/7vDiXFvz4KijkOsLQj9wGyE5Pa3e1ySJ8d97mYkrfRBl
xZvQjex/WmGKniTdGungxMC9W5YWXRoCXKbXOG7ChSqNiPy7XkxbGtY8vVgj6E8e+kMYvcw/aoQF
k4A82F6tqbkCRuETluH4dc+nddGGNmVH2owV5Hcxgz/dDqbubr1bYfNSgzdVbfLYEior6g15IWyg
OWIRTNYjQU6/3K6xwPu2HiUBYDrhXoQUDxhPCOCmHtIn9Nyh72lBkaFHzt8Z/TpPP6mc/TZsR1H5
ah1lBSqWqYkxqrkE52lBkS0IzSITamAXF05Ldoy26VOmpiitjL1/o05hL7MwjOlkGFIgh/nWBjqn
NoaoCyCjg7j438yhLbJThB6GoDR0frBGN2H1Borjze1ji73Yc3o2fc0BezarxfYHNrNLithkwul9
0lKZj4TjkBJd/tQ6PSolh7aUwRICa0mOid098hXjA6zQeoAdRyIhAKZ4r5mxV1QZwuCGStTqm/Cz
POg85UfGsAteMT7S6+H1j3DnikGcKlJf4ezojH8EHhCm7D2/x3ahHyZ5milcaMz+sTTzpzOpmOk/
q61n6H4GmdpUv8vwhV+bsgLAKyIdTkiYot11M/r3ropIcG7ThLLOCmF6FxEnBp0LHYi7m8EqUP/y
xRUlFBGtLRFzk/i8V9li4ZxbQOyT4VOkth+Ug1c7Rv9fKlvRNUQTOYnZGxfY0K/bG1OgeJOyB4Ct
CZdSPH7ek7mZ73v7oSiL3QLx/G3PvSy0LD5t5JtzKCeWB62SXOl01Au1YgQXJx9hTkycs77CApX0
g8GZSo6P4rwLktUEBVPhWrVNBDUM1XDLGS4dHd3tTTRX3r+JaKv/tjOevWRDsHt4wS6mP+ajsBo5
yIwIzXsmX/mSdyjxxPcRX9ZzKO+sodsj8slX6uKEqnh4DlsldnBak/xNq4Qw+aA9ST8/l+AN5TFq
/hyaiaopTAxdxO02VapvKoCnas3R8JG1DLKioBXfYqRXN1u/blGRfbDCYmISqR2MRih/+USfaeS3
vUjrSwqMi+i1j9Y7OGtcloCZ+GAOoCt8TXM665L2BbJA1JkpNIZ0JF9kLhUAUPTw7uEkh6AVU5Od
/NOsKHxpqCxYXP8goX4ICBnAGrVcwuX0Y8/3o1TPFeHSo9NvDCZN7q+1W3MJazCitYrRhKiPBoz3
fi33pt/rve4VRVEkh0ANxQDGqsARoe+/8nEFU95GTY99BP6pMR7ptthEj4qABBFQcstMPs+w7UpU
kqYjryoo59q4ysRuOfy6Ux0t8kCtL6RP5ritOQESpaR3D0YyXuZxQECNJwbMen+AhKKNhV/B8GdZ
NVHANgMsHScZDcQgNLwY12Vq4c7tx+jeN6V9mS2bFCvX4UBAE3U+to/cpO+zkcFo7xjSjNDXlsyy
93IuEB4KahmGSEAD1rEDYyzjLCyRtu68qljP8iovSyKvtmSM+YabQmnR5oL0HSyls4kEjsXPtJEZ
uIWCe+ykrycPMPw5PVDpg4VsoNRIwOhtUaV07cMbs+RhequmpXHbkuu/mypvZ7ZPa/NlbIIb+aQO
MpQj6y7PvYRU42TT3iH57q6KvNgqc//GyMD3FYFfPAT0I8FF7lGiDiU2rOSMczlTB3YMYoMcxEoL
D9fHGHj98XB+PYkmfZyt6Un8kOsdkKX0+UnsXkz0PbLT75XP6LPFePSKR0szTFFz6fsmaQQP+eQm
F1lHLoi3oQ6TIthx71Rbq6Ci/z28RvRn6zEKJ8z0COy35Qu6fYy3OsyIXmKPsiN7pTNnURr7jfof
J5cO4N1bsclvjqQQFWQSrAJynA8c/y3vG2ekgY6PSR6vlNSytUJmPBr2/j+qokht7JOVb4tBxG8D
Nbm3Y24M4XQSK6tdtB7dsx2djXd+RMvlTJyyoEWur3i1f2Xt1+DtEQhy11qqlv137I16woNhgJpF
PEPc0NMmbM6k/QrO1ztXOvSeZIyh7r42VhoiM9Vu+hs7LUp/G09kyJarz/yBPg7OArSjd6A0GTfa
ItlixhJyUtuvi9L9tKMzoUkvUt1XIpShPeDaZVucBSWVNA+hmXCYMTQ1TDs6BD4qfgwhbc2gCiEb
pUeME0QXlXlUmHD6S5gXBpl9LvdBfJ5WBlL0HGYTGTuXVP1q18KsCblcSm8jIAAlj5bVbiaTFvrv
niYIcUcdF6IZOP0wGVLmMuyXiSm7Pb3llyze5oLrYJNP7dY3x61zFVh1ZtaPvzJ7gut7hPsYgg3l
p0cQamnDpvFhbjndRH6tZnrPh2ITOp6UTz/RaabEVU/9Pq/CBYjJVZtrr8UyMr+mvHw/XgAnpSBm
9bbnCttz/iUB5J/jmjInh3kYjQb82OE3WfcrvXMwLlCnk4UM4s7QTD4Wv5lU/HyJUHs6pN04+AEa
ebjmIj5YzxF9k29gcfMd0vqT/pWYCkGsSM0KIkKvJdOy5SDnoDB0hlWr4Dn1t2kbf4APwGq36/mJ
`protect end_protected
