`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WWOUvIk+KRRub+nVQ1Xjn1bxLIzlyhNmdprOvPJkZNgxLGKVYNGJWawOC2vhIDwiQXdMs9vtSwaV
4SFD3AJiUw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DEKTQXmmCTM73HZTX+rCaJTnBI9IDWyFS4pS8gwmMog73PdT5vgkB522mRcuFtfV6V76mgFeWQuU
fTAOe75yLr93ky8rjF4ScQqoIPo7JWqBKdeMyvlKj7EHJ4DZEuB2iZfZeic0svKcVnVdbv4nud5o
aQmMtIDfVNuCWKZm0DU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
h8kezR+zRPGtthXJE96CCiSyKKqstBQzTH050UWz/WuH+1FS+Xca8K7o1tgVhHtpMomyIbb0VnRR
6IV/of/uBHJlOcQQUWPeUsVI9u9hJvHLeT0gcN2l8UBPBVD2rv0Y0Sohw5znB1L7OjTTlXPGrBRa
HOBPo2mMFmHcKuJ4wsOaBBSMOTaN44LuTpWBy2UQeSNQlrSNcFAB7WzoastWbQ8UBeibiYNuDlo3
rd9+5CBT/56vqJsfE1N1p8gTsLVcELCUU5Ckqp4snIwhg2SOnwlqlPYGiziqcm15jRF3EXxpaQRX
SMDpGfFfIdx/MMSWPqvt5GuYgauf/omuiNE6aQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fxkVUjEOM0hPHq3R+6jZOnCSAYHFD5tNZuuuGrgrNKVvBWqa25uuZt+TasqoSLYoeJBu3Tr59c7/
5MOrlhFdBYoiByoR7xooXrlW58IBjj5/sYXvHIvrSJaCnb0d2sGJep/0nxlqHQKSZvQBxpsTMpCa
y1qX8P0ypilgoj+UG8Y=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tKFPFsLDOCKtOgP14WPzVEg1hqU0HL498RNy3/IieAD4+9kZPXUFv5lJ2PjwETeE0ZeriK6JwyY7
bmuoVDbhilmKfaYQvnj2oje2QY27t9iy9ca6OUAI/66HbdFKyEQ3dqdaWliLqe0DfLfwu5TvfKkC
1Lih5WVY92nVvPDm0d6boipSGkHlgAkToO9dtKNaZ0NGF7ikQolkfZz7eVkHjRrklk1FuteLsAg4
9ErST80tr2FMPsF7AVGxEjp32Y5MGoh9/4wPNVdR1t4E+0bV1oltXcP4ohAfUCQ2rHjZX0XL0YTw
bbq+3568snzRvEjY5ABrCjzf1ufua5mDsp5YNg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3248)
`protect data_block
sl6cxsms/Uz+pq3XGb871we7NsN4UX3VfRNU3QSPNV09DwHBCqPt8s43fV1KIw84i2AB8em9obUm
OSgddNxBdE9b9OYDx96T5INYtBPv85AtinrJ7Gi8+B9ihCI/sNAEdXQsEyz9NSSh2+4pf/qJOOII
XSqq8WPISVg54v9jSniJWdx19+7X/cWKkQv8qxjm/jNUa1Y7r/tWXEGPSmAdNnJd60tKatrHeAuq
54h+ymaUakQnWR8/vEoPfB/7WQ+Wlt7J61Y3sADqDyByl4cTyJ84pmm7OOMuog5GIKlXzyNAjFHk
Axe51HKeLLQXD8l0g+fD1xkZNG3NZkaBNR9LVdkQSJnnvfJvsApyFjgN7AZP8Rzcx29NjJ6bvvAB
nneYBPW+ymlpf3ARGwEVVPxQU2oPDvxSGAFAbZKQZv/13z4rj9C7sX9QQmN2FW8wlMzwCMO+9kW5
Y0TZPPch6Pu7XgmRvOPO3JfrAqT/qprDhanzswlc7COMH1aTI5IBQby1b4V93+XsyYrNw/F5JYxA
ZqDEPrEhe90cmfU/52sc0glB5ljKvkQ08Hl9RFebU23hoGJM+A9T8t4prWUVBBjYT4GE750CU7G+
zvk3H/eMB8NXCtjIggsbRyoRdizqF1oIr30QYR4jVv05YY2UTMHI/c/MWRB+/zwmWod6VCSQLCMk
2eiXpIk+LY3CYP8rHrCeUpRtqPtvUOn2aMcxIvBpSTdFnGaoDgpTxBGlO8qYZj0+N0wChW2Qo9hQ
BiU8643FeegxQ0v7pTMglr5/Iuu6ML7hsydwkGDVj1J7dkejc1YrbVY+RifUgZW723gwYQ0gHgg5
HlM9hm1WWgTIvhmF8kyaRWgx2OE5HqjDhAaD4Hs6qu6BIxRFHi9MszMsar6NmYD58Oytnyueit6S
jbHXVj68omtHNHKhWuVZ18yvLRF6ExnZ1D6jpAyAc2bAXQWrBQrjLrIJKKjKD69yCin0W7Zcz5Di
19vViT3+ZuxDAMFpewvhiLXe6DQCjACLzmdQMK6YuL5n02egOzHyqGC+DrEzP/zS2yKFXf4v1uQG
5rP0ecltRfVcvcGy7fyTm9QHGPs/x460auVQEXM2F57NfALUF/XeUYZb4Rzj/NlZax5PzTpL29P3
PZE4+jPRCF8oRMFMCb7L85nHRT5AMpB6r356lvZWR8qZpa6Ba0YLxkjtOKTKFYqIIasE5IvGLSMc
/jiatte2Wt8VGCNU+CMvDerbUARaVxUGnnQ/OKWJcqdop3GWDJgoebRNrBIHPv87cWMOuS7+z8Xz
D6nK8Gi1ZkbT4n32TEjxn96Qbt+xp1LuEPuT9aZPrrJGosW9YHH6MzmFGwzW9G4xl3oJXbWhsTp9
ZKP4CFoKwVkt/zWzLdxXOqsSQdDf9KqLnnVhZ7ke7m+FD8oBIstcyKd/10WLCAJayU1hC6B7q2oU
43yCEOucY8HF8HWCLkOHa7jMChsWzXH7BVV+Fpsp07Um+HYhrwmXPkHBc3kTD9fQGlSlWyFY6sqp
ijoKdkGhyNfDcShXJvU7jxqqKjmDCxNRLmRNz1qkm6r6JmU5nDJsaNx2TlgnvDU5sMjIXLOyLDU5
kq2evpJh44qKnt/U86n0mKNEEF601Rk+Pm6U4jDBxrV2hT4L7L2CR8r9dg549fbppZtot0e3XyyQ
zaBPUaca8R8qU6PmYva2G4BUPUVTStmjgkjdfEymulJMAgkHZAnc+QNUIec9Xe4URhUxv8K63VIw
zcD6+W30K4SOBKHwhFALileepeiCj6OFoO2K/O0Q9lARa5WEaYVje2j1nWXOeqnhq7RkgcaF7le6
xX+s3y2C7b8paLFAeubF0/sJPafklspNJ5EnRzdhFyeE90XRRdUR9KrZqg8weqmI6InmNu+R6cHP
C9FMQ7YuX9cpGqrrxCqbzmTBMRyRLw9t+VJuYnNOUTbXws7qp+V9UKhqI467wEJQ00I2wOqAOz5P
X0h7WAUkzMURADMPHtjCj9+UysSITAB8I2iQSzATlbACoMIGK2/enQEo3hejACKs4VT8jmWa6lRv
bZwyRgN7T3lerL+8y4r/2+iWZKgvvYVRkvm+W7XmSdFrW2x5OS7ncYddySflliJo4/5/eg3VDTp7
dv1Z6Esz8lMqUBkFEYSQSJJ4Pk9TFph6H0MssbB6leCTUAvHuQIflL/Exl/HEpjeNUlkQiBP5H/N
fgfskN/4nvIvPV1Sca2dqR9rValzAfMi+D0kvicJsuvUnSEzZqAu2zBAW2qobe4Gp9NpTzJEs9gI
U1+YGDhCQdviE/L7zHN6H2lvPlxcDtMSqK/YqOXpRIKe2I22xzi7Z78fz9lvEw7J7g33XWIfzVgD
yH875N7HD1gOfWLMsl3x6/Z0uJBdzALC6wjg3+XGhPjkZcw3RkPnZ8bw+4S3huuXGwaltGj3dw0H
2gui6XNN3HPq+lG/djAqjO8MNkXAoD7Fa7yt3s6HXINSi9GmIsIdeFSwGTiyNf0rRmADb4H8wZBQ
rkN4asLZ6RmyK+NDV9uCu5gWzAwplVs7OBPSEBu69hEt3H2fU7fOrZn5fdxDKucaYSXLzRvGb2Ua
FxIym6u9axhjfQoHzTmDcLJ1fw3ihBe9LPiLdQv/WAH4c6aSlbICFekdtBJqOD3+QClsAilC+ODl
fV0M1zqprrTiYxDRlb2RCKJn5s+bj255n2aCNS2eXj+6kPH+foAUQfZFbQgR8/QyoWjpKWjqGoxR
YWdqLEu8auG7uGdNwVa3y6iE66Mmr5cys/hpkA8JcCIABCW2HnPEZN1Vp4oGN5Z0Jqg+1dMwi887
kVFRwVFsDXs+ExqNLHdmhtThWY693DSvylARgcnlUYVu71/c0jce+sQDSNVHCO4bEJTAUUt+aILv
PyER5fMqEpTj7FdOTPqW2FgMlimKGw140vXuHX0Rv8ycof8r8pcDZYh1rnL7O/j5qNNTX6qebzTA
BSPG92ELl6TS4h2N4kVjJRLfrP5VXI1GMDBZoV8IU/LKip16HUY37H/HWyetIkerp30cKS0W4P5C
NuKLVukhGnMXmc2iHyYySnelyfLUbFybIKJ/nEXQywePt9QtccVq0UDDHHv7NyTHOwL8CyasNicX
qjgsIEVXILzOT4qRsZfDh80/OrpVKPsmdphvvf9P7tyJ0gtZlmxSFEOHN82gDbN1ydBNFclmInnJ
X2EcXsTcgcwgyNZhbNnLsnvvCkDa/57Usi1JXoYuGnJijCwdd9ZGjkgrVFTMcbNVvAJ0CH1bJ4Ln
lYbIJNJkLp8aw1mfVt+UIUujsopQ50xCQIp5t1KTi6tcA+4I2PR+i6AoGrqcw2EFINH4+iClVAoU
aWO7nxKAYSbTtgA7wOyAhoP3jyCdY+jOY4klJoAG7etsg//wuNmjw3OkBh2Dmk5QIJO4IwEhD6+e
NVPV14CUKsNaoLd8YB5hVj7uL1CVdhIcJ5sRnj7uic/K8zxA+//MGInq9c7zoOg9l/gDUtO0ZHUR
bF2NOYUtHc4M9nEGKBzu10T2Yk/jAKfZhVcC8NmqOk32tm6cD2pkVFLRmM9HUJx9NwrntCr3NsiX
72cV9FQXzN9DpgLVq5viXAEMjj8jByV4qTTq8P2oBbU8A2UbJpnHiLKP2dHHmmgiAl0kOdPv9n6N
zYPID83ajscINiYHR20pMehH5YlZv36mLT8+aI3pTcK+p45to3lC9d5rpqGBtEooj74piMZUFHiW
JskPYO1kInTHusvi+tYmHXsMVIpGP82jizTfwOWWQdG8BCRGaoxeOozagiQM2e/s7m6g2si7mWqP
tJGgRNzo9s9mdcFZvrNYhaDGyMcQjDlRLW6mG/q4cHHBom2V1lHjuM4bQk8aI5ymwYitV/1EOrZ2
rkbVaSn3xXhH10FOCWLRmvghEEFusCzTRsNsHmiToQcjP6StFhfFPijdAfq5AbF3qeRhHkLGhG5L
36AHAFqUY7AwV6N1uMxNv/t4Jol7UXuIqLoePw5P7OKRzd2uFSP0D7mk3VeHmDR/IRRYHXUaD9rx
yBCuNmmrj50Ferqn3T5twvAbBL/bvj94JfpNudgSV2ScTsxk9JTMmiAso7iYuIpQDw60wFUFYE1v
tPFLYRbTBcs0sk0K7JsZXuOJygHWCMH6wgZgrEf0lM6rcEXntUU4pKnTidS7A+FkxIyFquUClwDO
wj5xJSGqix5xPTZUNDnT3KUzxmcgzqI9C4ez8YFcI3ehzTdFQWW4kbqn/NB5R57nvrYxHPYShLo3
QeX90ngwV+ee9PatdQOl21wW5EWVaJA/IXg3HnjehMv2PgyhmY+4JyBjf5XcQ4Wf82mU5odtTi8=
`protect end_protected
