`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Nv61Wo5nJyM+Mpb+NNDgsBBvIUnEJkpyY9HzwVD6RuPuHqs4xvF07Iy2EOnqvpg8gI6Sg49y3rT4
exDwUp5Sbg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XlqoxMmNEA5NW9h+NwqGOhtmOFtxlLFt+OLfeb5WudSPjZmOesiRU4OkzaHKkkfuLLddPvrQnejA
5Z2oSKAaxPgl9e7WSaWTzxoxZxNL3rJQxgY+UcF26rRV3Yeg1pGZ4BS27Z3glD+39jElPdiAJ4Mb
N5h3/wD7Ea4PtRS2iA0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lLOYoJvyVt/yVrasVQeLEqOFi/Yn6cVS3kjBdpih86hrr12pBnH4cH0F9+6K2RV1Q9aNsA8R217D
rBID+drNllZB5h1139V1Tubn7mKCqOxWb0UKQFYtJMxpNuhyXjA/nQfAtwOkzmfyMbljhW1Xx8bf
7W/I0C3PdhnKO2cJqB5JQ2n2HlfEvvoDLcgvZgbtwTJVBZ6Xb1tywJx0CBCXrs+D/mXZZyYxfJxK
ugSin8QZGfnnRbCyhUfhwuTsCpU+hS+e9HUU1Q9o1XC03eaBbYeWgpNaN7hbwfjxDhI1/AtYjmyc
HwvG6ykQenT4wBwWENQJQz/bj5gxVLuod9mozQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TFctFa48s5x0jlTcOfmPy8vEcJcT6hTOQE89lTA3c+YN0+VcGM+fmBBVliBpxUXlS2zcIfhkAlO2
x56mbP5v6hd/LIpH7Y1EqnhaT9Fh+aN2xa0pqoWTk/hPVNEOdB4cB7TkgKhLcKQld0XWXne1ozlB
XOSg/XVW71PoqgIQkHc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P3bwPCrmfsUv/qCzo1XB87Ut77Q364szf4gDsDTULx12erXRAEp5tOtk/C9qrwnSwxv68CRAkLyE
dCDqzWGSLZOPuwVeNPiUDJaXJk5DSX5+Tfh0GUMRAU48X/Q8QUAOTOCIYQlKfmmgVmIa0094838x
RsPpSiZjDkDuB+R1d3sHccVxdllHCpay/Xt2aGCAq1VVEbXDA7BvnoYJRtpGz7mf66KsoG20auG7
FMeljbtB+oLBFYbqlRWJtXJwTUtc3RFm2lqETHFyvZ4TImcYObCKKN/2ukysTOcv5kJ9rcJ59u00
LlnI2nihw2qwz0zrNNd4879E/YCnk5HGQlqS5Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25088)
`protect data_block
7jfhZJd3Wo3toZzxEMEG6rbCDnKuetbJ3R4ogVSdgeeRUz6kju0AK5Zc15GzTI/3XkISAd0Y6jgA
V+Hnv3/4ojhj5j1JW6YOZsLfmtG1ohTTKf2bbt7QlVJGOf8f9AEza1HxRreksBFNmA9QT9i/45Sj
Wq3HSZKiYkmv31x/lNxrEYDJUfYHhQlFV5bCZh3bn2wFMgkv2ORLM3vDG4FrlfpCVwiRb4Se/qFB
OSn+3h0w9S/YdwyQlwn4KCp2ltovVCsKvxfliYsyvSQZCA05A5boSjzgR0jPJYn55MLb+gXmQNTW
U7/470GzzZN9jYOXYvn/Ar/Sgif7Dj+VXdmnicPqznnTJyWWMSxO/C9dGdP13ryyxNMAsmydRTGM
Fc5y1XfNCmO2P5sp7quuNZDiWebBx9BtyZ4sjGOeLgAdcxlhIudCIfDd2Wu26ZY6PO5c2MRFjKai
23fJh9GIrHyXq4OcBriQgljs/0VoivKue+o4axsI6EzVtCjEoi5OYIKDxDrrFUs2gaXILPQgKuWl
s7nZJ7BjNZaHlpuZ8mHmYMJlveiqbz7RBzv44VhcOZP5sZJwc6VB3vEesQmbVJHeFtyGr0adUghX
JoL6yhdYoMO/1zSsPJAhk1IeJqE15plQENYAVWmondA/xFqodPrQ90R//9gqfqsQEkW/7rahWaNH
+Z8dctVoJwN/n905GTOqOV8lfYbTYZA7ZMiLGYPrytBli35LXqedZrxD37XtnX+++j1t6mCzqksf
Irdjw45gUbovpqnEJ+0pMRkMfJXbnJe/Zxu0cwG1Ck9N3JBmKO/rEzJV4q/xwQHGOZzhP1LZ4sKE
ftacGahiArWvt/yT3MGOBLmM2GFFwE+a8yvLpffbeuh69rDkxp2BQjrxVzRaO86ETraLqsOiohKX
s/etNJcve3F5pPLMb+D8PTIu2QbbstIDoftcSHrrrauN8hM3KjeseAucNiPXnoNQLFpkB+AbyO1X
iaDZ+qRoB9h3viZAOuvjKYxFLP7SpHoh8GonVl1cGY8LS128G9pd+N27FdDNIP9OywfYxgr6YZmG
8yG98kNvjI/WSsR3t1GFePBKUDbFR+5tmLBnMaO5JeKfSFbRUou1c2nB1Xdyo1o6yTfCA6VLwRga
BRwL58Ugg0GAyWBgVxgYVrGGAsYjIzI3NU40tQEhOeDjlRZhp3QhmA0bKQzWRXkaG5yWtnaaxBE9
Ty4Vc5unBnrc9NRjjmMek/lynNZvl4P9lnMfgd2c+2ljyKuhbFC8xzMrD7v5kXs4jsjMR8X3RvRp
ASZrhjkjkS5/ZYqz/gEPnnTP2ptxagnUebeLZPwdwn4NNhsWu1cw0ZEke3jUWPtadNi8eEQWkYYB
bGVVkx9A9PiLIaiUNFe5kWWKk1ctAzfXR4sAhZMgLdJLEZI4it8Cm4UgvsHabkEfLvJHLzIHTzWE
22UJXKRQUTZeZnNWGIBMjGhh26l4zSyRDzirTqMEXQvE8s2ZFgZXnt4c7rH9z+jUQT1sGMKg05KP
xh6jLca8tWSLK9kn4FDsuhE78NmtIkzg6Zxsz+ohDk24at3O/OYTSvZ2YMvSp1DxD92PLsqa7pXK
36YEtk3+ixqUIqKZ53JhZKWqvYzohLji48HQecTYPZuOozvOHYq7YsQwxXjQIcmxhC1Cr7PTDKC6
vI5g+iJhKp9GPl8hFD39bebUJxSr5cJXY20k7D+GHryOLEgHopNWVpeYLj4WMMxpfkvRGoYEmwwB
PUYiecY0pi34trD1hGkj54uQfwSdGqAtxzoefi2i5DavfggzHCnpQmHXZZPPJ1zJgyCyA0T05Y2Q
nDoZ7pe3eVJBC2TdMgdygHcV4Md5eGxyG/9/R+tMaLvMDYtfbQnsbhs/U7/8K/N75jwITp/E+1/n
L8it0GUVFiJPgrijbKwGcoJT6EgIdj24loz61wrVWSro+17ra/Zb2HyoZf7EMEUrELLkrklAvsdB
Ws7mmfGbpK6vxpCbkIhFa/nUGFM7dzp3p3kX5pPg1Z5M76kpp+Qicab0Q+A1NcEexXd8LCylUndn
zPbKeItU9QbdOtlXnx+CYiHW9Nx3hoVPKYcwNtDd8a0L/G2EkCnyOCRjWy13MuJkSfnHw8YD50Zi
t9+zr6NLAHs5MS4X44PcwJWwXIjq5R1ge2gF1GddpdfA8IZJmgOZCvx2aT7S/jEoBuW1pGV1wjZ6
w64W9DzD6ZobUEjjwJwIO99nmg6aRfK7D9gJyMLKfxNG33MgA8NyWLtmmgYvvmImWyEFt/3WjJ4o
8Z3DGEWiJYq+Zgm+Nqa0p+Ze3M02rdAw3arFBBTSuqdBCMDYSFLxAfoEL1JEd7UG5S9bdeOyPfe8
mc0DSKzykTxBhonHjJyNMBP7xnQDwQYzL80bcVQ9XHDdp6Q0KGxT+wbr/uMN6Nv7U0BYA0aXkyar
rDMlvP9nj4Gm6r1zNOV+ZgKXjpWiD+pCs6s0goDKfOhK0KiLXWgDOxgDFNIygTz2J7Kg1zw5Iw5G
807V/aM+G3IsgtJmz+InVIQooikwlmZeR9cQhuhNSCqjrlrg1uN/wYFJLgom6DEbT4YQfIvHdSrI
ZmaoUsSIdPdhAfcS2+rw4ITS0nR+z43rE6kNj8kDzSswqAdF4Naj84zPnLSipMkLubyjaUc3+2LJ
K3H3WO3W4Oqa/18IVEqEVY54WbDNedSWqQy857mEB2KnKWlkmIeA23IyNGeTUK5yeLkuLYJrgAy/
8fH8yzDE1nFg5kacZmYj9QIHx0BWSVR+Ed29g9gPyvTS/wWeLAMm6WPA0QmBqS8QX4TZ/1MkthGx
pkC4VmYhgL+gK/+at8VOFA9DJHxq+rAOfhDEfxWrYE8hKtNbm41hM3jedmW8A7h2HF7BMQ4EF0dm
X2e1gj4dd9WurPuI6+6OB76ojobUY5adatJwkcPsbWVSKOMyuwRDGsMjMGwrBQvek0gYdiBcUYWW
YK5RLiyk3DQilWIZHMtuSxaXCkX1zYbxY19GWnurjU8dsDDFHWiPgsymyDw21KKB7kex6SyRyDFI
oMfUMjzAFZqyqjajT28XxFlxf464H8RN1sxUme0PkBV0fi7EmfHuXqBqDkebBHQE9LZdkyFyKsY2
6ENesPFAy1KlXZbeV00njRfWmd+dEJ2Cn93aNkCs9qUw3ZwG9jLMe0zTZBn/fzWo448b/UxelH93
Dlfv8rFgeTr+DHFwuOhGQZlWb09YV/AyN/LGtVUIb1xef8ZoyDaO/7O8eXM3AFKiotXW0riimCpX
qc7eb6/6PlLk5L6j3kqJ7Z6VlZRrNa9t525KXP45ipDSB+pMfD5t5GLBT/iAZfv5BJMKPb+j2zwc
hR0Ijmb6KWs3L8w7l9BZIikT121eAJjeELAMPiLIW2fl2fStT/tMO45IRie7pw7w84ZD330WkTK8
FsWglalgymu8G9BzEud7QWSsYe0xzasbSLDqetu2CAx+bxJ2PlwbsbBnaAaJqV7CsBkz02Cdsiuf
yxQ/WY5Y9nQH/X/jvUUxMSQR15SGVBhiFJvj7eRP7pBQRqV/AlLmJElvSzeAgP+b78QN21FhkZZk
O5NYoi2jSviZAZUEED+987TDm1/ko+NRxykw4LUeoAYFzUAbHzI9BHcbIASqlD3ob4UafDi0yPYd
IvX62gGzd2LHgZv3fuw4C1an/y2xKwGm+ojlq00XozQWcoZZGO5kMwLxwCjFxkcG77hOYjYZ7mQ0
oL048uzkkk9xSsxqArHqUTDm5O/vlkUFpa90uBZd844gz0e8MKEoygCbOsnASMqLLMJyAmGcmrN8
xeLXDDPku/CFRfWuIxvZg95wJ+JoDC8Fchj8DF+HLCCMnM6jDlJundo/ukqtko+NFmaxwmWtZS+g
LUNc/Y+VyTnTCTYnLr3n0bxFpbP934dLFtRHaqVjDWK8jqSfzNYpaU/zVd4HgZfP+goHoUl2BVmT
jtOwxF00GS6CAjD/4H/eC57VMiMaCQU9QVNH5CK7FBB85yO4b4QRswIYO81YHz9PMdlf0wtR+sZX
V6dc+DThs9+5WhIQ+hvQOJMWjiTFMidOfjySt8QDeRHH6obw7M0wbixE3aCd/sYnJ27ionSpbk4V
mjSr7c1ioCeLF/+kWOTnv5OK6Nau8SZ/NxzmGo/Y6LHIbRLkPNbU05wRD1ZZKkvAC/dCxVVN9vbo
K1YGokfBzWXdVnaVYH/0nAEAIasIJmuE/b7OPPVWXXAXqoJUiFZmUH+zmUgJntsh8MJxQcDmCb9n
LfwvO2pYT/tIAZ8JtrCODfUduhYWF8nwkClpTL2VzJ/rTf+FaiuOayd2ry9dtPTF0p68b28a/Wu4
drbc/64FE7lJuM4dCZJqF0qhR1+EolsWABCmwQ7XBTaKlmOeNgUxMM1OSuIRPonLvwrVLg51xoxe
eOugVfUJxftCl+8PzOOVDMXJM0gtT+FHaK73nvjomtLXmt2QG57EIeCZnF8R9i/iosct/OVMUd4r
AmsC/SyFBOuX2xsN/1hWsXqPeHflWhx3kM9bGwifuImXMiaqh/+V0xtyNIVwIzDsqYkMD3Q/dGB6
0g7Mhy7fTy55EYamz/cHs2mlEt5q6QBQFKc5EqVl48gOnZuNBnAJNfybL7WmRbpBG48+LVn3SJ9x
9KBiAxUfg1MEkMPoC3PIyccGuS5eLu1kwrKfIVKyGP99ASThJoJ5rEbeENDtvGBQozaeyaOVUpEo
Hhm0WNMSYW8vdX9Atmq/BeTSEO+GLFRkKe5Dhni8967yEpL57kTdCz69A+KlNyKLfxLZbciXQ9WU
W6hYrGoyJeA/bYf9DT+R8jQmjQNQW1ghKMmtLNbDOyCIcLotP+chxWK0SL9NJnHomwkDIr0m+VFR
DpnpekPrCJH4LLJ4WuGcoUQJY1pxqBIPxEuKXZpnoHEi/T8vae6G0c0k4aEu9Wf6BzyLxMsJzjBn
rB4PX8skphQDftfOcC01cK0ya9USnh7HKrf7V30YmOLaftaWE/bqQRnNTHm5KwuNDCZ8Lh4SuEu7
5iYI+v2ECd+OJ6HjFnoJ7h8LlvSZy2324IjwDHh69dIISTztzPaZk24vDjCgyzXbG3fol+jeyplA
EDITQC1EFRaMWf8iX8QIqcpGHePg0yFXk20ut4lZMtuwSo020h9wQ04enJTH1PkhaqiD9yxNhQWw
493e14O02DHUCKDEWErK7dTJ7P0fu0uMXOv2Uhh3TnREAlDFkJE5um6h+aVneUjIcHXm/gQL0HY2
O1PsZ/ydgitxuVrgAHElGQ73DKCweoBtZS5PcWZSZuth/t6pn4T/HRN4aSS+lbhBNjQELM5r1y7B
LYyoYljtJKEaSgVQY9XMmpTs+iU5uKEXYPQ3fptBycF0w5eC8/FmrCVt2r72YYXiWSS87CS4L3LL
TSptUkvEJDVq4OEwaMxSTFQpGTcmD+gDXOCcA9g9rFFWlhBg8PCbxxwwCAReoJj44BRwi/YhCkE0
oQSS9DiAVUiEw1zBLmPlZb2xzUrl8zjIra5k2i0IF16R+Uf+FXwUAEdgj18SOKbHIfxhT43BD6ZL
s5PV4iS59oPiPaXwfbp4LuttB0IIuAY9awtRrLPwCP/cc32kbKhxhX84GKT8cSQSyGLISGzFyX83
DuxhQTiAiOteuY1G1B6HizN1oWyledXm+BAuWFgIdGsggLxlt01cG/gIvmTn9mBnkwwtd0nWTZQK
wrUPZHgKW+mTcY4P/HFG9/FX+6EQ3JRHRo3pfNF/q8oDN5uKoqITg3DeuPIYFbXi+p+FXN5GZlXv
ry4GqbQ0+FDem1hgbpRWc6ULJQIPlgXr43OeAwcH1G3YisBcIFtLzgSeuMHa0b4uXwSqax2MO1Lu
FFUDr8ydC2HmdveVo3vqQno8C/U2H+eIPL2hVCrbw6bncSvUK5LpRIh6CefT0GaHSvd80H0gFyZQ
NJOueZzSwpeSV/osRM2F0n07dqLTuCRmbjnHgbfv1wPJvbWt8m4UjhXgvbdyl9lDPewSUoCAjy2O
FrfeS8AaAQJXOq9KE8NkKHKZpj7borQjFgXYtHK7cj2UttSrObw3w4WwUDGt+mSKqx84IcSq9COa
915gG/xzd0USHR/ZkRi/mvm5WxzDzavwTtzb26raWJb2yNqETpOfZNHuj9iT6AO2ky9U/+4hMVM8
rgm6rfC0z5vOPVCK0SeKKe/9NLnErTRwsevIUVU7LBYII6ECRE84mUTMxFcX713a2Ky+S7AWwgs+
l2UJj4Umvj1m1HANjVsqaPY6hQEC31ttgMQYyc5+AoETBXzhcf6zeqd2ngxyHmrN+DiYBZxH8vSJ
fDddyoqGdriAJ4PEIixCvSy8jHClrhNd2KlczUD1Iu0NAJnIgWkwAYJlr5VzUsO6LrZtVHYpaIVq
ZC93heYSY1ohOr+gS9Qd2//9669VeRJu3PZa2MdSmpPd4Oc5p7wmthdBYq9FX/6IPOADUSZ9NqNO
7zjgdKCTUI+7ScmFkUGV690CHxBQfT1j4PH6dQCP5Ul7a+5T2K9JdheT0NXhrV2hn+JWYhEwjQaK
7wYJgnaWx/j3gfFCTXoVjjIf2aE6ZnF3vOld4EON1met+EUecqdndZ8SQXz3difN3ghWwSeh7B+o
0VuD8LyUISl+xnF/XRyxtI8Fg05UYtgAP0KmuhnHiuragvXE9izDGqe/ogfkw27jahBIXwpy6dew
i8SflQNqXyLVrdpW8ij8/JldtX1+CYZVZ42Juolnp2frIRszrlvntOkzDCX+IHWGpiefX9bQGJTr
/+4MIgiiIQN5KmbelSnjwS0JT4ZiYzll0H3UaSuhgeEjLAd0dxDXcUt9rIlfUD8Scw6+87j+p4ES
vTJsJQWOo1U+BKECCOOsjCUBLmXOAqZcwgV7WCpAbj6JjQ61fVBm1ZHoYUCszBmaFYpSREIUeVTU
1MCVlvaMF6PeU311wrpM3WF1UJ2JMSHK7/YFMQYdt8OMZcyVVbD+zzoikz+XhK8hanoNDoflqmiK
HU9iFpnvulA5SIdvuiSr3IHZXoQWjI3HGnLnKEFeRnB5JfkDj17m5Y3NtNV3e6Af5rdAz+HtwIa3
kG9dVyNCiWyyb9z/Yu5UjU7VpZZsTyUvpqB5U6G2zVNeWrUu/IDvfdlg+uP4XO/OvqA+6rRGocfd
lvqUDdYtnUGGcek5r7BfHv9T/+Q35wgQKOsZRjhf0zZuHilrMUH3c6aG8gKm/y5zTLYvbp443DkS
RQ1fJWL2EgpTzbU3dyDrm4sy59ylnma0AtVauIbcKu7k8Q1Hqk7lGlG+puDosG5avie6UwI6nwKO
PErNZ8UVGcN57cVbRTHrBQVS+sqF4FSJgZhTEMbGWcJLyBcHRFX+cG44oSjO3T60F4K0hqyNRspO
3kcdTo5axzL0jqZ1pyLGgxjDZiCwp2XGIFN1xCSzXPd2SKYCV3xegMUuPSWkcweW0SIJtZsdS//z
xyMBwNpPTQ+u9PAhHmh3ymZs7fi9j9tXB3fOipvRbF/Tl+ygqfTLqmji8nDEEE27x+IF6WnlGgbe
wd5iK45KY/UHij8fBd7TE3pA2z4erF9Kq1Si1NJxSk3xbjneUAunVraqIEkLDsB5BIB40GSqSoxV
4v8YuX+sFfaEau0ObJ4ruRveWVDbIIOiou/hGp0sZgkAWxxxp5Fzjw3jb4YJ8OLED+yvVMJRmCru
vi+salPZDVzBpb2ICjbLFtXomcu8BNjpZXlpYMv4cDgjoi2OO0vRsLOlG9D3h1BkhrrP1rMAs3e2
B2HEkUbhieTAsxrUkywkqBe+FzR9bEN9x/OR0nhUstnF9H9mGCP0gFe7JU3/Hz50jusK3kdK7obs
Hdx1l+EOkMDIP/SLRCeYRs9840ZBluiCZOC0PP8kXejhi9kH55SKbylYOSl6gQWEl2OQcy9aMao1
AWsE+kdJrxlxQIJEdTHIUmeoOBnkc0vUu+F3+i4j9at/E+7Ytr8sHiixMEmMH3A4dcG6mLVw+OyN
7I2LbFo1WGF8gLhLT077mTm8dYMkuZsL2ag38rShdde3q6uus/bKuvTkHqf8aKBBPpVWTDIeOk80
dUI5UFrOwMHOsTuGy69ivWiiptTV1Qo+BHDgHYHCdT/wUhUtrkApzos9za1KRX2CqUFIO8Ke/Dhc
0cIzMZVjz9+Qm8E0RjWnQl31Pl80htnVD8pq0/dZnwtqdjtxuVzEKTTGltLPD5O6flSrW1SopIAo
Ok1KZ1Uf4N1z0O109rllf403e0GHUautN4cpv0NOdBHhkIj7cFaP0gMuI4wtCX2erazxjRBECDDm
zebiPUunwwwdgpoT48GYgTWkMj3F5lMg1sTDZh1bf8a3Xfchl5NtP3dpI+rRGSt5tDuBhLABRKPj
wn/9UyUYCCVFKmXlatogKUO6gOtlbul/GRH0/X64MtRmqJATKPyZPUztaSsVSYx/XHGKNriLlH42
Ohlg437JAiLkFsdor0niSjQCrLLkp2rUJgzy1NI9YMPuZhHs0CwFPb+xx2rhd5WMw8clDKJS1IYt
X7qTp0VRh1ZQd6vD/3XaaGlyrAlGjErTUtpXG3K4G/EELiX6BiKjMeo6AzUVkxtJcUqoEyDe1+x2
RRtTwqbz1MgLxHguyRsSN0cxd+cj1XQ8+PGaysTmK3EvkWAWtCG9V5EsOW4K8mQAdRXaLECHoO3N
UOAFdP9VIb4QloRZRbs2KBeoph3IvkyNm1QdoFufbqneiBtjRwRRngb3/VFlvj5R3qWdtTsmIkfV
U7iz+GiAeMnofjx452bP0zJdadHLeHpY08rnfpN3eHqYqmzUeVLuNlq3Ry22ZJGyDRp5aiVZAweo
96F+8i9jGY5S/QJ54SGt9MuIfl4wWCoOYdcUvMyJqHinRUCP3Umu+lOH4kONiYCN8K8ZkyvCcFCb
FMejS9WDvXqbp4hNk8Usc29pHhxVwdcx8qqmlVUi1a0l3M3gJ+IbBGm1D9tuEoZmPXJpeHix+jID
huG0ZDlMLSzs+RXKPZchSttdld2k/jOpswpF/hRxsd3N93WIWSRT4tmuWzRY7oO+kWhRS6h7aedq
HymVh7A+gjGx/AUoacyyPDl0HDIu9tZ0IuoOy6FdDY+WSBVLKOMFYRlFymZZ6Wwdld5hUccxCxcr
dhaGXwF5PHSU1T+uEIqMHREK1PgqG9UlFKX1VnUXvNe8R0RPLGT2smWXCyo7WEdezRq0gJ3Sniy4
O2GMrl9IGdGRzwe9jvXVqbXdPvz3Yjm/UiynZ+jwBSU08ZVpQtb23EFQ9uLGODtYV4KSAi4RQyuv
bDPCTAoIEgl+BshZwT5CuZs02aDjS+/n5bi5IbpwW9pBe4vf6Jjgktoofwjapgd2YH7sVUdHcgY/
SkAYifYmRWfeBzjWMbkeBKCOKZWJFIxSc15lCEjPUP+BsE6SQMR2Gw138lv3mYcp6cHRfmPR2WcS
UYTZYRwLrmeGbbxA229NkV7/TE9MRMMjswXSL5iMXJio8WqMlZw/ivj6b/+IdKdNjT5tx3Yo74nq
KGP5OcbR3ME86OEswVaRKhWzCGW4Gbw9+YXIp/18xPKk6jzFRq5fn3YyqYreVJOYB8riyUeHtTcg
CT5ZkRpzi3LLB25MYCkeIBoHgq5nUaHX1OdoUkgV7FmQif50md5Tzg+RqBN/+LynV8FDRnVq5wmF
95kGDJmHOj4ldicRKHCcw3tpbpGovCtrEwrm4NgMLB+8v2LuzD+a2oAQlrwt0XREsFCnm4eE5Mu9
9RurCkR+Rgy7pQ2A6gaNuXgzMxodU7SwxRpduVUkuqsQgGDrQU8aCXrhdOa6lbOC44Zprm67YQ8D
hWFx0KGfkdY2KSe49rwgQYzCyF5FejzMPTIJYYQjV94ltiuDObPYM4N0BrTcRopi6H+3FRw56Lg/
IChOSIGQWCChJ9oqAjsTHITuAdwNAm7oTC3AaN+HnekyQ/8AYPSYAaTOmXBeJfcQf/O25qRyWSEN
52/owtz0kxt/PeIjwZPm7GpoN+inbJ1triHaxmRvuf2ASDbWLQYtA7oXU5Ur5DBe/plGy7pRRMT3
VCk77OyUF6csqiUg0p2H3ll0FCc1cUtcrGslAevqgmYXhN3L4ngu03+34R4zGW0cvpuqlWMX4Mwp
FSXa9TPeiPZwFGGKkudXiLJzyCoCqMV3CaBVLkuwzqTZkuwC5Wre79S30qAOmlHfWvAr/GtyEmyM
zrdxmT8RpBWY8ZSi+TowcBJxxMJPJt1hqsnhEe9iRbp7/STShQ1Td5GPodTsnjoJn27uGwjarZfU
bWMW3m9LT+nz1afJ6GDmpGWAE3buytDfxw5eAuoZxT7FGbE40siTcgpy7ZRKgx1E2vg6PfO/Jvz/
geKPlSbnkpVJW4MOJDhL7prmzU4/GkkrKzUvHrDzUjgUTBG9KUJK5KbK9dQCUjeakYtwdeEg1/gb
sKHZ9OEIG/YMpt4Pvm/Z/3wMPSBi15Qzs9MHunZ935So1naGn3nQG6RmJMAa/4sVXOSFvZ7y3QTY
rCVTWhTr0Zwsvlyrt8QAPaKf+9d53upVilK0KCq20TVLT3f+ScrP35dS4DU9ZFtNM3WR9/cDCq41
LJo0e6ccgS69KrY6mOxgagJoYnIbkNeR8q6IvHNlsbWkFd20xlwmBiNlwWcKHmPPC8eCVQINZ8CJ
/bcfkJzitlzo1x0WJ07SYEEwOy8njpISAF9PBMEWU9aSQkmXfu3bjLUYuhR+UtrWO39tcUIGVAb1
nOrQhvqnsVG9D0Qbxz+Xh48PENP/8JefxK1EseOya9OIhVLVOCycCD8zhrSDAHzwchqWjE8/ynL8
zkED9z+sa4+vCntnXxrgs/TdpaP4nyP1bWKlriqFp/jU5YTPItJKy33qYk63iCv/I/gPQEZ2FQyJ
G21mS3fQ0vpTu84vuOrXoiU+wN5xzybDmWgApcmF+Njg4+pDnm6DdfKk81iA0sseGItfZ8TtauNc
POsrC/3ABK8vQIE6HqnIsmGyJvml1yCIB2DU4eFpO0sjH/HWX43WLfzSfw9l6VswIYQeUL7AanTg
VZmNB5wWXSswXiW1LPU1ZbP7QV3YWWOPi3NTFqC1/l4jdOufEd7B6PYg2Ft0pHgpDYZBrjZHd3J4
TZxHbFv2MOWjh9OdJgqvHukIxS1X4q7Xyz4fRBcgSEwb7i63rnWoDV2SCHQFm6bIYAHMmCrWjGF+
nRgr8ny1ivZaJIUoYTEn1SGMkuSQkLYHD6dUaAeG97TYokU8IcBYiF87BFLMv7rUeR9eSb4T+8kA
uhecrzH+fgQDHLkfXI/sI0L3OOynhYfj1EoMIXCa+RvUiddGRWrs/LCj/qWrBtOM07+iBL96Y/0F
ViD9QEh4hBDQHGKAUqZa6/FFqXc0ZR+8KkliZmlxj2kF3llAw1U/LeqY9zqWOAPBCrbAZYer5Kxm
KEDcoyZZJNBcT8rXkWSydqNDQ5K+Yy60T0b0JLJKDrQrLCaVdiJOeiInlxlb+4OrWWShO+WMdh7C
Oi3Ltw0Q/gD2qYJ09nhl7u892I2/IceCtFaGWmAsPtj9Hi/83ZvtpSLA8YI8SX9y1V5M2tTIbsi4
eVhWxbVbxi6+eMDUB8K7DjOHzlwxujnydQqU4CgIWlbzMrvVR6JqhgWqzwinqoxa0wuwn46UMuqJ
DIGClGHVG5IL5r8hRAP57qsmXAud0+jHXZYnTVpuq4Zq54DDSMkaViN381jepnVzUw598yX02LG7
STiOkmfehvEjvX58DX+ur250M8Y2dD8SIgg1kq3Maj2cukHMTSLravCycxvWftsOXLOfnsSMJ31Q
kI9T4rug4oRo+2qa+0ZkVMTTrVKm1+yhoXxBMX0NpzUgu5wMR5Ie3W3raiy0fBuxl7NJsHMMYpeU
VmrsefexgA1PejU6gonRAy7aVyV7e0ya4kQGqTljyTMoyw6MUnatMg+uqxJXi+4nzo+SglZuCTkP
cy4Z49viF87g3b8LUxnbM9IcEATkOY03g3vhEsSy7qBMjHEq7O3dtY5GMAMN8YFVzMu5zaCa/NtC
rO5JbelT0OL9prl1V1N9jyZZaA6EY+kd3nhzM6GcBzVG9YleVvkQAtTNALt0QU32BJT9IkxqgxeP
ibKTP3/WuvgJ/KbT9fp0hEcME0KU43dREHjagLv4qVFOUaCZoF8B/Ox4YX4kw20egjgNSTGt9MVN
Eil4E2eRGNLK3Ii8LRbrBt4xGr1l1vOS9AsweqnWPWntHoxBvv9jYygbZByq48EAqmuIlvsrCvKS
2MF6RA5orixzRsNQ4Zcd1ejHZ7Jwc9jd8cj3bDo9UHV7Fgu5mnkWRvsCLlZTs0AcQyLPm2ciWY7x
3Y6J1Qhi2E9YlA0oAgUwrz2fSK8AAv46zbignuFu8Qqg4AT1QZp272yE2OztH/711LtnjAOwHcfq
jf4BLVZLO8BawZBZ/UOdjnkV/R+Bg8Btn6vqapqdKUusDasHtyYnyGVqPz/l+GL6GWG61aj9Ilgt
ewSHigZ4WeKbKlDDpU17gSXpY+RLwRQ4c66lQ7GpWzVr0G0IQdvGrxbzGm0UBKpWlm+ew+VlWqLk
ud6hj3LkO9kz9PgxqAaJvGrdjUF0CKV98ENLS/cC6SVr8DFGkg51s2y6A/A8tR/28w8UU3xWIhpB
Uryl0fyRgq7Em/5uX5adt8mBft+Q1AvsK+sDs4HidPjKsQskJzxXS3euldrkitqY7zG4FH8x0R0e
Fho+6YLhrnvEV20OH1JLP6+PiyKsbnS59DGGUTEtfwaOkIJ6b6HnPo9j5QnTeJeDvx2nE0kcDzkq
LmofbnJC7vHEKDLfltvu4lrE/p/lhWVXK4UbSRwUNCqyWdap+YoOd+811IcQw5COcVukDYOHlkZj
GowiSSxWemrcSUuDTe7j9sTCl2Q+X4KsQf60upju/ZBB8EHxBxhjkfKItmGBeCE/ZyZa6i8bJtsU
hOvpf9tx8q/WMjSPVmoAvNtZoVuvj4mD6z3zACiNPBs0b74kVaCo0oW/L4ig1THcIkFVb9BfmtxN
LoRDNat/5U3QBuPklUkJj5cICE7pADuNtDJAvAkckqw9aEYiRx9v7KIWYuv+QBODIKTs90tOndiG
QgLb5tcNrlylL6bk5+8t4HOCPgZMGB2Kv9fiHk6MndnoX6am/KRyrfTHBjFpqNiiiHObsypdw4WW
OfnLB2aKCGeMfSSNl/miXccfp4lulwwKPSfciZ8WYF7r+EtDxPQBKMbbrKCDN3WUOs2gArzE5zK5
CkE0FlgrwuvKYIxr2gXEWj3MeWkuoLZYeEK1RchxayUsKDDgf4ZafFaaFzGnCn/ushwlo0xMLeyZ
TN1IdsMCuOgOFbj1zFrkYeSRFS4e3ysC+o//F3T7IGeadJXEa6iI83PchXadKGoyC99jYORpZxXj
wQep2BuX1teYqYba9CIOHPwb4srcsQp3XWHcEqFxtuaWSumPqVI+uVX9nsp5BrQcZdP2u+bdu1a0
oAgKl/2dYHWMMl9v5YiUTvJaXnE/yPvnKLBzaduErY6r0pDt/J/nBdWRHHKV5J4SAr5O5g3dmeyb
lDnI0QO8uzCu2fcM8ETK7AL/HYuBH1Cz0ilgn1WhkYdkNm7xvxKP+DJ0TqMhClozT09NbfBOVPzC
nZnx+N+nCjJr5dreqKSaMfP+Fu48LDy8GckVDLLqfXZcu+eetSAizUoWQ/T1uNUgafjxvRVWJOCS
QRxC1oIWOSkYSjVUAnucfFZoOKFvbWUKIa5iDRM11ZIvW5jyWoqPT6yzK5OD1PYKotUs8FIBwPo3
z9Yu4un8d3Cnr3desDXaHcba3HiFSBKTqvzgWHo41VLMjt3UwwO5k+7Vs8P0xrHaJOLYUPtM8+ZI
EkRKItkidlsaKYs1m/rDdHDYcKYL1fl7t0gP56e4Fg6yIansWYmOjzbWVzUjPt7JLkHGOHV1uygR
LqcI5YIJr7fQWA5/vuIkB5Sdt+32OKSl8iONgTI5QkmC6l2lNiWZZXnG9J1aqIg+wHmajtG3aX6u
LDpoZiM58cYPQONroS6gg5byyCYMh3D/Mgc7iY7vJ5tHKhmt3eVW77I8s9dqhSEknxdK/YJkAlze
V2mEct/7nF7XCuVU3LMYq3hPBvegFQZF7j1KqQyzRbJ3mM6tfPJgMAMKDcYMkaD3ZwlDvB8K3qoN
NSt7MvIg4o7Ql33Bq1cyPIi2F53JOAIjqnwV/ZluPC+/CHn01XYuhAVKRd6vmYYusyVXlKnHLrqE
gPQg1Rqj/kCM8puhE+Ki0JCWXNmQInGJUh8D8UKdVJQwcon0FP0zTnImOYiZL5N6Mw3StRoaKZ6w
Xhza02dIkJfoIlDipf7DXi0asNh8r1oigMKFRT1SIdOGVR9YQ1PyprstqXF4RB/5ghBxbM+nTKHB
BtL6cPFDl9Z1uGrczJC1tyaWNkLGN8Te51At877/W/jaL0abFqTBD38C88eyq0RN1A56GS5th7+/
6T14IylnZT2aLIHdV2S/4LFXzI0Gasj98nCps3H9th1VoXm5El1q8Cy5OuD9zBB0f9voQ5EZ0Es1
DeKSXB+3aspQ9Bt8+pbeH1Sr2uxT8qBuDDJUB+zl5zhTPZMQA+81xluudwasLOFZGGo7eT29qfZn
l6kiR1gBLJnENV8l78G3USw1lCqD1gqVOj9NaOCtZNrzsh8nAMNZx3cxM7Gdh6W1tV8VYRRWYaD2
E+c3PcMaF/rfmxY438VRVU/UxhHeOrN3164RyR81Geto7dvE+u42yj/59DYpDQ3WU0mI9Z3ByYkU
GhbN+EF+fomV9QkFohSUepXkZPruH9tRg793THXRhTLv3rmJ3qaEsl+1MpncEMM/cNv44qbkCO+y
19t0C4/0veXmCJGlsAjPCQYbN5WQLN74lMdFOypwDdhcMfAlbLf4LaDjCdXNxr9eBdke8ONszTZ+
BjIu8PNSDXNRUNsPDVj095APEeZWOipyv06D/LjnM/G4fOxT1zC3rRorcvXlPeqjDpEOFzDLRmrs
Tx75C9yDmNVbkAq/EXB05Z4dlQlSLDm0HpbVZQp37t7l3QjlocxBG0SwUdwZk5imfAVIURK9+j/D
SAFAeTxt+k/oLXner1Q5wE2lzReTvITAZdp1m44dcqX+hL3WuiJbi4NPa2+gQYWS9cKqoG3O3sgG
XWKxIyPlnyyY8MawNB7Een8p6NTXOf9Hw3jV31/FYlD/AQmGLH55dZ24pNhp/yaedrqwlMbh8x9S
429zxPvymR6s1tfujsYCevOqqXHgJzTMAO0ma+UtGEtQtrxTPzylrObc9HAw7/f8dJqoo/2h4Mo4
h9PtpuidlexVc5GXG26JsY370sE7oOf4qPn+6DRjnb2mw9c3F10PxbdHDP6X8g1QZn3DmM5HBQ8A
ApZIkDIh2Izql+ye3oBPAZF5XVr6gt4ZMi6BCJ6ao/R8MinRbGSaLMTbPW3Dd5yhgDPU6BeKlTV3
psCDR2I7Fbqqv7AJnvJZLXXe2PDpiEjKrLnsaZJDgX49kcsCNHyUX1VY9it1is1CmjooQIwe5sNW
7J1ipYEXwNySbIsBG8Hosf6++R8FMKIvCMcNUjB/vcPog4pEknLHnMBLo4prr5JkmwI9Mna2uspY
Gu7OeRpyuRT/zjb7MK9POUGEaS/GjgfRknOPZ0hlw+9nXHWjkYgEK2qk9StXm3hKNOwBzZi1/za+
qIy0yEMtXc3Q7Z1mvjCj6C/OrTnxCNwxaEvtm4gFDiVE+GWY/K6cmBmhSUMqiV1uJnqgoKCdvmMx
u3spmgIwwbGLBEtOfUmrRvODizxUq+ALBEOwXIc3+v39zPH7tN82Ypjb1dx/IJHC359VWOiHxF0w
HqmiWI8njH4/a+76LnRjMusJKPGbCYZju1ShtC+9eHHphwMN51GAOhp8VhudCXw+Z2bZjISlnkRf
pnYC7o+bpCC2ZucGl4QMWqsgNy03SxrMEh0Q5xnBs9utlNiBXqT5VeI4rm+eUcpbUbQSiiCZZZ5Y
lSjuR/zQNx1UQ5rehZa4BNyb0Zt9QiYC9BXhQxXdSk4+681YNIYy7b+Sk9vb3q64ZaEN2Tk3u56D
KDY365z/zE1zVe4+aBDFLEEBBjCQ035ZSK8txCkp+9vBit+qx9ilK/OpWGjclj7JRHkygKfERFkT
qNGJC1KQHmRoZeVeaQV8NEW1Q9FXB6lqQ8QIeuvULTJAaUeimyFm7lcj7IfVqEg5g4e04bT9YjQD
+NtSpxQV0bC4BKsh7BDho+lJO7AlxppXLmfoo9bb1bIbDxgLT48M2pGzyYJED0ekQg/6E5M8D8za
Vl47tTW8eI88Dh6SZYT9aiUyxOGJmwHTIFHo7GeNpN8oMrpIkf2IJfuUxqcPm9GzrTThBvvAvhbX
3T/wjGUAlmo3e5eVwl3OPTfp/Cr7dljMfbnPrcsuXNGt1IG3+ICxjNG/BxiLwbRNeFkJj1ftOIEj
j9MKHBj1yAI68vhHHJZbHOH3LM/MNB/y9FLJ2GoKy/w0iAkPItgkAQQblGRjqanfK7ha+pdE7eYI
UjKnkXiwPdyoD8OV+LbR/XyVNwJdVQuu6s2MtmzpB2/zYtAbz1wT+KUm1OGqLPy2yBLdoxLYyPZI
t++ZBtp+11YQcTKDDODsQDiWGLUSePNEjtsq8K1IZYSLbxlRWd81o/zvxQ+yyZ1THMh7Wm0kOevC
GNWKdkxJJL+xsfSiKjFQrzKu4I1jZ8vatCJArwxaN3mBYI5g6WtVPal8Cazt45U8mhca9BQQ/p4h
SLX0+1Jd836zFBUHgiE8ZIt2d7uqL/A/Z5IhOXVGLRu7MVjD6gEyNuxcKAtKFHmGOowlV8gr+bso
daY/VMdEjMaEWB6GS+rdCVETgufv4mOK0AHGbLE77P0I0X1GA2nl1BC1bA+6ipIeH4znpV2lruqH
aNTlZ96KK6iUFJcBBO55kkxx0pIvnwv8LW6uehLPMbAUyvxYvmiq5Df6txz8ar3grA49ucIWslPn
QBg7dcYOFwzkZm/yVHP9pN+aYIF1Y2s1BZsTS90YKQg8nZLkeGt7YyC8gcOeZAhbCfFGBNIz9y4H
w2cepJbb3f3LJGwzu07dNZlVoTbKU+X/7M74HP1c9vf5V8jESFYrgCJW7P05kc3V1Mlxl5drxkte
LqA/L9667Al+ldCusp6BI/251jshLTuuPDzFuKVlYVLPvrLzdOBtT42GLASoE0TgxN+3UI95vbCV
UHXC2ODSh5OZP0l99hVnQiASR3UMi0jHDk4L7NyKzPBs/sUOGEwPK+COTVVdiG1XvwyTR3X2MxZo
THYRDblX6MhrbAbISBge5b2abP3mjFeamwZsEkdCynG+4R/tyG+jJScz1aFxF6pW6+HLHvmSaU5r
EE8X+Zfd4vuyWmu4+EzsXkzjxJacHfhUaCWjiSQQ2M4fotfJRjwqw7F0otl5/N+5MwsBsXr2iPGJ
M8W815T5cD9Cf9JJpKdQMHSjHX8d/NbHsAcYZvJJVV8n8pwUVQcLjYGSVvuafLuLNsl5MZgMFnzl
LXsqLM55w2fTi8EtFsarr6e87Ct8XCM3QFAAmkMiFXqST2AlM5t1DWrmtH+5WQHTbiuuwLx3CU7n
rtwBdCSWiBwvl37PhUYgcEykmabthZVFj+rSeVU4/bqLb3TdXHAP3TGlvkqtH18SZKTQWQC7wK7R
Hge7BKqIMUq15GBJ4P0qxmpVHm2JR0rMjXQAWZt0jD913TAD7thqNWfW66UfRfaWrEmsq8ySnk5h
7R0tu+OIbhSiy45MkxWJYWedXefcVmKHmtMf1FJb8bTVoqGPJkX6tMOCr6ytoCIj/x7g5AqNFjOG
drGvY4U/Mp9ZMPpfutwfXXBy9344RSd8Wy18HugBHC/HGi4d1qB2XJPRmRU2mH5ZofHNm0+d4f0+
fMxDx/lUnq5QiZcBKV+YKYkCYHPVIqwkSVfXK5ZzadvropFHtdspYBTsVtBQCOmk6oTLpNDHIzmL
qvaYadpNLrkWUJyTN5Y7ZJPzpOg7uluz5ytPcJsoLAzuCLL7k++WgK8En0jXe4XosmzxQg4T0GBe
H6lOyRteB9FP4dliLz+CWkeUIrVsxl4u8iWvpVVRe97mUk+5KeAe2NaVv+elBEY9UZ7xOBZioXve
W0SmjuqCzvAIh/IfB/PkRo3poLEyvCVwbCgqL1h037u7dBkeFvScbfiT3ji5iziukKnxcAmIEp8C
DMNyP1oG3CRJmB9podFqZ2ceA3jwZ92m4PNmH9pjDjqRVflKzqjRjtuEFVWO3tfxGj2h2EweFVrc
hTIXY80ackvP0GHSfQexoxPqnlDOcN1ckQRl/x8mh1LTMh9YfyqG0qgxKPiO8j5GD9AumweyHlc5
R1bvrdANCfFfF4yQZWo1aIf7sQZBLgK/MWJo7w4Y+c+6qVtgsCnAdC/ro49JSAoF88RL5Jsn0a0o
Fk0GtMfjXkTzCrCTsDwYYFzCbdfJz0ERw5YkvH6/NPhxjikWPRq5fTLneL3WneutWjTti0DVx87t
ChqSXXqlmnbJ0OvCIK4BroTtlIc1PyJqeSeQcvlJ2WfhG2ZQIW1/ocLbdAhZotSwQjeqJtjSVEsy
Pctlh2zdnuqIsdecGMoWG5unJWxQgXCkEBNHFFra+QtpySn9KTuobJfl24I83yShY2VeQrtI9gI4
4WvG95G1EIDUuaX1nJIlimaW+odRC5+vkGT7XmapNHqocaOCNkrmfbFEGI3HFZIWPUWF1wBGkQF0
0wIvQQhh7YTFHOgsJv3yM00pZPBlOi17Y+H8S4VxBxb7dZGPihtbtds9pNS30wpt6KyOz6cPLMod
7BcWmdid9Pfab5PGkDhh1PNVjpZph1GX2yw7CfzKosgbrmO3FBp+9mggjNj4ADNcK9T0z8d/zwdH
lud27MDnipHuuVfKlLNRiPLBf2qUgnYi6nHWBwNkJ/NLD2k8yt+Mrwe3gr3v1L9kzvNvu1af6XU9
/UvRNF1XdUep0Q3Ts/1AYxcj7VnQ5cYIqhM+xIpE0bsZb9O4cmJg9n8Qrxb5er8ECdrxTEcvucjN
UmLU4gog4/u2DuhAHrJY61/LEkKv4vC8oCCgiTBPiPqaQQuvhHXnZZ9fKpKCiKV7Ga0W3k820c9j
hBxJLc5B7eNz900coWxpKzoOUkAx8rYADwZQbbx/RkHsD00lQUr43oDDgPq4Fi2VccHBCanbLbSg
bZT7Bet+CqyQQZLXUCeDUg2F0LBSr1aslWIIfrMDEBBm/SIhF6Dj++Lta5MStW+sBzaM4hIptx2B
J/XS1WqeHeLpNu9nv/Q+OqCB+vxo99n6sH2HPy3+M7wKS6FRjEBWIkoj6X1VMqD8XPKaRQXRYjEO
bIrsJaDPVlY9XPwFgibKCYs2HIlpRU1kZB+u/9Fj/xjxzyrS6MfFu5+gr0n7GBo2ANU+yXwbJ+9r
watlehOANtFN1eOAmV878/CjzlTOu2L6MipBtDD6pFWfN6+ykE5PfouGK5von5d3rlVBH1Y3QRZ6
aVzK/EiBDaX8FWgvje2XPW/+AQxdjO33nHZe6SQnKnaHL8SMvcSbKy+NZGv3vf4r3hXJLBeZk8z5
jjosdil5XMTz05eTkydy5d9Bb/dswC9XFyzoVImZDzzFCGmrM3XK1oMlu2+Mc7mFZ3+/4648akju
yRwD8jfLQpOcovyqi1YuZXFiI6VrY6vF7PUzuxS0zi2W5hVejKwQmAO57xJbkZLg1EM2BTIqSbK7
v5MGm5VG3U0Sf1eZbRdktpqvbPPILbI2v3FpQeC9WA9eJGNlbBOtDGjOVExSg3FTKLh2POMiUFjY
PTIzAJRvcotOC7EN/ACCNp1ZdHO/7cHgjet8gNQENdFzTSvAbiLvALY5MOTkaaNalZrWdGW5JH4X
TWUs5j2ggNL/3AokiACAxDnDvDsHCFMXQB71Xm/BGPyWMveuWZmjnlsmLD4gV9KYwHe+UVmqYquq
RgRQRHXnpNwCuzE7lS6M9I/xwZ45fmjq5NySctn9vKe29VC81zxpM2lWvYuUOfTygeFQ1SGmFPEj
P2rmZSE293retyYxEYcpu0i4ZZDODRLQHExoctLeL2uCMY5YZxfWYwcc3dFGxegYlNXMFr28RZtn
MpZ3Af9nWx2M3hXojYPxfg2R+TL/2a/eOwIa/SvI59tuGvUtn5lW9DUXnI+2Aw8dJiHE46yWzZKA
9wpOaZMJYwGYm39DTPcZ63A3fE8spzRuYtAxGAevt56HHQrB3DJx/a9sQEdFtPsJwssaVjq3Bcww
gX0SyUkgokF66Oa4pzh2fDnsThkw088p3+o8MR+xXuKMs6RawXbiR2zwUa2WKzdbf5cRBFtT1xn1
dAmf0AHvQTVBkbidQEiMbHIrPXz6p3DRw83X5bA2Swa8wul9SLKz3+KG0DUDn73HcqIl2CodpkJA
XrzBdf5FtOka0SsdcyFxKKbyKOSFH6V69unvB3Og9UKRYVupb2XGY/My6sM+J8uw3DeqMKFhh3NI
hyGH5oVF8KwTQBaKVTov7TWHjJFIsUNNAd24Rwz5Wy1hb3JJpOyseXDNCtseuEe2Pao7hgjsXOn9
f0SWYbXTyvoVoIeB6CJTfbXY/oBf37G3Tcm9EvyMY4rHf3M1P/5nWTuA5HLHfOcEe6JblEVaG+Bi
QU2KPd+XnABBg1CjoOZ6RhlYE6byGME/eRP2qyskfkCwzqNSL0Fa3T+Vy1TrwbUVkwSxtki/RWPY
P5aYvLegJFo1L2yqCm0Pw8XTKXO1NnHNT/8Kyn6UWIW80EkqZsEJxXFrS0mVn4FZaGBK65AFkOO6
/cKdjvdzNUyjfwsAdST99uQY3PLbt1gr4c/uXzgVuNhh87gxHClLvEfH69ra3BPIq6hAxdrgHp+0
9KcrpL9kt/YdaPhDpyYzlXIcuoFkZFLlF63jHM6BHajgsyE/1eBdReHWTxds/gA1k/5T7y4d39xp
Vd7cekEQChT8RMYWp5xTgD0VCTz4lU2fUOlnyxUWnYdvqPVYm2BaW2w5imOrFIv8UNb4mEhwa//c
AJIp0MzgOoEqiRXTjMZbYbXxVJwdHePCrsK+s1E5Mu56sivmLLbmlzoIMoDntpEzVf9InCBYmO1i
TvgVZRAgYX8aTnGOJiVf4bkdqFpIxzGtXy6qk9TxTpW9Fmh9YUNeFstv//m2md/Dp0KJC5UPP39b
SpcDeFGUBdzndY7OyBacKqY5wFHH3JWzFVDwXN07mmKCbIZBkRxC0ttigCEJhXMj7AS6PHudOQVa
q9n2w4/sRKqn7PybSaN0yb/MXmg+tYqkjff3lknaEpzVfkxtRc8smrkobvZCALNmFNOFhHsVYBA1
0QU0Wq3RhRkVDhD1tHsfUEHz8UhPIrbuFpveveIeeoY9ooTG3BiAAIyyhLf+6Dgo30MEJBaPriHU
MlrNI0HekN+Fx0MW040Ze7Id10WRkh7DCRrFsORQpMvQ+yGaENOXK8iXfeiB9N1x+5ocVjo408sQ
87xvfdXPxFwdtiEeT+WxRAC7Y4rT0QrobrNs0QgziFhDPcDzlvBdbSlCmxwT2AlE0e9AJU2eDo87
PX17b2YZ2/zRPehaxVH5TuOjVlPhhxqn09RkLN4MmAYH9YaN7pkbiIgOAk1VXnqnGx0bAgnh/8vt
DoqRQL64JoQnMVOm5d4z9EsY5rvYB7YcePjl49pyDYCHF42p97DmbZPWHyMQhnTbVK9p1XiKjjwy
28FgYSoI5iQWqxytvSNCXMYWkFI951BUJ5s+1P4fLDveIA8ad07s5ImEIYJ8S3GMD0nP8Isepidc
JE8qvxsUFZ4+QGfaQsOiD6yjTFJRecEjhqJJIGFqznAwML1WHMyFWH7U83oumQYw2TMPUZRcVKZX
2B157HGPmQQICbPAUkwsS0IMk+ZYH141q8TQmS5uJgD23kihDVYnMLrygCZVJ4dHFwB/gPUnNduC
umdjm2x+7mY7PEfoP7zmRU72NCK/1kHHGieRLUh+aQaL1pAXBdDHC8xqSTQtEEoRkglnMnWvLtkN
RfnK/ddJuM42Xm57ADqjNa4Y1nSHaMWvhL85wqamCQNZ7bFineXOWbb6Bu368wjiRGyLzI210ZSV
ws6jt3DzkGutCL3pFGAR0Zg+tNT/R2gOzNwxDZEYse6DDDL2t2Z83UrnUu/bvENq7tWUTm02dRC5
QGNS9kTd34PFf1vPcVYBmAi9/2ulvyCBr1DePdU1qSefKbgBygl08VBwToHij4pSg/TqApkhGFlz
mdz5RMuSz1hSlfttrVIIDzmMtxU5JIv+pDDMRyTSD/9KfBSxGcI4DbJLHfpadV79yDDTfwYM0lnb
z7P3q9xkvr32oYpZtrXYGIgQisDwfjDWu8J3u+K63KLt4FWtFazdEzhEtPFB6A/aVOQRLjYyfU4A
QMaCeu5VLFWANRnS4/zeYb4klP+/RxymllEZPSecVey0O+8KpmwU1u8H56W35rkvUVXRBb93rEPv
LFDIV0Gjb6gfCSlPtpjbOsfgrvmROIKi7qt/yhymp5ZeaxzRAuL3QPGE+rAXcih9BPwRD/222/bM
E/7g5dhZP7/VbIyY++I9j+yCXdZGVipC6Jfc8sS+jLdJf1HPl5kg8Dzb2Gx+Vyfh+uwnHA2p9YLw
vlLk1MVKLDq0NZDuG0bSQqFxWMI91blAEvPHgVlQIJ0aWrm2FFeZXk8fgrg1tCxmfnhjuvTzX4+5
zkseYoUozSqIUAKiaJfdiQ0P6cvSvsQAlYgv6jYGSWUbuMpHGhGTKUSC4MkFpgcoXFyu6axYKr+B
cCpweyaixo16UQ/4VC+7BO65NF4pq//rs5w8IAfK9nq3I00AmC/TyDsxOM25P4+YRH5Kw3fyGHcG
Gz9HMUKA/VBPoug+xVjK+HGSrQ4vdh3jfKf+rVAL6JX/VoOFTdfo5YelfvPTIblqoVW9rrrj8dLn
pBpq27DXiqG7sz7k+XEBfbb2YqES+4K5L6zmMgyaGLgTGAscnv2eDKd4txt2FpMnyZ3T9ZCF8+vK
6CAIU4C4JLqTt5DG6J7u5JGlFdVdaH4RighkY4Hf4GzRFu9jDiNSNVcArZAFM6Oy4Y1fggs+rs90
9rba3Wmj53e4Os9Wl+Ja/gqiN6rRxNye7CHT+axBv8N6QmWLCnUInsPBnVGYW8IWT/hpljovmQW8
FnPn0dwfr5qeg56VSBAiuFDHz9peeiXz1QV7TotFAZLW0t3hx55GeMvhiMDCaYb/bQArl3E7M2g5
Yhblor3Giu2nlIZ9vCLhaqLyXg6Gyw64WzY0OSbo6wkhKug051ZXzQVNViZqtTiF7Vz2em4gXx2m
hIBJkBSRdrrHAIWSFJpyteaMAoIbJGcs8otgM4b2NpX3ljplHfMGDk/I1IVp7MLtdcMHOcxQ/0sn
u2+Ck9UzESj/BE4bn6sTpAlgOUt789MeO1Mh4dThGBZh7Oy0ADau8ky0Tg+NbctVfEhhUQXrWeE2
t+0KBFsrtXHCZhL7G0zhmCLILk45CU/Wn8uj26YlEb00DbOssuLwVCN8LzKS/79F5oJOKjgxZtFk
4bW5WRpFlNugjkT9walY3AzV+ISB1UegarJk5o3xkC+Zx6y+532FmkIXiJOvnyizwKXebwGGkdmz
LGja9aQTNNNp1e1iqZnKxdhZDKBZaOVHeJ3w+B8v1glNG3VnJDZAlnQ106/smaImzdj7G1Ek6Drg
Y2rDlVJ6/48frYsYnnsLKpJa05L0RrhS8nCnGuLJEnDEy0V/uG9AIIoywfQ3kOcITfDM/d4+xeGb
yeSr2Rs3uHl0NpW0AhQSN4HcCnsLyL1ctpqRiM0+ycjUHK9ZDzGjc4zvsefTsrqIOeQ5+6ATnta6
+kGvh/S2Mb7KVyrd7GZrLde6nET9PWm1lAx1kLcfuoloEnkcNFzyN7XsY+tGAy+4ibg/syTPr4Wa
bYfyasuVzYerd9b9qjj4BATnN3K1ZaUUjDgsEfYJX+Q05c4vRovZDQIZvHVsNN4ZUaNNRJZ/SQNM
bJkxItouOy34W/TuIf2OHBYUmdCC8iWtPXl9NUq2jtHucKenfayr5Q2khqo3weDqFgAQ5pRg5fwJ
vTRTro+xLnlZtf7QHMvntVhrZhYt83RAswQ0j/Rwo1xV92UN8TfezoSPST648TDEpZZBneCVVEYt
hNbU3++DWjSu4DfJuh2jAjTCJLKSo6GjzYB+127ddF5HeblzIshK4BLDDMaviN8QKN9no3ZT9WYR
Gp3UugUMAzzTbnDtXmQS4+Di14GOwZuPvOK79CDd8Yu9R7aVZ4zGBUwvx4ymGIOUxxINu4NYlF8+
zrHWEwC7g5XG/ctSnW6D27yJpR5+QuZRlwjWGJiqdfZpe3WSDizDRUxniqUu5DvCyaqr6pFATpqR
OQ4VvW8B095Uhm055G/3FQecFyCQiUJvjA7jTJOOtJ1GtNaYy/8QrXtWCYltFKAi/lmfERvOl+wE
Xv7ccUM/WXPOZNTZkjYq16Voh/77YldGiHRUWvt6NvK2i9YK86iTKYtyRAo7FaFMt2AW6h0FlKfH
2ZIrFGnGFNqCVLDL0+d/gOeztazftRQezXeafBhexFpCQ5jzJOfpJ/hxqqfzPvVPlENVoN+cL0M0
bVUGaRwIUrX/sN9QR7zqIdcmuwJQJYMxTmBBumaBgKSD9nYMoJ/kuwlBFFGtDLcWXNfC71nj7yZL
ZTz6EZOMFKx1aDhKY6ynYlBhm8fa7SoWLcJ65Vj7u+pC16RQv2SrgbXz0Rzla4tLeYnDFjaqJYFd
UagM69v99LfcPHTRaTclAZNK6jzlAMuHBO9FFxwPDPFr7A1DdYg4lAQ0oDITPDUTnc665QBnwFmn
9pVOnp374c7U/1bEjvxBITpN53X/yKjSqKN66EblfYHbwM/GLzBPVrD5ZyPHe6Vry47rCypwmUeU
QH71O9wSXzC+ZSFOF+BpfBXTD+Eb3YGt0koAWGT8jCy73VtW5rsYz5VS3iRqZ9t2BCU/pOIb1WZz
vk3pXS8uzn4psfQTenWFb2Q74s09xB2NA8YCuRlHVDQOZ1nNqIUxK7ZQNGbYxc26oMkOupfVrKMc
t1GKZPUqBe2gzLjFICUtMCZjLkDN0iFeji5fyRBzja4XG9iCpl81pzbWXuRBiMJiCgiyyu3235Ro
M3PpjMu6zHNvSPtrNys7otvrBc4fhks2uLXjBhsb0rtvHGoaNmftmTRtuQLA2++++idyjN+fVNRj
MADDvlYktRzH8KxD5rheWEjJ4Hlg57DcHCkcaWmjLUL1VgwDpartxB0yEUDgmCmPMm5vlF1NB7lr
JC1At5SOECO244naM2JibjJKGkNnZkUAuiXbuVPQF7DNoOJtcDPTFNI76GUueMGc1HSwdiio0vbS
c6ceZpFmcUtVN3VWndbmVUj/xrtt+LoX+5hcrD4Kdwrhoi/Lk3aCmDzD/mE4vMn1ERGW2d90XTwD
hFxW6M2W685yMGn59mAiGVQLnhdZrQvPASuseEhRHxtg7QS58XvfRVgDLrSi80CfPBcgG/Im6cSi
7jMqvH/ys4ukomyYqhoVRIWJRH9i+V0q/u8eK2J72vso3pfMoIsIo0Kqo/0eJ9Ort2O5BZb9JZby
e4mdcXmLHpqLMT0tW7vNrE0kEIgmy7kE1SfB8R2IsT/uwW7h1/BY0EhlBTty6dRyjXEClm4l3E5o
rWAOWvJ2Bhwh8vmAOgb6/fEXR7U9TK7XQohKein1kAWehBChKUSqX5zJvjHgPoXnh67N/ukja5Vr
YAgRg5UgWLxmmqp2Gf6Gz4N66iegb+Ns3jKnP4K0IRriww06le8AZ8Ra//4IDZ+9PT6ks9SP5pCi
f/fOtfwRctkEkqOouqcZTCnfmcFi7T1PJtrsKO60mSrZpyaxNr3hMARpeZ0A7fCmIIzl8jIcxjo+
3O1ifgk7i6aUETg0eR/xR0GcMOtjvJIOWw1+NLldb/TaOibWF6X91IXmh+DpUQf6z/fQmowp8x39
XHMguD9kFx8dOuDyacIBiirju8/Qtybo2YfVxaEiVvZUhzi2aoLE8aBijYFsuozb4bsTWIxRTqb4
/ZyH/0gawuGjxtKclzETRJBRrtRBE+ndrUtkYFkRaV8S/L+zlaGwKu+KBByvX580bNPrs02LTa/o
sOozREgWJrOiJo3baUKBKUydM6/6w+bqshOlz0JRCcmVwzChztBc/IC8cuUQfokIOiCV5CNqTvW/
9XCCd7wef2CQzSidZp+f9maR1WRrN5cjSiKjN/KqYrq3Ey5dlDJDc/Re0b+p98O0LvDsdH/6fbba
8RMUJW6J+OWbr4W2sGt4np/7/6eKe5BnmA52XhQNd8uD0en4V/4cGKoWfuR5/gQRy4WybNvF0B2z
l0SwDaw47C0p5vb3arRQU/9Rh44ktR2eQDXGAXs3777bsQ0RPpcErXt9c5Q0bqjsOdna4JDe22cB
uVZCcG0VC7UY8dI3YNS3GGRrqxQTSJp7yZcwk8DOUphVq/VGUcH864iUKAtB3YlUsHGoh9GTmOcX
oPMIIuaIMYOt1Gog4/tOehqZKBKUq4G2VawQZ/DizPkWpdn0SsnsjJ55M10Zd6f7lfM3fubFZbrM
KOxfbI6HgifLMkSEVCclEMY5UFIK4t2okvHkDoUmzCmH6zE7lxiRCzJ9OambGWq4MhL3ao8HN9l8
nca6Wr63d5y9+B7PF+4WiUi590SQlrZq30Nwg4GIuFsRh5hRu69O9KVrc9pDQdxAFGKP6Q8vkNgJ
LovNQ5SwZy06DmwFBQ2yINTwMY5H15zqUZ1scxv+MjWRjtt1uGnxG4ASAL4lb2EIU9xOGlIg6MRj
I46GJtveqzvV3FrnMN1dAtHRUm6FndY/Owu6nDlwqLj5DW3FpBjQqQoTchmvTfJoh5zJmMvG4i+x
vkfTfS1oa0b29W78Ih6hYuWtwhslBQ0QybfeFR3r+JtQBRNG7sFpTgvmsi5iTSVVYzamTss7ugfh
n47EVMVc8mNbKkBHGN88jbXoH+7I6w/D3GSDwCAXaMVVXykr6+tSuBeBjupFER7oZyisZt/G8adF
NgcxEN5ZRA49T3RiV52e+ar0F8EeBNWORgemYDA2LLorXDJIObiCxjKAkBS6ysmWlybUusNNtFgr
V0gQJ0y/TcUB0EMEWK6V0UbHyReDGgFqZ5oZFjb24/8/8bBHhVJ+6nCCRihDxk7Xw0X+h0OIN1UB
GNjgvaOoyLmoMOds88b2EPgXRW+4JM0QTHvfd+p+EHHblGmIn17cLlKaks6YPmJaNOTEYTBvHQth
HJFKJaNoerU8JAvGwZ69kmhHYpAr0hz0r9jUzLQANMi506qxSWpjG5rE+zvvmYyQUFBqGzsqCAcP
UDYYUmv8+mWFf1Wf7kcEEjj/gu4/ea5UXHq4m+qceKGvORGyA+/uKLq2yOJc+mgVbzGIWgH1t+7/
rQP4YSCi4y9T9XMI8VYuQCWtlOKXA3jl575PfMzPBXEvmZL5uBVVyQ/msLoAx6LkMIe2EPIdcL4D
YMXZoX0G6CdVESTNOxBBjGuGIPMIjc/zBnPPtk6GYMwdbhtwudd/LFPO1GRN722l7KpJqWS78W4y
U3WZPW9uPv5/8FgFaIl0YrDVAeM7/WX9r9smiR/UJ81Ty1K4rzowzs5SkOs5OaDv+2iYjZ5chlBS
OmQynIGG8IejnQ2IGQKE+SRRI4tvE96+wz691p+P9cDEZm/Injfigm/efUJzGtfIkQgR83RfE81O
1mU7OO4ZgVAyaPtLDqelTh2kl142mxDp+ytlee3E2p09kBDr710zS85c9AjiUZ3phVZo1w+cscL7
JdOgPFuus4NCWYxBPydbi9Tbqlno62ARMWizkc5kOHui7MNRXYx2mbFIGVczZi9XVVUBfqyX7Kdi
4mRk5ATyGbFZdzA/neG4yo58dTzWMYI2jO6ufi48D4wmOKTiiDTqWmQfZqUz9tFnhCOQD9mwoKhZ
7N0Hv+XCjOgps15Gd5K7PyEWDymwOL4MTo9GXvBJUYw0+NGLeekUhr7b5/j6Q4VRWW9J6QvgxIPt
T8WfzGs4+5L8abjHIaea6da6XmabB3QzKLdJWG70pwokkGo5X25ZtFeJpEEM5Dwz1oOOJPlmuweL
xosdZ6dqvfzRcBzZSIvfPjuKBV/8I5iPsnTxqAxqJjQpjmT5V/sZ3hQ6tn+cUs8WgUH7CPJQF1ib
F7BeNSHLzMEaHyZNx0vnXwc9wvA3IPqbVdp09g8LOJiU7YR9LUwoL24gD+UpaN5//jB1EnXB4J6f
IVnCmZQgx2fGjFWjgplenIwPbOOmos/oN1ggcMKFqkVo5zkxjTkhPMx5AgT8jEcAHyh+NNWSfIIU
sCye6I3YkaMcB6P+Xnd4UiENo9Or0RlhmhOh97ELaoiy+jQ+BmBosHw3BcI81X7QMqfbE8gqtreh
E9aRg4v6es6H6IXforq8Q+Df4W5SRIZOnBu7jjVpeXFbSM5YX/G0wP1DryNuWrIKGOyEl1KQr2rc
IYKR8OoRpIkboBVPdTwmGmACQnLYnYoV/amMcNZkFlzrr7hdhyf2oqmTm3qxIj/VW6QDfTDPZlH4
njtL0WNk/MXQrHaTvPwB36gqlXqYj4YKTXuBI646Hq1yioWjA5I18hBjaChCm62QOtnR70syZDvV
FfhlkftXNvK9XHk2YmPqII2SQbsQRuDMCE23Y6T0egKHkEl6mVdjC91Ss9heVzIs8o4lyhOY/mTw
vGnLrCYF02eBbtrdybjSwivdAe3EPzv0G35qAYzRkF7ffAyLRX5K+jShk0yeEORl74emQIPKg6be
SVRUEGfUHHHboHXZbzoPBaYVw5W8d6VderPNAonwMWgFasd3Q1ovCJJOyHkn6Yi5yS2BzrXo3bn1
3Z4Kt7zy6EUfMRB4sVn/jQ0oYwas6n3DqL0jWU5d0cRWhSwS5wMrGBrit4b3Vc8NbJQ+FfBC2Vus
/SJBO6XnK6ZVcR8NpS5+XNRLLwyWz7wJV8zuM31YqCjvxfnmzylUnMeqxzqVtsC6+pGWbg6KfFLt
d8YLv1W7m9muHAsTgn220asemndGNWA3P4T8rpXG7tmmyNtfEFkDTLzKeMRkPdRnRfPoyeXzhENb
RB8Tjntk3FkcBmHM4hb5ibCrtmQgjIAlG6fUh00bw2FvtgvnOFpy5kJUweBvJI1AzzcG0IQhoH8P
CI2Hz+mt3w94bzQqxtamsgy6RrRW9wL55D3lRjMoUjRCPRm18zOQiutsL/mJIJHySqoXaSyCfTDU
SIpEQus2Zcoat4WQymQHlwRj0/LFUogq9XapflNDiiXtphOas0Pe0iToOlzpjnPQ6diEaVZfCRiy
501hBygF5InoHIvUFd+0kWfAgfVXqpbL8cMB/VLpVC0oJTmOKUAbQUfRt+xUZ2wHUEuoAoRg9TZv
eETXQrsAFazuX9Tz9XnOv50bD0u3+RkcHcSHSGGU2BfQZK9ytbQjn0HGGrYCkguWxegnI8epu9tr
eMZibzpyQMaeWTyEXFf9YHj1+qY5S5vmo0y9ryasH5JLlB6i1FMlCriPuhacshox4+t8Ziv+xEKy
HTg8SBfdJt+fj3Ud1dHvK3D/sBoz2psZBuyXWqkzZcEoImgs1tpbirQY3wrCZjFEUkmRS4A6g/lr
LhJQsyNDv779ffWOYmeXBRQKL2X5gaz3WU9ANf19A425sB1X8a2z4lahWqsaA6rtqfKlzgn9RPhy
46K1Yj4usLSnfx4X62ob5EwwRk8U6FUM3IAAXkBw+7FnZZGdjQ5htbT0YY5B3wMeTqqXd62Fa5VC
sK8CFeqA2Jti9uI+NJW6nBFQufLCb2GwpKDgsjKM+A54BBhH17uMczwsYj6bKl3R6VWYmJWeoWaX
Gvda6ii9kuEr0UWXQe7xkogLJyAXx/TEkrRhphruQ4M0ZlqX035G0ghnUFKDUmFEhGPkAaWiUC6V
XitjHfFwbNHrHesYL/tRSqpTIoe93lzdtseTGD7VWxVhy9URANDZJKAwuvIjx7j9VOYC0a7cUIXN
s3ExDKxBe3Xz/lvUSa0ECCZj8fm5rWyp0kE2IMVpEcpVYVWdbk3sMLmnLQIXcP5leGnx22AOUgJo
ISm6WTmFg1C0yMUc/mF9tnf6w/1PRRo6zetxv4u8HaOWsb7N2YEdXJlKdTyD8lsoqUPxMJzUjoo2
43+6xzmG0KpsG8zhy1bWr16/rtOxBuF0ca1eDMa09EZVJ36kal202jwhct+ZDKaw8L4hwTjqDFJN
3PBHPjzxR+fwWz0xNR6U9ioT2MwkSNPu4tGrlI4YTyrkwC35gKFTesIdaIvPUa2yDFIQGWEt/bTe
OZ8hwXZHOjCVPamHstnnMYoyIof2uA8t+t1tDB0yih0VPD4lTGaNDPzmmYUCZ1BldhgPb5Gn3FBS
dOzm9/0LaoxkCDr7zZ0bg3A7khGCNN9O3591fHaY3w4VHQG4Fsqe8U/TxncahI5gQIcQ+JmEUqJm
TxP7uCLZqdHpSumQk5KyTeuNPWRGQubRsYlPQZj5l9mnDyWTiZpvluzFLEHh195Yoj7IVmBVbEn8
QmRkrj0Ad1TeZpJKPDGdUOYI6LRy+/l23xVefhHwGUHURP9nSaPE3yIwSSogyqBYtcw1yPCROwVM
8v1mGzPWgG9+kzHhzq1OPmmwOlBPW7tR4pOl54AFJ4iN6eYU/ZKUlqHlTFMbUofAAjjpoJhRVnLJ
5BcfTLqVXMcLKxPTpBDHSoypeMv1ma0aZOju1tmjNHCdVgdq/YXjAru5+Jr7jilogrRLxtNYNaW2
ybDzMa642zDAH5MGK1raA6NfSEcva4RPiKsLHtKQxgwYW+ijnkt6cmasnyk+S6c/YIybsD7Ebsda
GPd+ti0ulXmsUC7bKuP1ejsaj92SJI3pWEhNgpshfy/kcI5TRnlTss8763br2zks6FSbOqc6rR7O
WAX7iSY2sOaPunIzMr9gHxo93ZQkOZX2OX4XnTIxp1Qv+Fv6hJVhUMZ/AGuGV2smvWjH83xjBKPX
zp7jWYxgzKkIi6bbTn6c1gwmCZUtdrUOtzpKaUM3Alo2Z52hQpdCC24YvRmegpbhZwzh1gJvsSGj
ViFk1cdjz5rG7081JAixQgDOIwXBz8SCM5sGP1myalTBsQyhpI6Nvbd16KXgw/L9zH6riO0Y7MY4
HsdKSp+h6Hxbpe8TEK73/wR7xB/olWrr8kjs6CPrW05WqM+o7ESpOLdA3xPmWRsYsuSnK35jSKOa
FkbuWm6C1FJejfJbuirA1gEdH7I178VN+zLQrB36mHyZW6L8+QpWyb7qfSmG7+m8SccTdQKOfLKE
6Nb7e0DU/GD/59ghl4kQ0K/VVIsRLSCpwvheDrEtcWrEq6qOjDbHVZcbfTKLzCrcgHS4znOHbP0t
TW2plpFKshGJnbFKX+j/Qe/uV4YHv/yAMMuSAoUosVCBXNL89bNLSRL3S5pYpsFM3EOyWpGJ6/Q2
ILoeLSK2pxaGtsREHvAU9LSK2fILXxOFAeiTMfEeoU5nuElS1GomLFmjo/3gD+o+FRlenG1l1IPs
/lEl5qL3+WGYiPa3aup1XJ5G13+Nlo9ZMQUxKYa+ijpapLpGe3IMORX6Ut5VXgZW9ajTHpU6+y6B
LD/HFXOjdDlFmq6AO77vz0Jc9J/+15ibnEXWu5oAYiH85uOPe8tiI+8aDJrT0J+Y5aCd/V5HeLY/
oMtvl6KTvZm8AvspJAe42lSoZWzwEpFAS5umgnxEwnuWnzU54DN4X8gV6vTerxMB6aCnZVZ63YnM
XxwPUi7BhVFvCLissaISk/3wbAAxCiFJVI+ks/2FcdaEJ/GL4csRhw5byf1jhm1qF/IL8Oz7ID9q
ydtkkxK09EALTsbPbBiqe9Bg/maKmJRMT4z9pzf0N9wRgyAsA5kZWUSp0fKBeifQPEOviXEiBba7
QbNowYGCI7fSB7MdxYLbNwow5jcGd8nd22XNTPbbrY6IG+agAsuIdM+dF8IdAKNaw8KIFayYq5a9
3HjD1H8gWhEgyiDouA0NfljK2MWuo2EWwjgNZfVk6NIu1zEpak8w3TVS7PyfJoBO5Itgf49IPEIX
lnxokrjCvmyqrw6maWTyDgSvnFzuNNY9WbFpkvNz3fZdqq+f1UckJ1E5Q/9BL0DDjtpBUSCSvuAT
pzp4fAdk9fOW7HK8wn2Dc9Sm9LhLeAp7VOuP/KcbZ1/gP4GvpnyFsccpZzG4zjxwm3+f1ftw0JTf
VeCfO0GskLJcdtytjBF6VWF+RMjm/y/WELTuhiyxkOuobfaYCwCTTJn78JWLvJr4iWRttsy4osXM
WrchxSC+CZ/BbeATAZIDyTdfoyY3jo7fB4rmKkofk8Z9mogXDNJJLkEhSBVSitMSedo59DMmNJQ0
xKC45dch1DjgPuV70PZEIeoDsMDZXA+wgJFgjh/OCA74piYJSw+j+YoLEqGYiLsCS+3JGu8zMRvq
sUvwVu9VSg3NCFjPVDPPGJqGo8K2q5LX95kNbCgKVlOOl9bhi5hef2dUKKZDKR8dgBaBOiYjwXSp
cVG6iQWgOPHRdp3QtjhOpELgvI1BOAwkzyu79RNPLLOMQZNru49b6kDAKiwVMmYHebYBw9V4wdAe
eO30eKVMLlzcfm75xMqeb4n8V0n+O2Nwp3OHlMUnfATixjpxU+O0xyH4ZJkVMYR48qf4+rGkIXIT
QGbpivC+lZxuyoP/Dk7i3v29tOG2OEHiczEtcR/hTNcXSXkLMNJzRNkCHA3Ds/yM23EW7vb9rJFH
wbQs6QeussPZpq45QMkeFywW3aTD8bAkhMOhXhYDgu9GXUliYoAUX6NmAyyuYtKdc3WqqZrBwtMU
Byy1/zZfFhhHP4Lc/wc77aerJtHS+uKFyqXK7vtbJ5cWuMlzuVmr6ywD+c5bFTaIRqZOMCagPrAY
p28Eo4PENCXFPxZsy0WR12dKMs5Eoyi1AsK5cJeT4Jc6+wjAjPloxMe99JWW9r1czOIwollnW0mO
IYuBFQ+wVCcVRduDhXACAHDLQXtI6EGpyqVCgqKoWJCfCneMadn83gOU7SOcDn7X43HgDjRbqw1y
fsDjCYb2phptM83KmUMEd6PTcb2S/2tm4OX5sFFCcgLu0RXUMhR5ftjk9i5Yp0+TH4UGkE9dDFBW
CeWGMVJxq+JWn7osUwu8Q9aIcPbnt0EPrJU4VtopDd77HtjBvOPcBVsWtL3b+3ftBUkc+HeDBi68
vL+2bIAktl5kEtvhK0/t4xoQt7a+VATvPxPSojgWgRtGQgjr7pZO7FHyXIo8M0kw62OFljvquobR
UZosmqe/k1a/vVJAdLm5V852dH1xVh/AdJSsbPc9pcnMUkEffhY9oB1PHMcA38jXuvp3I4QfFJXf
GXYqvUCT3erZA6FeKX/Ut+p/vecqLwiPyomqlE+qJMWTygpomDV0xHyTxacadSFrHc5HY5Rdr/kr
bBUcOIF9X3A9e1ekoZPCUPTS5GQsRe+1FtxD3JRvtWL1+wEUqOA3pUPrz8FpmXX06Za2TD7GYPpE
D9K8bMab+yw=
`protect end_protected
