`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mwx3IpM1x16Zh3FgAFy3z2M1q1tVZ3so6sjtCnsRLT2fff1a4xrEcVpLcHMSHpoI6ADEAiND5Yf8
4kgJhjNn/A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RdyiBlt/gW78SKhT5Ql+H9N120mRUB1Du9vnV2jPooDfjURpEaAkvmmveTupr7MxRsTlt9PEiHV8
z8So5YpPEDXeY0InsBN66qwHhwakqOHRyjkaaS6CC/PTjZzqSXCR0VRIxQz4sg8d7bZkiVTFt1hv
eKpvPSB5SxYWv8bO5DA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EJFRV4g9f6//tDpjq2n65PW8hOgUSQU+hvqF2ynXCeZr0S/4ll29AQjx3iMjDA6HYWGosdxxm5Xf
i4mBcwx9MFbN8vdeTWHbGUwzaxcl1pt2E6eDNYRfPwJzgE/2A/IGEkoJkbOH1baaBAddFwgiF+AB
o5Uuur82/m9DiCuS7ZWAv2/80emrDW2btc8YTmdr6N+jFoIspt3F+gaveqwNEsplz13I7db4E3kL
sWMhUqAySmZaTotqb6YzzbaJZzVR0CMKBVLGZCiokKOauETsA3lQN/b5SreP9htH0gudEJ3odSM1
RBtF6+F6EgSQQQMdqdBbZBnMACwDhz6jLIrblw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fx2Basn20pIn3VxNdaGyCB+CK2SsSkhtD8j25zi2U++Y+zTQSmQpJ01W8Nho6nM0VQT18zpHD31H
Bh63oassvMaMBH2KLVGpFCqtd0FKbPRkZXbvhmdyut/lCCUZUHz4pet+Ck0d4JvjPE2Ov2mJvolc
L9MtMWr3SQJKmSTMuiU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ncMXD4xXCtaU0Syz/N7ujJqMVNKqelhT1imBwP2YkX/2RKlNfvF/5V8TiMRD2a5RaRYaviRnVVEv
Xv0U5eJd0Ubj6PVys91K9RF4yx5ITJq/gnRywYodZbONBbAxTHVymNL+4h3VSpMUHGr33b1pO1cU
twjB4s87MHlaaF/2dfLjiwODcnjwgLru/uGpDQwJqCQP74MfrKy2FGmYYfcrPC1s0aztexxzNhPM
LxXjerWALJTeGHOW1yq9ezsfFHF5jXEsMZZvVBlNPfy5ofeYGkK4ygKemwf+pvAt17H54GS83jBr
xZ0r9+kKB7Rk5IBTt3e9LNJrxquE7pKJSSlVpQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74544)
`protect data_block
Nx7UIW0U2a2YSX34fR+bX0HY+ex6yYbBSrcVoCEPKtpRstn0ZJf9MELtRj0myPPQLJ1a5OZw4i1F
k0zsqsFur6l5Y5Z7pFyW+WaW/1xy5C6IozAB45yzy9G8HMCnRefByIe4T1Fl3Ymh9YXfUh776nyJ
OUH9Eo/Fi56Y0FmGrRX42PIwMfbWNXMJ6v0Gw8l8ohf3jlWhFS7u+eXNjVfiwRLOtjgpZ5wMJTHZ
mRh90FM45WlqVRiDIVAnxqZsBpdK3TT9IDmIHuP9kWYJZvgzfu5rNwx7fEfKIkmV4ucczyxetS+n
Mtx3SJvIbCQtRdZwnJR63uvGYKnW4PRrHaFutB2OnAqJlGuiTD51hQ1JaV7QAvRNPfaMYgtcBQyY
KlvY3VU4hI0syaKIvkWuk2gEyS8wneX7/4LmLTIIwo7WMWzcRHWzhmSZ6jOb5nWUp4ZpG+HIkVUa
GQ9tjVhlCdH7xeno8UHHoNq9zOB1yISyI+YysmVoZo0+qPmVM5cR2E4wOke/+k+7mf16toTKPifb
BEV26Mt4zOA520BnDYAHC9mp9yBwCIdmly7aPZZLWTaoPND1/4nkFIcP9LpqUVUI24IWqSSRA1pX
WyDX15KXbIYcb1XaZ+IeCBg5OfcJYuoRbDwjtxEGdUTcVYIdVTzoVPKxYbCdpB58BX2UwzTWoR2y
yBztDZDx3/HpNyqm4i89X0G4yj/PHy4/juP1Oj2NT+mwqZfFRzNN6X1pAkreq++WFKdlpEU4Qqoo
MuThRLiZPOkHm5E4t2JY36GN+FiKXWdvtM0dpF2bucg6jbN9Tbb/IL029OzTwWwNnFtRcORxRGIx
jmEikEK/22dGnzqqlcnIz69jos9/Zp5V5apTsaBmsS8dqZePL1yAJ2uyxw/tMWERFrtQWRcp4h7F
LjjNBzGWX15L996kpn4hVqGP3UU0yfSqYB1V4AIhGmCgSdfYJ1tCPFS7o8O+OQPk/oMdIqfqKIV6
nNE33s7D9GjqehCcAUQLH0PJLgfPw1G4xWckjheYjkCDMAkm546rs2e2z2mT0oRdytQJpl00755A
peZW15Ck2D3KgH8j640GVQLtx82XtHcdP+0aECG0riI4eroVTxf5i5i7fBmYnhyGaz8VuPGPMvkw
XdjJoncbRvem4lB6QetSJ29T7d1NY+xpVUx749X+hprmPzQnAlSKB6mEi5y+55et3XeJGY/s1Ov/
ss2S/uZhWInCSpeaUErw4gpJGZKC5NCZTYbAOGTMh/EYF/tHPJzJiO4yX3AZEZKdonZw5n0VxzzM
rBJBoy+eJCDbUBqacxYDzEutAXz+fIElYh7EVuZUl79ppxLrHofHWk/XC/PMtrLvbSF1cc2J2sAB
A89O13KgJYW6xXvla7lJ4l7ab1FAy7pVYUSIql/veCPfVkF6y5s180SiQqG0gNEUixOKTp1zwcB+
/xLZY2+bLRiJt7SsGjwjj8SlYHVQ4fIp5GjgDqWno8goAGrGa76CTr9z194HkEs1caj9meNDDb4R
Hp0jIHBW5gSYoKRLGgeywK6fJ0ZWODi/AhbeCFhVJlpA4dYtt6yHta45My1V9+MVxhNFGrr7eqb4
64YiuzD9TB3gpjYMmr7oHKqKMB4GqrYwXCmrvlEzLzA1SZrp2IKfqKI54K7x2PYtx6ha6KNqNPjF
l5IURbz7zz0CgsZQ/3F1crunZI4nh9CorC1rLxjPBDORTb7/qJTVUCiVUwAxdikXsJGwgbLtuVqz
OCmSJDdxfg8eMhOIV61twI9xLqvBCK1fmJNbipO+In1GdkM6D9k0/u44IaHGxro0khKNwZ7Qxrtz
PMRHZXN4oee09JCTMWuqqkaOks1RUXLTJSle4m1iHPQMSWI1rKxCxzSMHBuAfZFukLP/zesVOpMn
9S8+Oztdh9CJ7NNPPb2tHYG2YbP/dP8Xr2MvVaeqIeYXYC0IQCGg3Jn13cNiy+SGSlVa+kggFHbv
enYKvyh2jKqslii7o0b6EEl8sT0a4fFZlsHJ56XRfd/Z+wGZe+3GHS1b7MS6mPFm2xR0wC67fBd5
phWEU/YyqpsIxp1UY/wHb8pCA7xm4jeLfryJn2s2C4Q8CaRzcDhSAu3qM68Io0FCBmArj4oINV6e
OM13FLf/VRU09Ce5I3tZXGpvk4Wr0sidkhi8kYrVTMdXmi/qKWw9YohWukLUpg6SB8ALmUjliEXh
738UDBQHNKS313GIvgRRlGvb1DAfZGOhq3m/yEDDqCCo9TsrxZ2OXhkry8gplEF4icVg4hUkOmIZ
bHN4DGP7gsHCRI4u4XsFY+2khmrQmTxJa7amDA2sOQ+HnPxZoy1g+QY5TqvXiRMjQmNtfyoZP31H
h1WKlnPuYvM4NyjpPi0n4S4PXLHI/GWrnrwxDhdVBr2NRdSEBvzslG4JvioFOdyjSb+bhBgV2a9C
gObIUoYdl3XkkimKD2OieACZtWqufCCGRklA3WFnpRaxlGFB+UlmkrB926/YTDhqGArjxbhg6NZ3
+e7iXLcy1lCdyUoF8G7GkGTewIiO1IFlRuf7qRiTJBntdsZLQTI6xYKM4Q20a989M2uZASAARIUc
b17+YWMNbu6MAuYXG8x/RiMDWdqddwiuHlZYUMArBBNDSn7CbvLoBlJKx60oCdsYM0FBPZB+HinH
f9DgQrsIC9xr2uM8gCzOGV+rFcuLJ42hWjPFncTEt0+4CfT8pgC68sSa6xbW0tLD+hY/2IwmOgOU
C/RQNab4i3M12ho5Cs4X1ifYid5mYS4RoQInQsAxf7Yf02P2MMljgx2Ov9C9y0LK5oThVo3Pd7s+
lG+5K+jJzsDLw689f8rpQcCkFrJpmr3vtRwJADgXK8dJl/uLr9rYEbhr5HBuBvN8kqO/zTkAuMUH
ZA3Am1dVobt0G2dV/ASb63IsVu+prol0XLkjdFtB4cYfIh235n+Y5x2jBARqJEu+F07DccY2dXiN
4v7RwvXm9pfEgY/AzNUTa7UZdxZETWs2UogJec4vhcPnLjiBLz8lEzVXjzEI+EysXIfIxPYL0Jcc
K8L2LR2o67MaVLd7YkzMszxmJFcLO7hACdpwGpn/NwDo3eVVnZXTyhjkNtKvUEJRb0KFUKQOW8aE
1s1vw1LNLHPLWGv22UoP7OD/UuKE3e/GJyicL1+mlyKw+7fHyHQR7zDiQRKHRtYoZQ+gM9vykDpO
SY8FRygSRmo0j1EZGz5idierYamGvs4q5zyaax0eJrSMW/SWhnasMDQufnfNdRPGewsdGti1wMfg
OLmi7ArUDZPH+rYmfbDqEz1+v6I4cm5KFTQ0kwgcUQYX2R/JRDI47MCv2bqLfpPbM9O4hhinteWS
sw83HEtnNNUni/yzKubvoBIcDfH5xkyJ8xwlv6DBa8TrxCduceKrPyAJ6V05ITEfVq6AnUt8OgLS
sBylpRz7IRPbMPck5gbITRSyTp52+E4Di8/VZg/VqTNbCma6rQqbsmA6Fz+LmJ1PeIEkKukhX0O0
c1OFbD19oNz4PNdSYTJ7UNEsyK63Kur2fLawQcNnOcY5nB6094i2SzqF9x+r6SPyvo2ayYLBnTjp
dRnYvyFFVeo0s2Wi+PHsJapQqC1BW+yL2Jh7R9MrHvj3P3FN70lwa3oE0vJg7vjc+Vib1FJ4iq60
b9xuYiXZvOxRB+GQrMkjhWYbE4zTuYaRANNZi1TT+z30bRX7cxQckyr7dFpDaadLFVadWLFsUMcO
mBZA1JaqJWFaJzyq91RaMYtLyEiNDFsgIu6wG7t2kbfpgzasMZU/uwGgMaE2I29aMwutK1SSkM/T
iVnaiUVBGNF3IoqdMI/cXEWXxx/JKcOBDId6M4XNf8oA4/k/b8NQ1lHX8elAuTP+SSGURDHkDRo0
ZooUQmEYF8EKD8ujiB2gv3zO2cSyVkj9umSAHirxyl+FncHoOyubHgfC4OT49Ixs4gffg1JTRjKK
kfIgVD+GlPob9XRs8Ql/B9pcYAtmh78zVdF4hjwXeY1OV9F/s6EeMaK6yJdlkygQ25OrmGbuILK0
3wr/m5DRkMzbTHKw4lasT3+J4s63he2R5rXlTKmypQ6JzhONaSxXw0GJZuQpQE9Y2BetZ8sYu8+0
/dUow1YTycqAQ9SqgSaBNI6mtyaX4A9Uz7uvoEm41+sAWIhf933JdPvR7G3WOnnP8gKoqT3sdaTm
X/v6BDRTMzbPEJfjoUHkd7T1UgmUX4NLaxIcYWRdb4iQ/qlt2EDuXCC9DoS9cYUwAEitli/Eh0ZV
h9mL/O55GeX32sM2IlkdfM/6WJKE6kOePwBi17XPI6iKH2t+qgsxw48iNRTZpW4Jm6PyQBvcRpvb
Qek4QMEGQKuagfFXDHAnDn+4KSDGHavQYB/dHHd00wz9CUm3VYq1n0hEsLG57SKROulxXpsRUoE0
fft+RI2l5dvH63MVCw3KKr5mPYQwygDpu+eMSffYfbcG0d766KI9mPwnht/viKzMmeFhkJeaxNRN
rsn5PC0Mi6ROx++rmNSFkmZkjUkubORD6tJjhqEcp5f17XiqwsY2WbdtnlaOdkTx8lSqgOkeH+t9
h1JZIcXcaPP70DkD/PHQ8LUSDNf2hYCDnYJXuiIgbwJN/n3CVjdjzCWE8FvHQnNeB+CWkcySkiFb
Flu2ZSupbfqBhzmD/9tXzI41ecdkcA0TYUzRBFuzB3NAZNKqj00TeEk+ImUPOLqStu3FFBg24wZR
UicOfJ1jtOtyTfZy7uGD8IjIsAlVvQvM83THBGxQw8NsLPq0zcMcDruYb2bY5QSMkMAiCPOkLRpX
7zc5wGIoGOcfty2woZje9iVCVTcwYdQXPb70io8RinHaoMepN613aXtciM5+eZ112jIirWUFIh4E
FabzNRl/UqSyWiQr5R+gfAgZFW78Q/ZCtG1IZOCTFR82DkPt8qcRmGVqMrrIaOz12RyM3QWU7sRR
XAP/590lMvTDpLXpUPesbfSJLos7PaGMONs1YBY0Wn7Vz+2XC1AWot5NIsjXZeHPadxa9OqJU72u
jATMXDY2oHLIdKS0Bqd4TrT6gzzYSxUROkzgCVeke/XZ9IpvQtMOkIW3xqciE2gL7Gyw3f4gTimK
+7hiSGriV38d6GAd8xvUbX3bLGkMxMQK80GBZ1pdFu+zvKwyvc7h5xnsQaN9/q3UXgh4AK2A4u4j
RQZcvOg2Kp5HGwXjsy1Eu0EIatJBFQ4+BoI3DdWSSFlkkhZNIvq9tvRgRTyVZxG4YZ8yNWveeeoL
Cxpz9luEfiFPXqjVL2M6nGHVI+508LuB8shd0/v7dZSS+MXTgZHcxcw9e7fvWH7qXjuZ4C/mqNKR
ckqDHKgNfBquTmTDo2UlaErGrex/rzmCIExkzvkqWRZKjnp5/GUkFPXq5EXyq77kDDciae2Ce8JX
2ypTldqeJ5VA9r0qDxJ7GKhBbJDEyuJ2wY0zqhrhcDTA5TWGHt50mqqHa07PtCoP88GkvZSbsf25
yyY38CnuUgBg2ZiM/z8dGAz6sn8pEje/JXarg5U3rLJyGqowBD6zUMIoOL83nNLnGGKDESZUqcle
d7Dr16/p6XhSTUKFxwO7ZE4/dVFxPR3uyY7wf2v7lLdpzGx1ILpLjgifVPxTUNRw3yRBelCUs3sk
iH/xuHDGUySsmOJL5hCX4kXCpfZTTSsQydF8VwJPsC6r3Vo6Wuw1SqTV6aSmXJEFzVD+qYnC1EBg
U0N4CcQhsWsNv6G2pyZzF1oX5RYAcN4dj4S8lHqA/2nOgz413/21TPwHWHFIV6PwLuCYuPtDO60S
xv3r0Xw5gPmfmyFQ8o3y/pcSXbxu8cWns5nD8A8l+yWmQ3H3ZodxdAQ7DfSuSCthl6RQ0jJMdT+l
pLTutYnF1T20s0j5eT767AplACqQO0tbBuryv5raCxtTAEH6bXgSoSGZUwrKWf2FwU7aHHFbQGne
70D1j6sNI6OOwCJ1N26RsDk6T5J5ptjlTHDYKA7KoBcVst6kyo8MtuyICohCp37gbzhnnOpApJhn
cLo1AxK9dYzdqx+jOhcC73gp9P4mM5VQ/6cC5rX0Wr0IFGEYYVptPRzX7Y7+P3lddhIyZbtr055X
rdHKpaPYg16gyZY0I0h3Dcw1hrE6bZICmR63g65InQfB1Ed4BpB85tSXKT+RPVbm82i5v8Xjj8Jw
0Txe/aiuQrmVfS5FFe7eDVzyV4Mr6io1wTJ6ThmLghMNgQ55x2DjjcFRn0rWxkWJ/4PJPb0e54w5
8gDtRFpaE93PA6vGRhzZbBe8ValyifbFeq5MQg7+oSu0Qkw/GESoNQU0hyGebPQyb5Sm0FgB5MjY
l64sl4VhgtAQ7Vj4BulNQYvLkJM/gkT2GthN5zWh8wZP/MERVDr90FvINoW11MmEjvBGRakLpizl
qcRovtXuii9jrEGNvmvKYIHfiERB0PwBS+L+IfvD8AUkhUFILuCquZm6fc9+ckwswCqkPCwDshZU
u/ofd96eTv6xi4q3T9L6FIvKwwfS1ET962yLqcPhBeTyvL0JQwqSWPAKqISTN/4s/JxzndBNMwlE
A+OVhUt3b8Dg7iGbPkgBBlkrZ++l2dX9qcy9b2V+9Pp7t4bhZ15SRNLYPviDz6ty+75h/vEzKk4C
q1TQUNCWCR8Y5cXxCtSUcBvdI0qV+sCMhTp/n/ljarL1nrKv1cYNGUpXKTvfOrxWuwB2Xs/4YVZa
hn6sncmHGLLxxgCavwDQG6vYI/vhZIOPugia7U9dpP6c39oeUepnKArhb5Y+DY6waOp87irEWojc
1ytMLnRjifXTiO+kGnAYZFlrIsWCFdr7Uy6ZgUBCj4ZEDKQESeSPCyqRjECXagV7TCOLrtLf6mn0
TxCcuXnkwxXHIIxzI6cLVWD2ycwaOXeE2cg7o3xVSRISIGAb0Q9K8HNFBIm96WnQlIpWjC3uSdt7
7i5ixe6DqkFinh3lSIf+VT5qm5enE4IJ99xEw/OwYJda00ggLUPMfoaAyD8+iAlhVWlaXS4TNXpj
ONPWMt3FLgrvOtmWAW0Y4tglyxITMACliRTF9kRt3IVfVW2wGjVbYyXMsecRmYKXqzOT+W4+tvQ1
nEER4DG3FHNmzkKSsdW2G4ecrZ1GW/pmUJf16rsSeI/g5iTtJvD7Zg7qTp3QvlwuUaVG+YM7DV1f
nNwXxkvjhRYAVTUSsqsuQ3KW70VaY6SZQMFilGYUwKhD8zkbHEkzO0aV/NlX9fM4XBHqVj/O/96j
KGsTW/qE8EW6U7qdFWykNePnbRwh86Y1sxrBpTkGqb21nFvmEjTHZbNhiETXaH8gJgrPa/buDI5I
Nfmifh37OteIQE6Fl8Ski8KPhiLF+y74v2Sx+qNnWZSVHLZi+zy0oQHGDr+S/AlDWiyR8lIU3W++
wM2FDtLYzE3rz9/peXwVp/Z1xA6OD39H++Ys8LKczx21SB59Z7jQv3RlcU84VrJbtG12+FvmOK5O
VPqnfgueOmhtLLwITlACpNh5l4SrH1rEQebDyZezT52wvWv9qpkID1gYoXkrGqKd0gkseFDPYLf6
OUCbfwMrZEVJ2ryPVp1FbjUwLnqqubCoPz9kHioeCz0qPMflynNA8Rgdg86K4yfNQ6AsZ7AXoqSd
MVHITR9dxp6Z16xhUGTdk79JG1lkFp0JXWegypLUHJMHbBsfc9R1d+ORmgap5ta5TjgyTbKd5YxB
fYtSeUr0sh0FwasnhswXGCrfmqz/NnWIJkwvEiHH5xAXUNWxab/XraeKBFZvDXOEzMHcw/unR6YM
+ZWeQmm4kNa1wP4Ju+M56kCjIzPxfBfbobQs7SruEuHhLnnpWQB9JqopfFEILR7zNbvMFH9/+bbV
WGMyBP3XfGYtpWHBQ/Gvwm8uvsNtJTHs3pYuEMtI011k8e1r93HdoEObhvYrEhgFk2T+504bNQKO
51bvMzkQduttyeYGVLRVzIhUMrFzu5372hudKjjOujpoF90JVU8aivyEqQRtcnIX9ga9Uzbl4+uZ
mu4xuRU9EJ9pmhchbQDHBK3uNg23nlMpy8JwIE0f16DR8XN8rTtrszTTfHi313Lq6ii+2O3hQ6EG
khAndJC7PhfpB/EpnSjvOJEClRBQYWGvpInMpWs7IElUzcmSoqCg18iz+3WX2NsKYQCe03hM/BZv
sP7hubQhaeYizwmb1juSmSwdsXeklGA/Kx3BdKLoMi+ckoC0RKwrDvq1DUOCyTawh+HOlv5ROyTf
DZf+fYum8g06jbpbE9idEWkpmqeNBElFG1XUyoP/UJzAjYALDBML4aOMUlRnZGWaCQdtrLbHNtNT
juaoFfj+fWe0VrhyigHVVE7QZGf8kj1MIayEQBbwgOjr5Zb7apnb1V4dEN5eb8php7k5DuUI5sKy
LIfGeDxviPoWP+gjc3Gr64EnAux/Rwie4Uy9uyUqG5cVznapKEz2Zd8w41QSOo9be7t1UEXimj1b
Ymg1Ei87NsOfb09ej1JVugSaVbhxqEE/tAPEr6C8a9/PEDFY9YZZEdM7ygOoue3OV4dn8Q7KwFJu
1iYLNsDjpNYFqoHCLfXW0oPZcqK8ev+r/1/pulIZFCSkaAt1iQd/qLQJHSmJ96F9TKm/3qby4FRW
aWZBg4/2m0OwF5SWNtEaXjwULPefuGZOv7vbUzWZabatWmVjeGHt1gxuHNuwmDikLTVgHmStTmsx
3OSrV52PFqEdH9ONv3TG/7jmCNgMw9/jekdLYKmb7uW7jcpyTVUVFCpHWDjiwwP44UoUYMwQxky8
f/D9eagDK091KchxyObu3G/Fq7F7xcjXEMxjBkvKgmeEMW0a2Cu0L7NYzD7G1c9v0m6AD+BhYxcd
5rMxMxL8UuBg0ilHrDlYju73AMA1hHAHN8M++VGyXntqEKiTZVSNAmJT8Zge24GdkDNoHprS9q/G
UsHfJBm6QR9u49vTf/y5akl36Mh4aea33mMQFG+Ed8iAjtp2rJ+/8qNov/V+enBj8kZiccXhq7ng
h1nL5U8dEIwfuNXBxWVi3kbb+RM2d5GVx5c1Np80fxllwZ2suZU5jGO4olcoFlEKia6lkDZOE2Ny
C8kjr0htKp/WXK563KywbWenDWpsSVUknwBP11oB8KlxtKvhHaeADt/0wydclwJam3e5++e5KodK
uGigwLuFI0NVxe0Gb8nH9N60Y0ob9O/5NF3W6tzMlL7eBlHYj715MQFGS/s2wTOQ+f7Uy9C1sU9G
ekUQu4v77IHDL8S2QiUUGE7uuzCEHDWT9FOmx9LgHkEDuvSuaVpLEWcNdzi9WFlH7BYmzWev5xqI
EnpIZo92M5QIxCw0i3ocPcSx4hmCITJTyyWMe5Jo7tYDugJLNaRK70uCZbAz4L33qVO/rhH3wQng
D3iYkmUT9PnySZk7Z9AgiSk1+UEcx0skPhHh/hVPSMO7DAL/Pl0BnikVc+kAZlAZrBJC814b54y0
na9Y3oMTxvZTezyuMQaO/ZNmnYBxYJkOFtkHLCPQQTVYH2zT2n5HmYm3UqGdof1NuHgJHN3sgYfp
tHrl/DjHd4bhDY1mUagvWU9LrcFVR4IUGbqFWBXYoSiWz48nITw5zEdKhCSLEHkZj+VxL2P8X47x
vSTwn/ZBqKrll/SDEXcmt+QbnOUGllLxVTa0XIv6orIZz4W0K6ZGsoOhPYTIAanbCG3bfKxvgbU2
OJ1z2+LO9F6nY9w11GTH+OiXBw0CzYHEelsz/AhwqyuQlQs8v/JSsudz5wou5yRGIC+iZZgxgsQa
XJKf707VKFxQ6IpZ/IyBcsYt3XGKT2qLB8vlhNksJWE7yJTkf9hlpH5YD4UHkiVQmKFUkcC9Ekfl
fc2y34c42BnrF8tpIOmEz0O+05sUhkxdot119SoUmlCz9YkMeoYyT+40NncuCWB9legiXpkdHjwI
Vg61cngyDeOFwtGsZnW7DSreAHrn21ISelrQsrqE+ShptnKW1ejOjha6eXeMaUdMA+uOCFohxCmB
G9GKiWr7hnf+6H0955XnEA7ME6D1Uxsz9OF0iVJQ5wfIWAAZMKqqwvP6PCvcYBBygI4SGGuU5yVQ
t2ZANxJsnuy49R6rb9WJpOfnR9AXBi6zTWR2heNg9ZwzxacCUprIlk4hUcUq2NY0op2/YPIm/7yE
sYssDhCQVKygCQa7D2dfN4kJAMR5mth0tgptu/orSyLa/NFkAeOCKeDol6fSnufK8gh6UCE8eHR2
3Yqpfav2SGXSf/+pjocHZ16iMsy7m79RPDGUPp6AkZo8vGG4nVzgwaW6F7GzRMi2a50RFOXC6bPb
Ddd5P7uIxKqJ5rO4sgkCaBs4pJd0N9UXtJ/RsDKsL6LlK3ZykvB/YKePGlgsJgVvhx4h4O+++V1c
VatqMm0QZxwlfTevrJtheW+qmIFLiUwxs8V+NFa5xjdHQxN+fZJOUkEWLNubgrhRUUzIAanwq5b8
6zvse++p7aAS0wjJACsSsylhU+Xt4KDbxjFU7a5nY3zFaGejZMQepLy72qajm/UoiI5ZXRao82Zm
zQnIYH6yTugjJeujiMHEVcsf5K6sYGo+RNYjZCPm+TRMnUCH2ZTtY/tTiVhjaBbdOSaIjOkd6kkS
/MUFYxeVn+E7zwtttlQJBlw/Lg8Rv7h2mp9UinuwWdJ6555DSdJk71WV/RrkBTj4LUA/YlxM9MJe
HpQjVyXOQOpUeTrQRe5bYNd8ABJee98GIwST2HU4nbEYvSWrw5AufSOgDl1bu3tkznMQjcmzO1F7
RtvNpUK1EGYJTgppS2bAcS6qX1iN2dm00p5XAqZPcWebXRbmNsVsMIOtdUsdIFnNJ0OE1GwE9fE4
+pc6YArCJL+Li6CueqTfA2xnZphsCV/ghxO+Iql/xoTN+DubaSO+WO2Ra4lw0oWaKtogC/sPrO8n
ZWhoDRBGkHzyEosbi57TnVLtW0UBIjArbUygcg7FU21L4mdMnHy3DXmsFOJTR9b3CkvAatnPvVOX
nuYKlC0fmM7BHsJr+qDBxwj2x0tlzIJQI3W0W8vyhIK5xX/d8H7QASFStJkH2pOZD8KZqXKhq9/6
rSG/iWo/bemsUB89rlWJjY1tt5/fQrWYCHpylg3Gfyrv7j8HENvRCdYqhhC4MuAUZKreOHTVJO2x
Z6kjQXGAznr4ClZsFq6jlJmE88FZ9s8pyisYgMf3FLeEVpGppmARqmCxqEdMSRRARsAm4/iAXoUf
RG5rBXHd3B3zP83cMskgEREpi5e0uFORYS+CSNncVaZhhdnnwVojtqnOefx2+ubuuIzMPVnbHi1a
kxEbzV+ztmOt1IwHyNxOrctOMeVlSWChxPBlvnyvqTKdZku6BLeFBU5568lrr1i6s9/zOo009TMu
OM9Yz42kaM+i2s3j+JUOjtjY+eNv5EuSPt9Os4bhwF2ons36XlpzXjup1+GY4RivSdPhU1mlXnSh
PSYZHVbZq/XAIrJzU/TfHN4ygKREsdooEYwvNQpVlJyuMUYwPJemCvyuXiJV1aBqzK2xBZEsCj86
BiCtoBtTgXSLaRHX7jh80/b2yebfcVOvaaJ1dXEmvH9IXzPUFXNjyCcBO2d9OVpTCU2VXe51Nl8e
uw5AVN5MFybVcxHtAg6iXl2jhyD7pAcRHdvkX4PvWbxyQBH0fZUFwWMPsdAvLQy1slfQjSXfu10o
OhH2ivd27Bhjlxwcrx2FXCAVSKnUtkbx/DFzHbIq+tALROMICzU2dNTGfoi1epJGRyymUnW0NXfu
qgNmS8+Tu5nnHTLpK9bFqo8fF4DGaIrRseOC8QF5XH5jpjBvO6HF7Wh3rZlImUZ3GW34QUW8PaD9
6WDQu/t06fNvjP18/KZ5ed32dSna/PCtVw4K4UopLpRqjWR8+Cmr6mnfMuCli2XsDtfD5+hEoxYq
jXegOKhKqUZ9r5xRtAOEj/DNOSpl7SHZBm67OAiRZ7jRJ/vKszOSI3g0CqKCgNE0il0JTUBesSSo
1gIdsTF57ez65w/9m2Mjg9FgZkdbmPffxkjc5uCk7iAEY2K28Uk+5/XBZcSgVLiaESCtwLr32kgH
JsGqt6dcOXf9DIkPZP9OGbLM60QCHME2BD9mTQXpa9DsBAq+lNU7+Z6ZON9M29WjKB8AzLy47Tj2
hfjfGE8I0g/D89ygLQU4x3siSy0HC9PsRK5TGwfSynv5Fn5w7jjVzf7SfP79u9KsRD3Q7qGW54Tb
fPyaR0sBcdFfQFUrJPZkC2/UNUsuw9wUHeWkMILmpiXOXgOmVq0FUYpYadFZ9jwtWhSP2nWdAbCW
FGZap8sgGCUa8AwVQzjXpeAUro8A/SPCt9wS/bm8O2QrruncKZ0DHHw60JKav2aDeqqsRSZMaCUf
ak97nG0K6wfeKiXJY40Q0oXXh/zXbuoTy1zJ8c5V3SWzJLYL5l1kad6vC5lUZfeUep+xHfy3NaRY
k12zNpzzbco37o1Q6gkfhQ/2Jv687UYt+Abbw2wqEV6tp0qQEci2ztlC8pEQyQHEjNgLdvj5m3PV
eiThLQOa4AS6wmTWS1fM2JjuBkawygXtBcUCH++7w5oe+uTW2fcu0hpyonQtt7eM5Jfzx0+HsrpM
p7wNMytj4Ch8JhtCOItijAx8Y/0+7zfLIqFMCu9ASfynS9xONclvsitGeab/Kyby5rXZoGkI8C5t
uEUO6Zad9V3/hmOOP9pRpD1wO3LrzeugF0PzATndPnA3yS5r+tGsU9wJtbgOTKNWE2aMNP/pxukk
WQ3JzJPeK8UbH1MJ2sJB+OysIFPOq3sgwja4VSwBxMEVgMIK9+fVNxUMWshiZazbpcJW3qeiqsBc
kEvjDvlHg6/jbEa//mekKYKqxgzi2mcPChR/BlHde4DRsNR0c0q7yL0PoceTv7QHNvgBcyfzA2gP
q8RBWQKu4Txfxn/8IGOaf7ABf0f3ZDUIvu1dBLqeaNpfdhlmmF0/EfQW2cJ7aktxdPlBdS1K3Yt5
rJYay/NQYuJ0m3WdluTmXpdF0jSv+Xk6BvtqD6npSjhuPlbqNfATwstTV2EKfBm/2WangQVhXwzo
ASimVaWEUocq8L/UjOyyfbA9uqZJxQPegRb9gHaDTwCRMsK0bx7U9k9uLxXF5r5hx5dcQEQujXCe
Tnhb6oCbUE5aXLvIEUZi++xqAM7+tcjxalFUKoLJGf5xmHOnY64+qjp4pjS0gjuvQBuKhCkk53II
eoiAl30Uc52fT7GeJBUSJG9i2/LqHBrmd9sPkjz5QmDHHwB5LsnisAqN65/U9RnH5C0OtZu+ECrC
BeLmoQ5cqGh6/FZYmutCZHzgKr5t3MPzr6+ych87rm6zfiM0mQ9yEgxHHEduW1WeEmagQ6Fvu/aa
YdioS1OAnL+OhfSG8+EwrlUsFKrHDG97qaLZJ+HUXlHfzVXtLQR4g2U2Ix0SCdiv1DGgApxEABUf
DZNEc8NTLUTRs8reiQAYh7MpIJs7aqO50Mz3SkR9qet887s1nLq5U1UqOuwxXp2zJ6KGZqv7x4kS
9oaBlYIBRJRX4kIO1VRT4o/ZWsWNr60ZsNTp39LVTefLbbB6gOJBWpHTbQo36564A84P9fsbQitO
c09EuVEX2lmffJsc1oRVEcY/PNtAUuKe61FMunljqEq4psaSvY5SRg6/L44CcFL+ogWH64kg0N/L
8Ya/G1/+msfa/dZwqCs9AM7PmRuy+YsdgSuAKhVU4wjHa5exoXuue0KHkt4gfDeyMkIFVRbBAAVj
Yjy4iqOcodCXpFv3rxxyu+QzUnEfEAEvdddSNxf3hDaTPpIuZLdBsJ02LsOS6mrDYHKm38l7LY35
T5W/MdYaQET4FUYwSevwh0XI5chfaQvQPPwiVfg9iruWLtGbu7fjX5r56w/Ua74xuFQPbl4ZHdt6
3vxALSmdyZvSklbBGyPjv/shida9rHbfVnwNY5/99glxPjLzdVBPtzS64H6wMT/jV0xkHteE2A51
8asGIZCZM34im+i9/vBHFMIc4uO1JZS+IRG8WrCdhgLYOwQK9KEUbvAPJc4ISYlIF+bR6oUkpw3+
fNz81fVS/6TeqgGHgq3nwoMx2Q3tmrAxCd33AlhjgwWuHyEVwZx8UZ4DENzG8h6mPtfTYaqZJl2P
9tAHxuZacgxP4wVl0fUZFilkAe7vgho5pb/vHnnIwCFxUY9nNjG56wbCqevXUXB0Wjjypn8UbzJS
FdpL/mm3eJSnpeB6umU8UEtB8dIgZsRXAmBXuDxzFfZ8t7nZ8MSzmtK48Td5oKtLJVPYarf0p4dt
UmS+s9keQ35YIlaxe7JFnWUym8MfjFk89X6bYUFM9bJ4VJ3IwmorkjbIlsHiaK5DlcYgTkKxpNeU
kKeyEGJc2NrxzS5KwqbdyqHbh77T3ALEQ1P/4opE20TUlnZfPOp9bGm0N7YUhnxZU4MzfmCZFkxp
VCEXHXFpbOYQ9Qqtqr937Zg7bvjzVwGj8SJ9/b64w74K2LptH/X5ZccsNUf/QDnJnywP5Qd04PmJ
9sHE1hljhIaDWNJ+Tg0K9aPWxQiseY3ZeSIDsPKRt1ty+u0wvZqL1v++YaiWF66hxMyiVWp/3wod
sQ6M+Gt63C4K+UqkYDWLgH1y7MtCnMohY7MVomOBVB9M3TghG9lmqMesufTlIuoksgoTWTKrTRzH
9eUnHn63hTKvJdmD1j40CYlGXTmc7r2+X4X285qqf+vJj4lRTFGtZyYWkceQ4tLGADw5qS5rAyy0
o571+IxtKgJscVVlalPz57d6mdq3fwjG0EExHQfqtuJS9Hm/YLrp+JpWgmubG3V4UUx1mMjG0SND
+X0mDMqhzf8kl6WuGumTZOUrv9ninP3wuQ5k2ArLXkEY4MGG6JJfmSiwln4+K7EI5G71uNhrXd8g
Vl28kf5ci9BNbM8oa78qdYtVYk5LClstrJINm/Kya0dJquKehjOuCqWQDID1Li8yA6g/MzjbgTQu
OyRC4ixFiFWUnJbh1jslS7BcFiiDqwFy5a0ApCCPBTQ/uIqhMP0vqvQyxl+b77/adh7Xt8jKnP0E
UO6b+W1j0qJkqO1AwRvERHrub3xdnWeMLrBPzbOzq23Fp3LGawpVjl7x4xgMz+7sNUcEdRK4Gha6
gsW000AwhTbHBxS5pMsZwpYkVMBkEsuM5bU+L132S8bixuxD1On6yApZnm8SHZj+Pfj97naHcvWY
CDZU3qquG/2ZZWI7csnz9WUUiAX18KE/4oESeDzdgBtTSuOeQcECQxxXohaYX/BGrNoPpz1IYBpL
X7B4ntQEP6DlK/AfFFlMjpBiFlH8cI2P5/F+RxwxNnbhxB/PdwelcW9DKD4ATPfhXTTgfYRQKKJD
s2FUNwLufSrnwCXk0sQdITN7MjIrcxGJMTN9IPcMT8S5Xlb1L09zHvHWyh5bbIhgPU2wYj0ElJXW
7x8QyKW716AP7Bv3AAVRb9mvfnY6f41UStN/ZlfkR0AwL2fAS8ngWvTy72lsQSxsvStsE5msuPZO
v6Glmr7hKXv8VkvhT/hA8Ru7kEUALby5Te0rXBMPnbZf4EjWsSwRxkltMixgPo8+AaH7vJFInBu7
LxGMBVV5Z4+k0GKC9sRLvPPTJGtxaKONXtg82r88ji6XZhECBTEaWIm2tQC3OdRhAk4IXo08NhRU
R+1lyGu1mf7R6ZNyG5iLKwSan31aCFrvSFjxPrZD4WbfBI8FUub3rWSrbg6UtNWtLEkpgSl57vP1
YSJcYAaHR7U84spW2zGvMPBLwDGilrqC8rnKf7o7qB90pCYjsj6rujppPmPp0dM6m87GGJU670K8
NaJ/us+yOSyCjXy6KTVrynbpVKH9GV9SIbEAGSOBMoWeeqTUAzJ9E7KSpfr0fchUZUwDFje9PgBs
j4IltIsv3fHnsyhQ36s3pWRxYHpHZv8MwOR1RuNCUX+unBVXuD0xuZ0VolJRF4WA6/26XYmTX5XI
Ab+XRDf6ho6+HYWgj8S+vQv8nqEV1nIsyJ/WQndbLi3N8eR2dd/btVq0teetFoyj4pCLl1q3zk2O
o/ST5wnCQqqNsSC8ezPZ/+hbhrQLFiojFo1bw6ESHRsxpx0HBRrP/ZaV+dszaMeNxf2ebOe4AE7s
ioDK03F32SjpoF1j3TPkmyB4ien1H/3cPBHjxBGlf1rUYwEcPqyxj2qbq6RmZES83ivVLz32vKV3
iqK/gnYzVAriV27tj6qGGaA9x4XCAlCl6NUsGPciarxyFC8H1uxTLcGYgcjQIkkl9KSHNg+qgazQ
vUXfJ8cc9Fj8cMONv8FNNl6+v6g0ogCB/yheBU2iIYar8eWDwPUIP03brJSc9A6dd9ZqSPBq2Pu2
PVUx7K+cDXnMtCdG8Vk9KhI2NR4j2FFm+y1nYl0KSvgiLCjBgyPGW/JyySRDmok0ukjHI76X4GJD
X3/gZnbc4i9E6y4QH6UZeXOD5pRsAYHM8D9WP6w5zk+PoV3sMJjcX1NAuxI4+NGl6Gw8hzHm08mR
lC+fnFaLrKK8stJ5uiKnKvKlDT/qtleK9ZdpuRIOF6DpmER4aAP8SMy/W3sLZoKrv9vsEVq6aiOW
Z6M+iWPuAtufQlwRQHhlX4xmU4WD+rbBtXOFpg3PkzbRg9IaAej9Ybk7bBwe9cvbEM/rObkYe7ny
d4cG18Br7bg26Caly/hlFIyLbkN6OHPU5piBiwLaHzEXudwUV0Cr3u7tsST1FK3NND4HBEmCtJUP
M+WHN9twt2c9HgtNRgz47X9r28n5rylPp1B/QdsOc8XdCQE/3YekFzawOXut7JEi4fFCnIojIhs/
M4QwDLNOWlay/0dJt7Xd4m0H7jltXC92J0I9jh0jtuqB1qHngD8BpuJ6vHhnb+KKdWu/8ybwzcpA
AF1kyQPVePFm/lCljTAD5bx+Kxi4CQkl6/JhxNYzCkGQc+DW+mRR3hX2qaTaBpflTNswu3VNJ+WU
r9JKk3PSNKe6W9EW6vhcP2v6GRPvj1GT1jhX7Wqd+w8ju/5QAsesBv1Gn4FX7tG47w2dVQWSm0So
H0BTJGrPraqYDC/iMmsMRXwOFWdm+JEEftcK04Letv+nle9MtT11unSHN0Eg1i/Cykl/1Fw70F9B
7kfhrYRzL+esJ9bSo0t5vgPsH69+juV+yzfgfN9+oW5QTjfYngJ7YU1t+M2lZ/VCX5ZgO600vMBH
xnOBNjeK2Yh532hqwpkUjyST7NG+pbGZF9J/6quAaawmoeAVFzhjaTo+LpFD4yrAhx6dQZ1atAQH
sKS4xfb5zHtMdRe7ZtBmieiIsWbZ41Muc5zTbdsm7ueqF6qRWk6BNFY5XWqXaX/V6HfMdCgTRc8T
nsp26+7ZkuCdKevaH66k44k4T2IwAvLD93rd2qS+nQxUUg2EqUmXEKxw41m/JL2XzypZa1aVrXsf
uD7UYfWbgyHqDLtN/qr7UaRn/9/up17E9j4z7UruqUpDHGn+Xb1v34Ifi9U4m4N2hp/tZPlSdfIt
L+nBafn/+JNupCshKqgsdBM7WFwx4RWd0J/R3IQko7WwwG2HR4hr4jk/7zjVmU4QzqtT6R8OXKR3
Kk80FfhpF8FTxu3ZiQQJZQ63Tw2lbQ3/WaFVOAVnpoA1xvR5CPG1h4bNecfkUnClZsJRV/h/zSl1
o/lFcB7WJfSYGQNX3/J+IaWj131idQiyGD3/SNHdxPS5PjBdjm4rJ3ugyLmEf6bq7FCps1ZgyH7L
jo2p4eFsMMdo9xz17+GZbMWXH4GVUcV9w+uo58EHR54RHpAaPjcQWteHvxK0dwzvpwLJoGtIrdGr
Wzyp+UPYyHisRsyZx52BFwaoc7w59FXdocs54rwo5bjq8NollDszl04mNYH27eFodbR0nGQeB4mC
iD5fNSlZnJqPLjJEokoI+FusDLtV5jr5ZPTj/Folt2uNFaEhwPfX0/ByBVrv/4X00Kd+kjgM4bVG
xs//EdDRJEWb+pd9PuNgCJhD/jVrtbCDiDtUuVe4ebdOiNGsG36cbrhkUL2phF/vmZ2WxWpfYIV4
DM4HQLiDOUP9jFA79vKyXe16HoZ108faFTa8bRH+e4nIMuK4Fh3USC4kEpiHwu9okFEL/wpAJ+Bi
U3quXNV20mZZWPLjUakXxEHDknadUUyj47mQ6xw9So5CwFQdXzKAAznMQvXzaAgc2GeWRyJIwQQk
qooZEQ7vnz1lwvdxGnOsgLO5s0qpTuA2cpcjDsInPLHXP1xWnVoWfdlnA4WFaOSMTf0mhGehtmxE
Gl3y2iuL90iOPlmpw8UEarrY7sPZdbIA4jVs1zaWpjmIFJL3JG9R3wAfiLml7q6YrH1e9yxx2adg
RKP9ceAwYCAsZ2DBKfUwU0oQXRsvfQAPVuGY7gKh31EgxY5VqD+yIkW2bHp4ovhFkueJ0sIFZDM6
0SjAaN6pah2bYKnQEo6j8zzUYYspPcoC0Y7gHmVZEsMP21xkFeu+NNsLuD3DYunlQ3/cT70uNA85
5wUjbxVQSjYzI3s2Yep5OqtOuuZwjyfPgnR+YNzyUtZaf+9HHGhMdxEtf5Mc57ZVfl/kONpQMUWn
xGHyZoEoLn0Ck/3F4KXbQ0Nsi97PnTFuVEY7OMo9zK3ccfmNvgLztJmLI6Nsaug/BxnMQL1QIPVe
xab8pj1hzlqve0ix9REdD0Wo2ZF7Xhe8qntS250qWFD/KpdeLWubNs5ZjwIKtpS4PM5aBhsBBjL6
RKNOFlrr0uU9XS/il02PxfEFT96DYDMYerPpta/PILHbWiz3vXxSxJXRw7jbY1eBRhuK1euEUX7h
mC+5zsr0UKuXjrkRHDsQP8HsuFUS64zAaHxM5hEQVt1Jl57xrcqIdpm0w79zuaaymeqn1qOq19n3
31C16vESNqnGW6puGxV6y0L8MIDs/3buq8+0bXnDJu96GZSouf2gxDTMU/LBUCx29qC0Yc/VxpS1
Qj3mRDqXC6HLO1WcM/Hbspz0qcep09fGe9IcU2jd8ZwAQtUF4kG+WvMu0F/X673OeOrf6MhilXIL
laCmuNZqbiSmcX0b4Oj7vLuZh607NDO7zE1kQxtZrrDsqekLcMSgSfl8LNQUdfhN7krMSxvIUYHI
xMeSF9nRRRjZknZjQdha27InmvcbXWRSdYgQdHmVt8NlCHC1L4ZfNx3vgPIs2oNjF6XsAx2QYlr3
TlxRqqLWZxjv2kX1qak8xfvJdy5ay1WcG5XKXT7B061HwWfZkVIeFeSVWAy+KcLMt/AbHAz7qxek
zBnIH+ggqCbWXchJV+M9PUSYxiAk4nRZI0V5W4c3YD86uwD1fRiocTSmIDMWLevLh6Hhua2ApS3R
GtZEtXQE2Loj3a1ywKba8vo5WMqTYrfAgDyHgSbZFPYHKEE6Pl9Hd3fxEtwWU41YGa6L9VFYR7Xn
47Iou51w1HHGqzQfM18flwaZxt6Nz5Vk/xAgGWZSHyCdAaJa5+APdMUOr00uvIoJDMu9ouJ79ARM
gb4guLsNORePdmKlckPtOlN0juPX9T7cdJ9EDG5IzLNqA61gFrvE/a/L021RpIpRVD8c8QYEbKTn
CBIINvdJGnacQdg2U6dLlGLbqAX39+7INZiC7h/KmoaL2eIDbkpEQKXWsHClw4xmGXEm66N3frc6
2tRclrZlzWhIxjjKcK/lOiPXpCa3v/SFRW26gklzZuhyoSalBucArFbXnJVx3W1BXV7g6mBY7H2F
q/6RUZ8HBGBdqB5+EAIJA2LlNI1xFNjDdcjR++XNHCN6P/9uKAeiQ13TK2XRDdm41hVLPt3PmobC
sDokUbAeehcmZ6JrLch5YHRsf08U+BdclNG8APPnD+bMX5J5wZ2viIxcIAa/x1Dr7esovWQjdfuT
GChhqwOvu0xMWLWaxVEhOp+1ZA+8DV+5sHsaUdDTKW3s9bpVdJJTyzaZHlUdGGsW3M1dHyC2AYOR
Ev5+gWwiY/IPbw+DnIuMU+cKCI/AjIA/1G8kU5RWqe+EvKJ+SdHHyLSgAdg26Kd4p9tSDSWcTDZ6
vGvXIcaqvQlG4h4qlA5Iyxi1LBIe/N73d8HSOwstdQsyBrKWtIWElMEL3p58EIeJRmVyaZJYtPu7
SML/ed6QiNwPrbr+ZjaJvrRpochAjuy5C3rh1aDgEIiQo/sLHacXlH/2Mf8o2fz4D7ma953Av+J2
H4ys03zZiocBcKbZZ9hlj/baYi2RfZ/Rq1TXfIvKmZaGunrUpPCHN2YGKVaHtBATuRFFtiEF06jh
X21cv47r9gJqTWl1kF4mn9qWHci/F7S6jOCyLakjP8GY0qgQdD7EjQQwLPWJh60udImEbwcZ0In0
2sy2IZLmeOtq06LDkYDp5FnZX9Tp/XpaqbWZw1AHxjPFEOpwCcBqStlWu3htwV1DAJnTS1fI8ZHU
WelO+IFZSF6TNIzJwtcsrFpR3J/rFya88eZ18usPFhg6km3ozSQEJZ7lBJ8xldPmTF1fu6POBALV
VJsE/z64MwFp36vBgEfeHQxKeHyTaxNeBU4nbqwwmYd/jVazpgKdtSoUet66r6Gfp0NcYDpZDJQa
mX58GOvs5QcvllBkwU9cdAje2TtXcgXuXGuOqB+Fc6F5/g1/K9bsvQf15a+MhePKmIEihisZKJLe
739/ivEKR8kPv9XhNZGWHPMav/ESiWI0r2pHENrIUmkTZhcIo1o1E9qRkVZxOAk8oGYL1ucatU03
LzN6g+/Mih2cgWKfFRelPQec+i/CRZ1LKTs+A4YY0fJIHISwh9D4o7d8U36AD/2FjNxmTIjSTsuG
TaokWpQJU8+y83mu2FO54TPckRtcK21XBK2fpfjl+wzguP3Av/B2OGbSl2nyeVHTgA+L7Nz6qGGR
TmV2rE53159uNniheyci9NMzKpQud6p1WznEOVvMSmKhbSSTagMSBU0CpEiz3VLMD/3DeFtJ4915
yxDZudZe8TcFXJ1pPb6KJE0BRDWY3g06Bmtvumh20rUaRqAmb7UO79BwYHddYqpclqHihC1AbpUI
5BVv940f9okHVo5l8ByaWZfa2WIXjEI+f7nOVsJHztAkEfQY38Xa8smUQYDJr2ZN/cVWj1T1NQGK
fDj/DYD4wPFEqsF0BHDdPEqAAKYkSMpg1+da7K7Pb6TQjZ23nXT4AJsei8JlLlBgT5+WH0cmTi9D
4f+NnYzncefKeKcJ3DOCSuivBiLeDwlcgWq2U7wLKXKx03CmVpZEszaQ44yVYejgm2pID9PnS+J6
7l4f2q9aU7WxMvPZjT94rlbYz0x+PEOV3NfdAxEBZoG9Yw4M2ouswWr7tNyyrZ6PoYUHf22/k60J
HSB2xlfeUYOGbW722mOEkUxqoF7DWMPeMoGi7nwyaaBv53TwveHajWPji6oQ6jDmp9ADfbz/EU8f
hnq+fSB23LqiCe4nT88tYM1n+2AviL/7RbzkYKqawqVfj9Ltp+XCzCIdmUi/WypwlMLQC+PP8DYi
lqtC/YpPyD24vgEPhsg2qiu9HOdAuL08/e1ewrjZGIstWGq3/T+WkygiVvUV26mQ6qNlfhNigeg0
BargMhNc+8jjPeFbBUkN7JG8I8oZQ5AEWe1f/xM9MJ9AxCTegwYP8cMbS3eQn76snPj7i3zJFbAz
twBSnFiAmhCj8yo8Yqz3+8Yjy6YhPDsXauIT9Fna+jIXJ2/gwrJ1j+1ZqLh9CagvEIZBBsUftP23
WbW0TD9s07BigZYpsCK1jVBgNqVVeiedkCIpwvg5fbm9quXn6aX3bkVlJ7oszEl1pnN/s0akTqRb
Jz0vvd23jceNjywEH/Q2GxcdNQRMrNx2pQnc8h1/WQCuZ6dKQP59sSWMuRd1J7tbtnD1JuDhTiBx
uPITB9HSjdaz0eXVv9sukwp2gMCi7SVfT47mOvYLBadhDqq0c66cZhrBjWHzlpZ6f+OerIigm5u3
qT3Potlw5JnQYK0Qt/j5EdTmwGWyhU0y5CRje91CtrCw15nP59a9Yqg7VbkoQ6NRsaWgJaP7tzid
JZQnoQgROuh13mKLwKsNJrZnbRUEKfOmA4Vv5Ir6OvtNjvLKC7Qliup1nQfojHAGhDcPLr9hi+vc
wVzKczQpSwSU439S5UW/15dK6pFG2zrc9wZLisYlBoIi77v7ojmWpuocAtqKGWpgLvt7WGbZfmzD
1Tk1+sp2NvcohurU1OEJDVYNTzqLMfbnq4+ng10aRkYYIGUeyrHAsW3MSldO9u/olZwulSdTqmwJ
VMCsmcMYPfLU1M10teV8piedJgoHwAgTS5Wy/F+qCxflLq2AjwDWfOC3NnKM+cQMlnjR8/O9xAib
5np/7Tz89QxcDLK7SlsgNiIkrJnKvrn2kVbzlMamiWfrC84HGcbDa5uOm+Fb1t/npPtC/yOYw2A/
FnrP+ffBwU63D6D0bgtlayLQr4/hkm/3v4JcvSEFvkapWYnudq+HCzxGOa4EkaE6jw3Ocs0SVAEQ
k5EGDS4cizv2Zg2DPGPsxwQ/qr96i5RKToQMEVOrRyPOWQILUaTm8Dn3t9Neg+b1bi+23BdX5GZW
GsN7PRGtSDG/eVy+azqEUROTycRnatHQdiMB49VwHDXwNDCYfKB315rPIO+eP2fzT1hvtDvit6JC
gaFlpmQLohs4bBzvTzc5pZ61dNpoHYUNSbRwkwtLR4MM5yTVB3dLBGUu1dOgsW4JA6q3Umh4zC49
SzVcXCkXpKJ+CT6AcOztb62mXMJg1uMBZp6mPKeAbWD/iuEQarEWBfcdV5OPVbUGWPx85pJEWTi5
LukmjSsWS/kzvhST+B/2PyRTBoVoYy7WqahXwZF+oLEOLFJNFKFyou5yTpEkXwytrHiYmv9IJisK
mx0HvkX0Xe2RiE07Ovx+zoGlHDalac17CIgXBmgjt+wjGwheFScIjSYu/nNwdnt2DAGX1tjC/4Fd
f1GFJUts1D7LEJ9Nx/1Lqw1zQPpdP4ZdxICPoMGJY2Rw/lWFr5ugHGLaQgASTaQCWEV1vueS/STV
v5hYzpqmudvPcRkJsW/LxiLV3tEztoSc813SPjwVkOsgbBIyo8qmzGSpHMhHoDcft8XKnITeUSqb
aMFLqpb/BpXIZ2I3zOJOT0RmGATIdBbiffK1kyWkecu2/pwiY52aQgqcZm7wV9JUKzzLHl3WReaR
qHzUn6iS7tpMBOj2E5JoXqRLMKSEDwveVxVGxlG4k2OX75a8GluoCmUXMyXqfojglSY5xEH9/SQ6
bB1+6ymzefde7dQweBL8kT9ZhPTRjReOZzkrCwPtycjKgdsCCEELvx/FOknVsIZJk0M1G6JWKuh9
tFDEhPQbNr7Cj7avTFbDoFgJ54W2pyzXDBufsp3gBWPakz/1FRyUmj8K8EqKEnyL1M38x2TprPPg
RTcriWv2fAmfe5p79kofMnc71SytiXOOL6ww0CbMbE0hpCfe8Z0kFZisd/bT2zjka0qqbHf41yk0
t2VwdEoF4uRcs2RqnwH1RMykZzJYRq+gZEt/ShMySm7oQ3Zum4J08pQZY/A/GfvnvPENR68nkXC4
tSePVa4XIEAZBHRm9Luh2ybQDiMyM5wEtyWx0W9U0mRJUvISKJTXOeuDYlr1IZf2LP2yGytV51qs
GqlgbmWX+0aSDJ6G7uux9b/K7oh1FN3Oe5VbMUM1yFIKMCmHXUi/dQXkrLp4ok3LMlS1LZn1srnn
MXm7qbxWFIgMFOAOGnaeELr6HcwRd2ha+udtdrMf0cpLgBAyslA0pFeOTIFNThgcJsGObbS7U9rp
P3/TOJENixfy84GcwNx/duSMQ3ZcMeXhiQBCYKj8RCGfU5NgVzofEQy/hcyloExIJc5rkq/JcsVS
0t1wwwlgjwn1PSIR9QvQTYzbjGbIMRHUkQNLMJUq+lyVcDfl1GIUvuejj8TURO8ndM1+88eHoxKd
GzTWXqiu4CBtVzf5ipCO4/B77ugvhOOx2FAFg09IPKuX/nOIi7ViRdJpPcVvlrzEuzFCX+K7tESV
QpvF05MFh6ecfzbvlUsR7a/owsobMm1JX5eQqtlQ0NsQb/DHwgIhdAOPJOoiF8BeodPT3YaV9Jpx
qi5/jOIqTe+YyBMz/SoeNO3wpz42eBMMS4P4HS0iCQZ21ZQ122dt6xgNqIGjhoPS623BX1598ppy
uwMBzZxNhnI9596uUbGsRVh7SNv2O6bIXFLFqdv3964jjqb5r7bF6DbxPNEMgmt0vXedhUtoap3M
rncijLe6Sh2He6CEmBMgPr/W5AEfD2XSfO2xC6xiY9iYodDokSn4/I5D2dP9HmYcBQS1IDw5W0tX
ccGaQ7x1z9qDkyP+nTJ6dW6lM72HvYZjkntGIA+QFNHLdVgkKmjWivOFs6EZMSbeCToHmmiUeI8b
rimBV3ggs5ZtCp7YcpTD3ZvhaZ6ZwHhhX6iQCs+3kZZHOq5tniv/9FBXxBiQcpGoOJxwQj27h1lA
tzCd985lt/sgZ8ABzO/6i59ImW/nQGeDdZd/NDYN68Y7FkdzTsTyjLmAa9p7vWiPWmo15y2pKdd9
5SIeTlUD+z3th16c34mMxQFXaH9PVE8K/Tw3QRYeYW10COTBFtAkoEBD8BehuB7guI8TqqXfEU4p
2U2Od9fTAoFTaTe10snYP39MxU9wMZOXX+MrY5QLjaW/oS3KOvxZcTsSqdlVf/GUUk7j0/E3i7Xg
cff3J+uvvsi/QQ9Qlp11hh7Xsx3sY9NCjqE1alihOqwtiBHdkIU72UsvzNYgWC9Q/9jW79UBtVEJ
dYlPAXKWTXkqqIEoo1elgLi3Y4eQWq5CISRu2c+Nq/7e66aRXSF2jaICAaZUIk+h3P20OraqM5e4
UiLXDzfQEjiqZhkm8OZHlEO/Y7d7t9dqoD5sti6ZlvM5Qbopt/czDhD0EF/DZAGC2cVoj7P1It9a
crym4Sd/ZNRFia2e3CwBI6rgG9+HFMsaMaM2oZDNCLc+jrldCKOg490zX1fq6+9S/lEFOIddZ60o
yYxZEJVLlNH8HxONQGQsknHFtC4kT4sR9ld9Rv9qdmFzsxnIW8LJ2Np+Hkv0nFxQ8ZanyLet2KC9
ZEazZatliRYwOrkkJoPomEfIyccUaLZJTCV9a+bo5q/b8ePIzdGvMdGXDQRFyMqyi9bYWaUkpTwf
xUKxkm+RhS+JlHxlGeMfwAIzZerddkg9BMzMEPRROVhs6UKE0Hdo69ZRhMYroLDTD9ALzfu4gJ7j
b+OPlL3ky2w+3S8PEAoSDYaAivx07a6IcFMQmoyd9v1vSmVibZwRlADfwH4tJkmaE/xCMvdqdg/6
FSm/mVe/pwKOf8TCb5cCskNG01rteAyp/MdUoRWQanC6NdMDhBcNNhmv+aOUZxca75CCb2CT80Wo
v+TeWQxNLNRW7SXksmqf12Zv94uzZ+MDsLRrVlLeFPCkRAuGtdJVyXp0Lq+dWtXGYpnElFoe353l
ucxkmKKCzFn/uguWWpL2VcPbEoflTQXg843VtajFudaVaMRsnqAjoKgyoCakNyWXDTkpcMhgGNu3
4QO26YXUyYD9hc977cUSujHAdNZ8rvKKDu0HaEEeC5Jgb0Am8KpEIOjnwJy7AYe9GfWJYjTXEfRj
ivWmgxxqatb7asKd6eu6Nec3z8cDu/MFKyN17/K9PvSsof3cG37j6WqlVzRIrDNC1kVUkfjIzhFg
NUTe6Chxxg/JZet1SRcBxEMoEBn68rFzk+Zz1dZe/au2zSQo07qmH+wnh1s7GaX1PYAjKPGym6A4
yj2CFYWv2qtZWAYCjZMQlD8LytzALVmOX1YfeVqj0qOhqqf2vEsolKJmwkQqRahgCgZADVL/IEda
T2h3tKoYgrbgQAASnuMoiMQwpyCcNVBTOxVh3EkL+IjxJPBYNiHLzEA2p2LsiXrQ94yewWEV7LSM
+cESY0LHPuNzdjvmdh4nLwyNDJxyjr8NUSGD9XZgNNohKdoqIKi9PkgY+ab53DpTdGRHEUy1z4iQ
/q+S5iG+nRj/c1yRs0zPDbdrb2geU0Xihhq9KI12zRVJYGfqBXAScCtpeALF++yz/PU33lsPSHf5
o+/Bu23kWe2F+/XxO/oIupRTDQkwA1yH6m8Yu/XZtncAkXdKQldxWntM2/XNpocjEP8QWvV7tUPK
xY4YlnTZB2aY9H6Jj8BzslvXxxHyt81H+xi+jWpzxqBwqzJtS7/7aM0dJ4cSz/hqbpTy8ANg3oe4
/cmg2WRPh08D9glw65pAF9fjVJ3YLUpz19GvxgFK1Ujqj/Z0C+CEpphlexr6leoM+Gsmz7R994G6
woxLsa48pL//2q0FplZg6YU4ixBz0YXVDEEOhsdEB7v/c16Z5HCrlQ2GA46G75BUzpUGGcjXOuMy
vkgyoXA2EWLfJnhY6lhOjkwF78BL17iHCkPv4GcrR4/Vf2srmaozuqwYlmVoAMtFf118TXwgRP/I
I4lNkhjpww8Q404xsuYjZp79hyyYoixabVcSMrydq76g4uLh7vE20TfXaT9FUlPFcALvcgl2iCU6
1fpUjrCvgdOPbILGZ50K+zQrZ5o1stw95/Wx7CoTpE26Oq0yaVwkRwQVT6mhXzG1/0LNDwa/GCz+
k00YgOTtd6P25cSIlnjBy85jgBWV+xyVySZoBw6/ZINplUlZ0vPkzLSNETYW90hMgGg+MI7ZkUkF
OM+kyy/zUB3bhaRzpm+zVJCEx2lqBCcS0FppuGpzWmPAiy4rsANhEKBx8OTQUYFeT7anIBmtLaaV
4VtHkdrhM1WR2Io4pnDZauJbcCtYDGpd1lPa5Vr30TX1cll4bGJ9hne0IQgCKHDFB6rU7LV40P8f
p3HYOgmFzDsoqFu4i53/p9FhlZfVnhGV4wd1J41s50Ef6c/nwlBJq1b/+T8Fs6eqd7c6OtqIlb9u
Wdx5LCOYQV1adMIpfPtpkyz+nZusBVRVXx0lJjrlh8GjTizXOktN+yDoepCI7dMpkkIQAWv2ETIf
6rK1Sgqm/Lz1tPRhZolsCUPPNNNBLF+NhtfRjZQK9EKgwTs6uvnjs3gEqwvETB+sSAe2frSioBZQ
YRCBW91gjpR/SsO9Qsh4Wy3KwMJeZGMOCkbHldwtEMrpXbOcvG9zU6bKphJjJIoGbpFm5szfW+NM
6LY64YaUImwko0DFIHnGoH/F737KFH/5KbEGY79HGlqUWzc0QyGAYEdsjS4QkwkssBdPyvQkl2Zt
5qyLglPrZoND63fXsNjrPvpTlEGJ4dLDmEW3/y0DxkWqbnwPQ583alZt5ksAdYM101bigHOqrwC/
E6024L8SAXRZyt7rqS4tC2rTjXxIvJr4mxwCOjL0FyZj1SvOxk3RNDYkeo0q4GCUuP/dppJP6EKq
04qcGViSkhiaH2peBPZ9U/hXwYvs3fLMBSD2kFynuOmYoHVs8neNBt9UVKACiiTjGQAcFnNjvnMs
aStuBRv3FNP3fk6dvryKkwfbFNBSqI8nawNYWTztiPG6188TjYI4pmlKwG77X4s+av7hQixSOJJW
rMQEF7uPnDfzQd3i4frWxSl6BM7fggBWzfk7A8CsJsiAPC//U6Ok8/7p7apHp8qhvsvoZKQ7ouqt
2UImvFq6rLUCx1gNq+mPglPnPrCWfAArhgPXeh9+pUXTvWMthrHCJld1u3wJvQs+z95f8gpc1Liu
BiqzziItip7C24wuXHW+Wr8pg+Ssxcwy9qryksDo0ha1Xf2mSvzbZAb6/7vfGNQHRTZIny3WQpJg
zVPV3aDUyVfjPmmK3sIdYdeiCNujl7heEj0iWlxwlgthRKXjkHtp+B1wl/mA/rAr5+70LT4ql8zu
5xwqsrBYQKanGnbct5gZaQ6AiQN/KfMN80uX15Drug3quj7dsd5YXxf8TgshmGCUGFMYuXwRf67w
XYU7IzFVf9v0Yzwdbznz2qE/PK3h3shF0lM2MfnLtXwxBbjieb9ByA1p8wBld25xYCysjk/jO16O
7JxEK6FoQ07AQZAlYhYQa255sLUr+4+jzN/gXN7dBM/zQ6GEhgPONEzaD65phSz4ok2xiXDv1GUA
QLND0NadieSIUKygQ25HvXkRzL4ZtJYxf7fb+9hbN6pK0j7fIR7rg2jm5hlShOK9D3ubw/PXvpEC
9JA63EQBC4RBVUyPtXeF1xvuGgoKEXG8cdYJmNbK7dDpwB2FLmgUq2h0EhlLe0/342ucG9zPhO/H
dfUqZ8vF7zqMvgTVJ4ZvK52OyEndzQWbpFbXpotl6XqHKjv4j6fgVeYAJ7jFiiRMMrMWMs894oe/
h+9hyqIdw8KYQW0EPz4j65jPaB8tYvC2SjUie9M7G0xfJcs6WPxToejnCLFBlQMbmKZXO4U1Tb1x
ff4IkUJ9NrqJkOS9J7BkbnR41335zfr++kG9Psdw4HtLPJSn3Gob9nbdrSZVuLC8kbg6HCa/Ozwt
4vaRkVYymLyFXgErNvKq5F6GxnfCqFQCbd6YsXuf9ZXNCEZn/JfhTJsxHbEBwjyMWCRnNPUtHuir
LAq4uuruI+PJndC3XXEqrOaP1tKFEnINgjnVG6sokZLLg359fLNN2oEgxSRZ+wO/tMXknS7y4M2d
Sbdp/NmlEItkaZqbs6jnZuhDwL3Xf+up+1SAOhUSBjotF2FOMoTO2tWMDgZgDUQea/Aahn//DZ+c
028QVsGT6lVM9DoIuMsoI0/1rueadaK0HjDKJjsfbkxeHWpUqIVhAW4y5JrsB7YW0dgtkcg6ioCx
Ldi5eaMFBe82YekjrZbpcj+af2/OI8/kRE/9fsDcL3+UkPJ6rD5KzQajM/Ud6Pgjq8g0rfdrhy0R
1ixNtC5G65Eb3bMQ0CqeAeXFD0lOnydWFXlNVEcgcQgV5Y1yKds5i9qUOt3qDZUfjo/IX4+6VK48
6Vi2iGfIHJuIRJpY9wnuguTMIEsgJ78rxYbz1ZEwwpLRhquL2D5mTOSJhHQ/PWzQbHGvjjOWqiAA
UxZ3huj8e9MuW8BnmqiuFuFUqId527rmFKBE8v+TmtEKsAuSVI4XQ4fDH/AR64nkdrrtlX2yXwTv
2GOShDpv/BkfixY5GZzwiedfzWL3+T8bVzISgncGLAoYLsEusWZGObK+Z67jcvwC45K1p7WV6+nY
U7jj6vIqn14CPLdB6FLi44UmOxi4BJSm466zKsPWUHqt8d2CJfAttdfeImZGzTKTksAo0j60REPu
hN5+F7aeX72gv0aPLrtSIcuscSAXWBo0CNEBgr3HYKFkI1k7RBMqhhOtyz1DlmkGUAhtYAbBC+Wp
c3G4nAtiMuqR8p+eUkM2JMbU8zAL4lWmQJSWm6aRMSfBIr1sHu0QxinTJU8oicCixc885sPTqBdK
uiDrUvE+lmcR7Ulw22FUP+1MjPKlR2RuXYPKBmmwkZ6BMy0RQ+UOR82BRHlQmEQtsrCSYLLyFEKX
0bXWVDaTQo44cpX47wu8SFPJlJEaXbkKzyE2fMjakHJTmJ9xXYHjxRZyNg39+N9og5JdwxLHz+P9
6P2DFZCSRjjra8jKCrUcQ1wenfJTia9jRDwL/f/FydoHOp2TitKmKYcpkvCrRS1I77rAqK1pzWlv
T6hCYcqgfUp7reMAo0CHwHP6Kfg91T94eugdywHOEKOFBUVEMMMYXQOBerXCjmfxBe5Cp1LbV1aD
cueISyWUS1rCVIQXEWdJ91cUPQ7ik+nqP+DhokHWRi6//aF6PEoKS1IaFiKWA6DHLcTDnUJhp8A8
JfBsGqvtUhc0zvJIvK/PcsDSQBnroaoAHUEkqcY8PU8rRtW04EQ3IikU0ZRK3bL1yE6RYrmIl/n3
pcn/iW1PYKXBd6ERta6Z0UwymBo8nWAs7IXFJZ5MzmeFJG6FP8AhbolkpYi6ucBM7bT0VSOKg8qM
X0QbVUotFeCgXhmNUoJadlL9flKE2SLkY1h3EjBUU+VhmKzreYA2H2PwuzAQ7/xGlDgW83kfEwxq
WOszrXe3rG/7yimQYWpt6as27Xd2TtNgbgVeESFMprA+tKydHuZrMrQlvhhz9WNF2EVauAV1OyRU
XRGDTalHBtZ5MP/xH3fwkp/jSRcA47+8yoIecu4sPQE4QJ7QFiS3iFgMMCOoxQb9mjRdSX+BHnzI
kaWdiWDgQpCs2d8U+5N2B+YbjYM8SkWUc+x3nh9FucrKsvocGNotxAZMMWmTYRbf8shqsgsRJhSm
5zAJXZA1EnPEeZStuQzGAP+CZbc0cmwBhZztvOTLNHexXc9NEJ9EZYgu1aQ9M+zC/wOkFYwNZP2x
xmDsdACKNFHgoNxZsvhJ14S2grQOxf+kRqGf1+2+RT6zJAmycmq6X2j7h83ouGt5DpJuTgSrb2QA
uMjU9srUlK5CY/WA+i/qQSmGq6/V1KO2g4uzDv79lMjDXQKCVacNt5Pay5iErT/77Qq3spPAl17f
Rd8k8F7n2Jk5nwKB4oaTlJndQKKUDnCmogFRAUTTcv+5k6e2fFO6kGH+ip8+4+WI/Ntq4swnmHJD
NAK22Gtk5BraHMkaA+0stD+/AzwExAHMr/VEHL7aMUS7zc8RGeGlaDW0XAp/LT10ePnSPuC3n5HH
/2nPLDUmMoxIjz49n9/TkWKqJ9JdNfH/w6fmXRdEPnj0vnKJxU+f6zJ7fm1h/4/x7ZTzWerjYJIl
q+qEr4fP53VEFWFHJwrO74GK2bgzMP7dMtrQAolSmx03MWe0lyGaCEsOzfU5r4ItAPyLIUz14K1I
uG6+aBs2YZpx05Ct1TS8SIUCh2oa0o9svNnxH+zB21rdWoPOsGN5Ghto8/MFwjPLZg0LXitrdWGh
a4HBKls1CQWusvZeOh961z20O0oHxrExX0TvQM6fLpi7Cpx2c2Qi6pLgjzXfdPuwsw8SH9ZEsyPn
AyRaa2+zfq7m3C+Lczyw6Vt/oxDtsKGO0pYXgRNcHPm133XwYVB6n9jCF+kJsWCWM03JJzFHATGS
gyPE6iyLhYpjignnitYGN2tCeXTZe2AfKu1SjFUIxX04rxqQl8e9vw/eKnLy5nDmQBOhCC0vpV7W
FHdqFCurCBeUj4m5ryMZrLUr9yRGlAnlZRWU7Wy65Vq4gP8L1dIc+gGUYMWUxLAJtblv4bX2QfrO
Fd+Da1YmvAF+JDf3F1R4SrWICJgu8mhfLIPElbWLOAV+5HAlK9emQIkuncaE2tX7iWfcTKIjy3nH
mGzErVR4eFXIvevB5JAL4h5FdtOFICYxbYjHF0BCl6y6FvKYgdeL2SkcEBHKrkRG9iaPlRtEELyR
KSYbT2nR4LwIL0/YjvT7lwZqrKpIKSuOWIql4NmEqDzjgNd+z3KrQsH50gB2ZJSYt2rFvs6u0hX9
/ihhM2MNb9z3oKAbxDCpPOweJiqblDNy5oHinuAzcLwIWlGLQX12atLWxe6XjMP6xrSYY1V27yAH
NWmxVAuwu5mEHunUQ1mXRsY1HSGtqgo/Zszi/jKuOE/RZgFJayknamZNZx2w1wa0taDg1DQSDLQ7
iBNROmibAHHbmiDLq5ephVQ07YpgoexHvnT7pxZvd5jIbMvk9GdlBPt2fX+Dh7s4udzBbdp1NLj7
pJjoYiJb2XKY97KQfamX6c7DxTYPKmQwfnnbiBV4CUNEc97eaWmpQmK2W0pnpEoLlpkvEv0CI4Tb
JckFP/T53Q3eZ17HsaXGFJLpy/pkkzySfuVnPcroknZ70tUoiubwwLCnGyLXmLgKN/GUnS652ANW
xuZ6KVJZaOwaUzyNvI2HoGjk3gJdwdU5/yMC6SfsLGD053Dct2iw3xNMnlAmeRpw7WjAeFgqOf2h
q0pkoSLZUGLO54ZFCpJ4/ebyrY6X3t8eh6wvqT0iU2A2vMFOMWazmKrd22ExhFA3F4alkR2FwTWy
hrF1+2IDxIFKNeATz5JCz2lCvZxPNSDom80up0wuf2WzvbILHFDN5P1UmO1aR7zLCyEswWxbRU5N
/pCWkoSwg0Il6cv02jcM1SR2h4VJPCKLGRgo2dSubTKopnduZa6ipgP8TABdBKdwDCABotxgPozg
FiyQHK13GK0HQ6KDfeFwEIwy21SNjWI8O7nAoKHQ6OnMkjTdChwBSX+zpJaKSsuc5eYoH+uSF7Gu
bql3yMG7YcD/04W4uYrEJtvCPg9ITfy7oZi6xY2edH2u9m/hBNlmvxPXWhSdsoP/DX9TidRzljsc
MNrUvk5ASkbG7ILOknYs8K2j8VqKluhq+jChvxbVhpjR9yx+69wtDD1sQWVumhcwCcw4XgQHulo5
XfYa3GDkWUguWXVgQviZCfkHddxsauZMrnF7WSS5zSrV7t5U1hBtvSNttIGzrKMjXie/hyN5ke8r
s/sXq7y91Q2r2Q8lF8lCpmNpLCO1If5Wb8PA36mDhkLHM+bYzP/RPvELZKUuQX/Hnn7+z2HYVEry
EHCihEIm36BT0LwoHa3b2iWcPgJGrZgUYENrcIuUtxyHPISXMDJVwxqfS9GWkripSi65nvfdbw8y
87oyvIxr0mEokAnczhZBcDczZhnAm8Rtvt7wh9tCepcqk/hSToDk/Zph9MN7o1rciJHK2LrS+XIM
oEAtrMAwXXZ/OqISp9VUkZAXCrA36u7M49rhyalQAFKrMCyoHQg7ScQfji9x9GDDpuVJN0TdCHo0
j9MSswxFdirSnoLGud7o22b3uhEeqd4FCW3+nyt5wJZlcVTjqoFtslKrbYkSVfogsnFYFt4+31oD
UqgFahiihpy6qyuoHqTTobnd5ik1yISh6NUI6H6v+aVzEH5xvil/ihDhYybwzcuaFbiqjBvw/0dh
bP25dph0g0bT6OrxN1WY0CtEAPDjQLfgraXsr2YEsUrQxm1bRKQcAhn8zeHrNTaLslMth+rzh90E
7P0+3tS987J8EdDWLaUl+3rg5eStFx/hLjgat6YBMIlNJ07tPlV0ud94OuE0OXBad+dX+x+9KcJx
NhxfCrozD0gxZREKNAy0cPDjeWMRZ+LfGCLhYnL2363PHEQzllhHw5W+U1whF+gz+lkOArWmOiWD
9iNnwmKfBAl0tMc6NbdgOO/wVDoZfVyvp7ExbHMPiECSwqsCI87OOzOPQWsf9e2OtKvmBXwyXgPz
RzB4A+9izRZBQfxFRJbbJBbmcA5K3rcc0wLDtIX3ePDOngUfUNhTsuJlEQwUlMOGU/zVONxLa1QH
owtwFH44QYgyIRv6rwoBUdTLA430SgeHrJ/7QqErcXBZT1CpuQbYL5drKHBinzKAZgb4ul2MnQJ8
PGFgtuA3sclnapQuWT2hByweLe7rbshW0Z7srdskfwJm8WceTJpKhIkJLssJsdvvQOsmXPWPMsl4
KoMNzjwnJb3er5d5N1UOYp/ZJe2S0LzfeIZ4GbVOjt6/59sINjdcECIEFOfC0grsu9PnW89If1Pb
e9izDwCMFIDR/nlYqe/ag+GyvXR0JncSoEmU++FmaiTy89YzuOacedFZcAo6nf1kr7LuEpE0kQtL
KMKpPmZMUG26AaSUviyl+C3WEzJk+EYxI7BWyE8KzW1kh9FIj1Suk9OzONGvTcd8vSlhi6ztxi/l
cKtB3sgyAIFMr95Y6tFSHKapk9M9hyEu5A/UfoLmEauvwJIt1j8QII3hDynXRo+LolMavH5Aqnoo
zm4G1zpvKNDeFR7vO2EH6SLnVXzIPOlXxpD/luFI6hRg+ed2ipGq2JqctN/sbSEKQcB39VOr8fXA
dj29DffcPf6M0n5m9u8MTdMKkhsjsnh/XewC3+IDnQVhddnwr+cqGHYAB0kU71eK+liQYq8/QqFi
izDeTBMfKVLNbhbNqllNHp3icvUcxsBVDHtdS3rE0ZRRh5iWQ/IuhozS6KmMaekIDbSgPnaOq3yA
2Hgmj7IB/ZzTN29bYVpmykdrvloaCwBhaD7JZlZewU4Ychrg3Pr52L5KDauj733yrmqyt7gxM5xw
qonyM9nSYXsV1FYcg3mi7nwrxW9KknsbHH9Ilh/unm4cX4UgqJpHLFsdBKnVe9K9oPab49NnbVkh
cAg6gaOOXkOAiD48Pa5DiQE+Vo51Xfh8h6xlk2huACy9NmKDJjOYa6MNnddABoLUgJymzqlGEqon
bJ7Sk8rmcyUnkWdSz0HQfy3TDjTfaIsuIxi0YOQfVWrJkOEIBgu1AjZRfZs0erIVrP4K2chfWJfE
+k4kSIis+nhTPgDykXNPzUrq3AoDmXLa0e+7t8/Hij1qFAiVlEh3PoBNuo77ex4scKlPU2IgeaHM
ciBPT5QviVCJo7TmAAPK8cmgw73GMc7J2EuB2hJJRlniIaa3d3bmLMPTaglNz3DdhMwOHeY8/QSI
wCK+qUg8ZVlMG1C0KXUi803z4QoISNxViGl8kirSKhRcHN2N6z4gvpuJ7klmhIgEAARnU2uPWTIH
Z4GtjxgeEHEEdxZ8RwPEGEsUF4nbRB0saT1CrxWuX+LyEvb/+4i+p3DhaOuQ59PK4PX9icVQRIgn
6djm0VX9FcLDQ4o0rxdZQfyyWitEJCxOc9y09QsJ2QqjNB5hI3TX7thX+I4RtFPRU/7VqCiuMa2T
53l1j7Vbh2zXzIyotfHvfJyUiXNfWSR4y/s5K/qUmeLauX/9Sh/rAaTXIyP7NrNKAEH6/qjLJsYU
eHOZejMfqTxOQPMo5Y8if/Cq9QlPjdUWPKbkguDuDWJtjlFGkLEmJxhXmxhYFL6fbW4S6b1/wfhR
ZmOzQ3X0fUGFCT0AZ+AEQ5QU39E/z/m2CQPAHUHZBPOByMDgy9ZKlsMNMzGPgCw5vyPJlFH1cv2X
db14sSAnSZaA+yWKRZTKxiJqUz6y5nDG9kgqbNDAg8KZ/8FzyjK4V3e1XAV2AqbniPXbtBHBA0Wf
AmPHoVpohBXqZP/wPIpAjYetLeB9bNUYp/gDaCDDSpklRONm/HhO6vh2iWFClJHFuTc63lJAyPWy
/9HXSzy+TLT2UUDlPOe3wKJ2o+mlEApoYFCcTE9AO0VVTwCWidu8w07WifoO2JaU4K4IzhuOOxKY
RtvmHMADI+vHYyZjvqdCbNcx33QL7SJpDyhoSenVH2FQaZhNm3ns+YMFj0G6LEic0gUxJJQ18nNh
L1qaD12+1XWYMQ68RaQWBKj3LEpqjtb4/1IYxzWIjKAtgfR+Wfj82YPKYILrE1gvBd0k6E5gn8CH
MfpJMSKpcGws9p34+PjvlI1JMSRpZUnrWwlP38zCwip5s5HwH8bxau4o99OcEsq49kGFO3C8Y+My
YFWlITgDXVIe8i2kdKqD/QFE4mV+rNy6q8HcNK4d7bQBaqOC0zH36Hxmz9k+OjsENUtQcGSWOqzB
PGKQTEyWKjZ10ScZuU6dSbu3DW7yxyUacxvS0pvWw7Ka/wT9eGr0EVvbY3QGA/8ZQSpfUrcKOKI9
q05xAxa0BoD4Cx+R0GBpAA/keQwhe6YAfGreeT1ZoFOG4PUpCLkesz/38pULOgHWbOrCW4K8OW0k
xaAoTyt22YKCu7OVP3HkXPo1zfQENCaQVJZ5g9PHiStVgY1ox7olSMYv90sHJIzoHO4dtGNX8OF9
wM8a5avNAoCdSCxoA8NBgJCYx8SRVhhRYdCIfPcOIHQHxlIJ14wmZm6eoVxpY+ceh1hjizrLfnsE
r5wgRaw7IFI7KEYT1NVjCWvbrmxG6juVJzFJPQdj8jEXVOKSwRGxEliFQiv87KMsoTv+BtF4tvjp
mCwL0TowO/fD/msvpjO21gfoi1U1eeYGKtlw9UJtN82hSlZfKn/NyAc3dsNpqxp5r6yno0ngvGOK
9ppjVLqiAlwTxcUADPqFi4oppRY8gMpWFslh3XagZJPNmOUILsBRj6/MvylcxvtMokDo7V+ww+KE
KG09QT8qxRW19vlabtp+Hz5W+P4KkVtUAgQOXhklKXuCXdhwH3KKq0QzcBDT5WpxTXEBJWQcmw2l
k1Sj0QOUo2O05zi1Ax1HJNUIi60QVhYNapJN70GvcIk4eSMakNfk2zi3pcrrJDxWqwE2HXT9FP6s
/DViHxuQmU8uEMXEohTMg8QV2fIVVcSo3xw8TTQCp5UntiXBuDALUxFbrnJ/4TUw46RhHeVdc+Aw
D5ceqqLq9P7gH9GCKGvynqkmxzWP0G7u26yuRzSYmj0eDAc/sNBrJxZVe4CzSgBHbE3Wf80E2Uon
WALLTDabGP3YlYFrjqme/KMUcfjhR76NRhqyXtNsfwGW4NxS/vijS5SDFdQU1hg0ZQ0In2zd2JRP
WoA3sc8tNEA4T48Kroy3bbIymboSgIlZQ2gXUOC+n3QKQQ/MZX7mUhAm3YsNcHqeQNTglmt+rUUw
qHlaRKyl1tPDnlDf9mk/UCTT3hN+24sseDJFQcepsTdwhtWEDqztixy0liuZh8KOfRgjtR0/d+qr
hd3LooAK/Tcrz02Gi9l6cfhl3PpQKN5X5q9pXNpDJKkVPk2afA4j09uo5a0CAJtqxGEgsQiVVnAl
ISZpsJUgIsWtwMFQ6VKpcMNNZfyxs096YNUXbgqCKT08uKffW3eyHONoXed02QKQsFgaSNTeH+5L
2QWNYXyFVbSjoU9vd/fhwLK/+EFQQMc+o83s0hw/dpRSvt3f7czKmWjATedS2qkd/L7Dhh6IHduC
HXes4gdDRSg4Er+DmNcdqpngUvENNkeViZp+2e5qpoYxL6pm8BrLCHDCkqEt+v/FPRWN5IQ75qrP
NCBRFMMxo9d//20gu+ZMCjTX8Q4VRJH3keE6C3mE90JoBAqcEoe7lNeZrXuQvwP2sq6bb67TBnD8
NTt31Wm6MzJLehGYrfDaJOdwTcGMzh3YCAaztIIDLNdE56hjnjXiJMBF4lsFNrBMXqpSwA5cxaEg
7ZTA7+IMFq0ubE8azMSFf4xv4HIfjvdZq2p2C98W2TgfecsVQGgsmLr1fAawvsiufcJYtACX5JGP
DyUbQTNR88v4Q23gsPXa6KHePbi5LbmdqyRln/rxPpF68Y4AmURb5PjZ3y1qVDqPJW3cw0KveYkP
4DAIHLIWoEfdFvec2/YqSlMa5z8kJpNz5XJZ3yR2551OTJUTHITNEXsTOPqpgPjgk0bHkPP9MXkc
lMUAd8OhsguwJP8apXAl+k3J/zApdGlETsJJUeteMIJVIriqTBpK6dbm2ZJUrq7b7Ma+me/inPdq
SSjPHoZ2iGZpiQUnnFkKmdILz650Unkkg960CrBadjVAEShymoHmOgC2gK5ZkiTsWq+4BeJ0/l3n
I9sx4lrDYirbvN2EOisHdgTJj9V4lyVyCNEyDpU4mFMOzvwXeBAjRRlGj6oSknbLK3I7U+BrtJ8C
pKXvEgiSjSXoTyAAZL0kJq5isLiiMtndymgC+f8UDK7YLK7lNPX6QSMIGX10c5vHRMWzx4prNWhb
mtLCvDXPQyPj8KNKaGxKBe7qUjaJbAn8RxHiX5x2VZakYWQhh3/o1+ZSsLj51Pxw1qji+G5YouoR
QdNSvX+bMFfeXvgWcLJGriqsnwO4JU3dh+NvFuYDUEwk46x19TxxkPtMXpLLXpemvWff1oj1+1ee
bxSD9RZaZxNwpvbkYzig1XfxO+YE4x0hsqt3uQ+S0mWfAF4v7nco1HuM3Z3/c1msNIOS/7oqDlCD
V4Lkq+aQcOS0EglgkVA/8468BBR5shM5L4SPYp4NsbNOCzu8jCKjW7RVrEN9S5lpCuZHqfe4CqVt
ydBOK6CeqdprV9WX1sfuUztX9Hl5Wz4s4u3CoNX7pAWxB4BgtijmHw21cXrRTpRJwlnoWpZcTfnx
vmPNWSJHrWmp6+mUlP5ZhvxluR4tE2wc+2mnzQE1LmeQdzJBpqODlm9wuFIb+8lzgJo4jlQury3C
YdDAf12JMunxeUQl8RyJEEwmIL/R4ITExdb7tpqsCEaGE0qiWojxLrEMWnFN8tLaIr8ePBnUos9w
y6XSLZdFrbFJY/B+4Az0TEu7HWXx8rpo+vpYQWbda2iU0rWZ1zHq0f/94DEXlsA0yVlfuVK6KU+/
d1dh/pRJmkNQyaAxhvjPKrDL69wJbbJ4fmdQ59opJH5LI9AFfV2pIDW96Sp1WAqCY4wxswsaOGuo
xQQyz/8X34fJW3uE4fbZJcuyKGWHZLx4NZ3vxx5YRdgPxR2H4bRSUnSlom3du8Af0/yMDUOcnANe
OqcSPgrPbFlrDAwALEkVF699VH6p+RZTroXnz0WS5Lg2vRYDoSlz+94yyCGdWtoa+s1cxTrx3SXU
dBABYtXfUlZAy+YrqfFIxWpYrp33nel1GeRqp6+cpU+oNjm3HDi44Onk8b5PWEqt3X0Pl/b9fpIM
rzQ4Zbh79/9jOLQc4/c7oz1cEo0xvS3RV/k0cLgJxoT6oSCmwqKo/79z4ZgmtCkcHplM1CYdgW0u
ESWSwP7pHCSfzQzin/m9JzUaFaKY7h+5IvCow8jDiXxSPfm0Vup6TRtvlXU2fUVyoPq1qMVNYQtG
Jrodfw7zhJb7oac6vrtEy/fPeXULjjb9sb3I4TYkhm96yA9/aeVh8fS8HZ72laU/77p2rWuep7M1
8Y7w6NvKjdIwHjg1w6mmQO6uJ2Sk/4LNO/hDgbzWHuxi8GDA/U6h/46W2tWxsWYTdJsImkq5jb2D
Q5K0y7qdwI99gc9+UBkcyAtN6XD+cJo08jhJJ6WlYUoZSZL8vpc4nVLvDBEWSEKGtue8FxCQ838o
OU1u+ahfSTDfb6pz+LU0t+GdXX5m0ktp6KrPlkimnrU6BR1fWwCsuoAEZkEzlmuCEHTM05Ayusr9
ePSEhyfTqX4ioa9UnLgU2PQj9WkcJlDyKvqtgE8+BojARyeTK4FMN+NlnWWnR+nFpPbZB9+CpaA7
GcW45UKJ2quioTpsY9zJKUTuCPuONR3eH/305/pgvxsCr9tb/b0qrUsOL7HcVGlrG9j7B2itXIwm
cO25vTP7tcxP83emOEn8gT5TkNWwhHsvFFO1Vqlazqwxkkfo9NgCTWcR+D+s7+POOpUUZpDeNfx/
bOk9vsQB+ygI9X4khTHUWJiFpg67jhv3Damn3cWT4+1nVHTBeZ3MUCNRBlPojkv7yMBMRPXrsmBi
Lyu3BjPtOeSsGA0/CbOqA2B2pHFOaKubATWoVXk2InQby+tPshlT5QhgaVkOOpwAvRcl+ff4G8Wx
CZtGpTdVFEfcKbnzgtJ+Y4G/bqaScMagEQMzWxBkPNPgt8sLJ93iUS5bHZeoml98lx3/S4Th/Q7O
i2iJi+pvrfX8y9a8W7cEcL6MvAoMN0FwFrpSQOujN+VJclD6wCGHz4yewG02UoXIGMl1rDLn8UNg
KJaKQUqedf9hCxSASV9b7xtsQUNqKjShfg+tcEjxfxhF88S3iklRvjLlfndOilfnErc6Z+EhJd8q
amlQnmyOeYraBrxzC7AQ/ouBx1lLh0yPiPIX/cB+bmLKDyJhXFRQsbfxGRSiQQPbar+Bz+71kpG9
btBuaZpkcfIvqZ8Dhv4edjhAymigxdHBuWkSbBnGG0n23h6i4U/0rpCNhj4z/+XREPmcVd0qb9Kv
HnSgkVfWnJuFA0Mpb3JdlYszWWK/T525+ROoP/TJz+EQzf44QIsKZjFwEEYadcckzyYeVPWf5FDa
8UAc53IGvleczF+pGevWco9lFtoPJFubHNh4/K6sUEcAkiDFve9YDVVNpv9Ju8LEXJ0tiBL585SQ
/0SibweMGuKL1l+ROFGjCFPfl93RmyxgSxd4A7hcMDsuiNTPg4zaw1Om7uR6mV2hsVzkKQwchSgh
ddeha6tSAUSzpCA/GMGF4X4Ckk9/OMeJemwSvRFZgc3K5dReDg256sek5Ii7wZeggniYkqtKEX3b
eDkdDOoRDfD0lpFqmT34YCSZes2X3rt+HyFsetSAy0WCudtmVmFtxlxrKtdOI7WHMRnlih4A0Apq
IzX3dURoyh4qxBRc8CLyvP8ycIx+MAQNJxMAG1Mdb0Tn4+cuXnmLTRPX4GhaDchUNUX7lLfk95ow
G6IQXvT+jJE9tBG0Tw/8TeeHLm8iPrX56Vr4YN4TjHgV1v0WmVjEFtIK62nOy2H5acKJp+8E1YLl
WMJ1HCOcSAKGi15XFZSbfeNavY/uCB5EPfipEvL15ifCfgk+Z7b17Q+9YinRMeztuwKhXt6EsAio
cey1ycmcJMOckMjJtMCOBkjf/tYzsBc0R6myVHBlEgzGHOIBntNKItKz2tQDg0vIe8A0ZkieFMn5
wLlLExr/Bt1LLUne/21fYh+14qYoBvDZm0pTt3C0Y18sT2x1YZ74qHF+UcHN9YNG2SUdl3sENCYe
aJjp0FZTYs5VrpQP6vYhUMOC4TY14bIPIj2qMg4xENXQhb17pyOYXxVbqF4AdJo+BjP3cYcboU02
PZjxxgBLBJAvWPNWZ2u4HyKRy0uKD4yGg61jD7O5YMs4/hAvvdzEMVLPQF3LOIZvNoiQLHebY64w
CmJDwAXqRyf2tDUdg5tE3LNj0cGwfvvrokUjMw1trr1wi7sifOvvTtfIBksAxKxpl1kS7EmSHIm5
DD/BUvExCmLlAV53NOPybxWhZHR5SasH5j04i3OGucenZAuG3htVOmy39L/ovKU9yXpXUbZhUgzI
0hHLvB0eAv6eJR54BK7fmMTARoM4QJ9dUF6GJZUVfGBzK5Usr1kgChHWn2KI62+R8Efahuo8qd44
FM15xSMz4qY8Fd3gVVYmm8fv2p4lo8hck+0HGR/vC1BbIy/xvsLc6YKygeq3x4yHWza3dO4ztS9k
PPhMnFhqjx4CMBR1a9wwn+eka6cNJc7BTS5vKAgZDu3tRybRrc5uzjlBq4S5LAOh1kbZsq8Wfzza
oX58dSdjeRlgOoRHHDnNz6klGBSaEkb/QQy51lJjgP1blxcl59e9gEuY40pD8O5uXVcMa37oJjcN
awLlxWKcByy2IdUHLCXyeA1snMxkeu5SI3Gst9YUa1qhQRXp9a9Xhif1Q4ZrB1bjlkuzltek081R
+wWGaF66Ut+2oJkIpz8OOvJgGcJwLwVLV3LezA5uNbmO17Xq9QUXzLDpQetOUTtQe1LVoggAvUVY
Oy7jASn3RH9Pb4WA28usKzBD87B9s/wEkCwyjSsWsS0+uXwxtE+Il6WiScfNSg1Jq6+vKHHuCc4R
IuTI2lkspJAAf8u9ysNxlMZcikcPXdw14JGzmz13k5RyF546edm/tSreNpVBRYfibdIEHOIL7smQ
R786DLlM4iLt31dAu3frxXMg77u98Dk0Hy9rfD9jaxwgifuME5Yk0Ca2gh5BYzZD6sVVmRJuDSIP
aycnPwBJVXCOFJh7asayTHi/4C2TjHrHRBqAmkAGaUaZHfywx35FdOHnh6jBRPAUqM0tgEr52iKI
6sUdJeGTQds5i/1BS5AtV5fgfTHJQ/x2mwmhUdZGYpScNc3eqeFpQa2qilcDKTMUPrBNJA65QlkY
88TrRFS2V/fNjU6dtBlIZOem1iI9QlRqHj5Y8Xbs57O9BwYnZblqK/bgyY7zobVXIclnyZ/c3woi
RRHE1Dq+ItcZQPQAmGod/0hnv2LNr/z8W/QLdE6yJYfnDvs71aAdHVDu6shaT/YKfD/TUjCVfTUe
c96Og+vHpEwpXzezwQ3eLaSy+rw3JbBHyZ3halRVUqXnwAu+0H56BcVEcwk5H+aviFKEBnxKA1jT
sjvsSTeET6QOncYdlzhcVbNzJbILdhpttYWT/YkPzC+xgNDxvRHbtgxQ859kiDf6CcFam265ssVQ
02uWOS4qmtoY/LMYwWBqJkjJ4qxQwHfMOcw5ada2Js3s9lqEPxAVEUruvsCDFuZUbs4Fyy8FF3jN
Ig1NsS3OPbb1nsMNTtCsz+n8bqhTlSBQ3i1hbNMCvHbqWcV7doNszfbYWiDglpuTtrGQxGOcQ1ax
7HBeuf/tY7qQlE8eNoFpLvxpiL3ru5w7/cSoZxqpaFC+tvskI2XE9BP6pOvTaTN2t5x6HctFJ+ty
YQwjBwMyJu1cLBMrbzzuAvGH0y1L5fhWOp/wc4uqN2G2MC9wLWVIlUsR52HuEXLO2cLTzly5TytH
ZUCGp4gj2mQBj+3qtKHzdp5UHAYOnJ1K+8e3wrDoC4n+/5l2eQYWIMjy32NrjvrQGAKCumK6q7KV
UPUnVZlayxJxNquUdFZaThMTQKkppjpvVJ7MiXssDNFK8R47TE79xNb4PI54Te3ZlPiekYfIG8dA
VEC1Tz8HXyBcCK7tAM8/VIy3FwYncuHHBsnn08lW1Mc8X5+LzhUTqQybW5ULd7GENSmAUpMhb12g
0ry+apQSX+YMPbXthVYqpj/72VbL3VajlgCuB6j5z5/ILD3CSdXhalSkyF9RMLjFKFpzgQPvmqQr
OpaStHSn2+xZLREI5d6KE0JPptYOTmMIeaYIPJtuhF+8/l4eOQ55hHG2w6agoXekVbnvnc9UYuvQ
a9bslDdq+UGcIKB8mWbjH3zDkDRJhHZfQwFReOCFn3C4QR027VPdMcwvttwKJdlsX14KFCS2BY8X
ifw5tK6u6/3WAZv40xLUvN3lbWpVdeHlJo44JSjSmogo4EqbGZG5jbOiRVJ+ASGoKqYw5uQ3B87r
kRHM+n2lY2lIJqaUfwWiyZ1FZyx/M8rNNjm/Zo8c15nl79MI8kfQiRO9LxRTePAilJEwbdVMivNO
ojRor0tfzVIuMzYYVRqUVvk+sbDJ/eYk1xgbI1nWrBQ9OcxmpnVxBpwKexwrwlW0ae5KAGlpD5Hh
jNpITzVr83jFs+1HTw7NPla/llEe0wfnEbmCzUIIjoyoZYAa/GLbtMTroCP4yXYFxXP7XaHL8DK+
3nZOm3xxjsMvIzRUSlSKg13ESQPGRICsUQ4zi++/p5xdEblztKPBfTvAJQ28k7UodkHQQFSFq51X
+qdnRpRC9Cz9l8kuXtYtONkrF1hC0omoERFfUcKpNTBVKnDdjg+N5Pk4iVRXk7RZpOcM2w4lt2of
vdCRC+a0SCUnTEBuJT4aMHcb6v9GLh5kSZj9RkPp1HICaCvvFxVLHHmGFshv1l8HU7cNue3pnnJq
OicPyZZ7dWNN8HGbZRSrqEVoqqaJUqaQUnn8itMTq8mvC3fRtVvGt19DbbjWL9JWXzft2Uho9dqN
/yRViI8+CAwNU0oOu1C2KzXMlS9vdgHLh+asFjv6momvbpLkmysaHJrHpU5Oup/OHgMeylc1nmZZ
9GRw4ePx9oCgNe53hc1xATUX4UlC/58hikAG57SfqiqX/DECYzemH46SugohMVWP+GorM2v21bNH
/a7peryUIPG2CEclB5rl3KJ6mB3vOP8YvFKT3ZKV8430EQI4M0XQoh3tPxQGyRUmi5FAZO553TC4
9tTa5QRlJRNsaZt65Q0W9b/w34kE6oVXRVlXGx8bq2vuCSL5avvOukPBAEPmh8rcV2KjUeFXG2Su
y2/UkJWKQuXxsfcEkNqZyxHIZHPrNIeiF0ul32/dC1wGiMp/Gt6W8C3DEpOaEU3rwb8uEFkWNaye
woaOYg1JkqBrfQ4mvnet9aqhV4hK42bVjlzEcSD0jMa8inodRRu7o+V5Wbhpci08AAjxVblRuSMC
inggJDeH9bGOE4O2sVlFHD0KxrggC4UFU28x/wB5jM2q94zkdbiDfAH0VBkxl4fxV5W75sL0o/2f
xXIU86KFw2hVpda8vrUewlSsLuv46EGfYeZXOcbYqwblxx8YEUjOaI8bT9oyKo1D9BUmdBCY+yp6
0pO1Fm4LoT3Vv3ALwLVicapFG6LE9yeefYDO9w+hYETmbmb85n79iKK3jswAEbxI5fn+u6xa2/YY
OoBdiR4c+u6ayrOuqj3x4hqsj1ucf/lz/xOi8Mdg1auACR8I82sa5VkjKPLojiPn46LOik9E8nkY
RjSJDV9KKzqpo9EgFPcPWuRZ+HeihVlBBWHgd+A+GgWEBXUSMPv7mDd0JtICkm0yfuSr7WJrMe7q
fBRww/gqWZmzUYL72C89tl/U4Nd2GgAka52ecMiRXNxfVTxJdq3E6q570wHGdXJR0O05lx5nxS9S
lDhyW6OTrIyUnslIgP00XCVQtiJzOFhGAZCKS+mzjfjlrKervBGN44IAgYGSp9ZQoJwuqCsfNh1w
lH2fMyacIwyAqFRPp7PEcESALQgrTG7yLARmudMPVsTwzvCh3u1sR/BJjlUfKswYscSW1uXQnbdR
jSympGCzIjE0U78S0uzm+m78fPnD2/r2iaaHpgctADyqcocmI+H5JymaPEvPJad8X/KkLNIJkD+m
2X5w8+bF0Cv0Pj9aVmvXghxmZQI9WAwOupMXLLDrUEE8H7Fdp++PGil+qdy/Up2Z6OcaV8gq1D+k
K8Mrd4j4DpQWCMYOHpOdDnufVoiPEpZtQ4XbQ9leA8iBnikn2jy60PflvfRt9kfAQYrvxim89pC/
pPd8K2KL3bAEtTJ6yUZOa1Q6YfY+fAZAf12KyW+4XvXiCzfvYBo+KceHG1jOLiOHmIMi+7de7XpO
BKSVLWzqsQVxtjJVgPYKVrO8/vq1tAugbzIrS9BHfIz/hHaTGsvqRK+ug5I+aJahT6c3Mrouuz70
CpZmzKEiqTTbblZzFWbKx5sYTG24lcAzxG6PBknuorX4KecAqQayoDdEBR8yRCZpu5IOstTxW2E5
TmbLY/bp0BIiT8BoDu9hEtCkQ/owb39WAkxwG2S8vMCTZnhu/AhZ4f96z3xeL8rpmtJtLiLIxY5S
o8w+aw7rBktlc6W3ECV+jusRw+U+4nGC9po+wn/ikzeYHHeQkqdBX1UdDtf1sZmbi4W4ekmEskqR
LvKZAQVZYTJiHpfMHNSo4lujzWD7MiJK2FZAmnbKXz3IafXn/479Knla15ez4FpK/dZObgtQ11kf
LYdbyLBrOUT6zVSU016eqiDmt4WR8P55SzZAdJ7/bzVIT2jOOEtwI+OZQtWqyzgbM1dfXzoLxFEN
5odiRbZaVxTxxgRlCDeODIZrATGK2n//kpB280m+aeILVHZDjb7tOb3H8gBEDboI3351aTf637nl
dKgd32Sde3aCvM6KrCxTCDadn30ykbq8oA8Doa8MZRe/fVO8PKMfpiJGzpBC4sJWYjnyLGi7f+vN
7JTNryolpaxoU4qkwRGmLwCtkIWZqXCiZaxbzZ5buTMGLZa2DDhiEistq0+YMCR2zBGCJ96OwHdz
ertgEQ6yj2L2p6u4qhSwuZPTWkz9L7qUbovn4zEm5HZMKJSBNKfxEmu5POFPH3ccORy3MqpHp+zN
fzvR4phvXfftNX4689fMsDZ0PF6dhKdzQ0CtSgRKEYDX6XydKN8AT8tl3URHOmQ1n28JvY5pPWK1
SvIa9n5Ik1Es9dbZeqHqlwJJe0vx5E+XdavB4D2aVk8Ww2wQDo+W8Q5qWWUW1SNDd0Ds6086qXmv
h5tkKnaxSHQm6NQsIqigLSbebQ4B7pO41OUOuiyb4XFsM6xHJk3jf7EsYaX9rmkvLpFjJw7DUPYI
9ii6NDdhcOM8llbhGN7Uc6yWjo6os2mNxxVGjEJin8HAvmCJTKB+AEnHlFh1ZeGET2Jd8jRVP+VF
SGZITJmnA0BnrEBqg7ihefXoFIt2mWvlWQFi8fPKxOynOArxrtjQZiziKhlTyaeyCE3unp4T5Wy4
S+MnwhoZxKVg8H5ob1n8edcrqyk4lLHuztBrMR9L8576iiaORt9UU6AsebrTODC2g4Vl26qE43er
yi8Jp6DIgylq7bdAEU2Vbpup6tX+M1KWSrwOZWMg2+v2gYOnOYLQUMG07pKeScp9d1liVXEuWML0
E/Qr5NACBKlP8x/63QNjYi1tvWvt32gJ+ir1IGUf6C+bzqtFEs7hNT9a/utzccNtAlavPrnUCbax
1G3cr8Mv5jD4KEkXMXyxDE0uVUzM8mr+DPwStlTRoH9JF9ioxfk/3Wr98CUw8hpBviQ9COUDUz53
y2uok3bJ7pyWAugky30xHaBNuCREL8LtBxzzOyqIc8iQj/R9KQJpEchwZgKtIBsThbPADHt3blU2
uoTMDX8x5DTiPVPMN5USd/Qw6Q6UISPVI2VIbEwLe5i5eOePxUPUZniqeDRbTsIkAZQWWSC927lw
ePrPPmvvWokhs8dFddJ40kAn3geVkciGRGlUCEmaVmZFxIPZl+2Wp4bbPxDUJmJaGDdgjF3ACnV4
b1t4N0Gx2RbV/+edFcSy7ou3fAd8nZsF9/KBoVqDr82GJ1gR0G1VQgPO54iDa1gOorh7paPePkho
fFDcm98DN0LcjR9KENvs2dRwU0W7hO6scjEULAfR1DReXkIKCQXmmgtY8xzVnww+6fq4dsMnGjOg
hlhrJlwLqaRTq1/x5BeDhM2nlkPTyb4FfLtC78ih9h0L4R5OFHh5SIScJesnRAvncWf4hVjcFAgk
GotAmNhQQYAMD/sH0DZmv52lXIY+LYOz3KBZXaWBr9EnSNP/z8VsZC7oink5bbGvqJc8zTILVZZ5
X4d73Eg40+d6Rmtlfp4j6IwBgcyT3vaX2qH0/Qb2+TJLOrfsR0mB2TaRGyMKkh1NE547YyeLq1AD
X9BhrgslBSKQxNsRwgSbipoWbzj4r5HKVxdPNNeHAVe2uixzfA5ya73L5PH3F8Wu1tQ8llFlTocJ
F72cRWOz9HD3y3ViDb6f8MQ6ZHnRNWw5QyTlksdjJjws4LQIQbr8RcRQpIwbzkFNfu1Gn+cDRbdO
P0lcY5U2gHdoJw9a//J37mcFLO1Dc0w9L1NIpXjCFLXONZrOacqIiVV5dC63z6/Hj6AIvcNAUyBa
84XULtU6cIefU4T6KZm2PqBzbgdKnLipZGQSn/4g0omXm7pThEPE2FxYBi3sHCX8a4D9YPBVdP+I
dVSSGC2KA2A+1mQXzLxyWsmuPS2L7LBTLfyxAABt+JZM3nxc0jpYbbO3vZVVbMFw8eGFx8JdS4G6
OXrJBWOeIxUMsVoHeWLDnS0XBkZEge3GXvPI4mHJc9xl2kIef4xsaJMEw01nO5QaeljqB4dv0uT1
AUaRIgh4GSPdTkuT/DResl8Qj4WGMbfhOn3U+mSW+dS5lvBScn0SnUHP5OEkD8QFbDWWt7KJkq0U
YQlKrYZCMZI0dfxNvv7Yg6UzySl5UiPRwfhej4BtDISmsfNPbwSVWcb3RZt8MJG1aS542ZhzuZt2
FjWXCodW9aS9c8K55tY9iTyVpiecLcE+AjlHk+eimzH7nnITKtQv1JUXqW9BVePdkNDXPvWahdNV
N1BlRlGmVoiP6nl4LWz1S5K2uTr4uzCKjpUseYfuNCM5Mxrxl5j87npsS9FCPmFBwdNHWifTVwKB
dJ4JOiSWbqmIXggrNTpzqYlQN4oGeCcNGrNfFUn9Pj4zZeCLokCx8RUfFgHtgTrbz3f84XpPKTsQ
yaG2eth8/F8zg/0jd5m0hGHGQTf74P2jI0W26Yxzqzjg1kSYobLy6TgBl/NWVKQSYvmfLR1Q2v6X
CzeQMyeyq8Zwprq0VFXdGLnEcyFPWiTpzuUNBhB3OQxm/66BwO01Mutf37QTTz47NiH+PBK062og
QwAMJMSdLa+N4ImgND3G6s2zQzng0va5eu1U7Va6vZZt3jfQMcy9M0+3zKWM40z8fZrRQnbcMarK
PLfWKOAm0WmzsmDVyqqIh5+H0uU2BvrVkT/Ag/SneU6TxOJoKCPWoN3i5XEAlOU7G3MkkZltn3Cj
xsUvqsnmhoSg+Lc93pljicnxj4IG2pX7o7WTlhotc6XNbKZoQBOzXRPoNPqThIdCtSVXw5GSrFZZ
h+gYq6ek55kMpnk7o39Yz0Abw/eRbeg0t6NC0OVMdrJLqcwdNd2Wp60FyLAHozMG+Fwxwnt6a92i
BSB+qjDWGo0WubEXOEA0wmZq2fCgo3QdEsV53Z6hHqWY0JNSpdk70vYl7a+qb5RUv2/hQfXvKUTp
Fhf99+QqTS8j2ycmDAyyXwIax1Cm5vRnzm8un7NEdDyw+WI1xqUwXn5iO5abqhMprE4cbrx6Xofj
c8ZuycT16D9FO6vTV5c+vB5XIQ9sBxg1jyAfVkCDIBTLvkTbpgng2X/2rxH0DvF2NIY0Wdct67x1
zbhVWkNfCXoTmIJu030vJrIplbxUIfQXyXi5YLc5va6hNL7CWJoTUUUK/5FeZwTR3vQBfnP24u/M
44Mahk4nkOVkVRXLtnl7FC7GUO5ALwyykqhUX5gSIOZnsfI7kWeJQyQ/55QqINx8EkOIlz8whZn3
bUGcGt0xBRWqBkeHz2AEZyHNlPfHKM/Q85GhlNnVaSzJ45vK0yTxAnJQZfnb8qofyj5CP6aygBWI
yICkPa93TvTZtOb2PJrCPpQnCO/E0Oc7XeMXvP2LU3o0drqLOJZQwopHYYAhoJ5vlmxDrrmuxcmG
kxmKsnc4OttPKA+3zJtXajdx5fclSNjDq8lg6sx2R6Ntvk2gxfG++TaEIEVNPkyxXFh5b+8wtH4l
d1P+++F+eDPmvRCVmaLaN0DygdkKI+ljZsryqox0K6MYWrWNiuiwbIL384HEcxpwPuLAbcEcxNBx
odSG63xi2rZvTpoJtaVy2VoLMdJ8oXUYmgRWi+Ku/qaadou+BLLlISfzgLHvwivquUSeW2XLtDgT
WWXeXNN77g2LSPiUALuuarlc/maknavmtsNzwLVxaFGkXC7lDqbTkdVSL1h9PAAqPDhuyVW13zA6
oPaRxvjnPdoxLLQy/tWcEzLVZQLx3+k6gWya2/0lk0KTI8QtiJ66xKgdTId9WwbCoj4vakqmoanE
n8RvlO4B8qcUGaOcTbCbZoR06XgJh1JqHtGQmdKFwJO/zlM/lzEh2TyYCf3Udvy9RvbGYHTlyd+H
egvZlTX0CmYsMhJaGmqDhMsajcw7oZSGPPRklqAD93cqARu6cLloHSG+XlRCWtavJH80mWv/j29d
35oOUcXjBRytJXsjXchNM0WPQto5QrSo2kVfxDOtArIEegtildQN/l6XFNfPtnxSOF0u8FKbOXI+
9JL310StL4TxABE8GOOLxGrnSk9i8oKAEgbfEYeCzQJjWhNcUiUJ4mNfEvcgRYYQF4281BHbdxNe
VDI9+CUU03YoDTbKYHMNsb1rbJ1zB4/mj7gzWZaVZe7F9Y/ztRxaSAv/kiJeBCHEA+3CnSqO3ZZj
/6T494aD1CSUs8fjW3YAqJ1RAw2tuX50DUMntA8Et8zg6KhMOvWVmwvKHHWC841PdWS0cjTvxjbx
VFA1FvtvLfgJMbKKdjQuXBbJAmRyq33yYf92pnXkatVvPRBmtAG5pHtvThN0pXx9UKP3S+qoT7dV
cpxALeA+pqoltwIswDWeMgjKfGTPIxJOwRRUikYzPQmDZsQ/61AAdeiys9LifCs0oWON8dY7zzOJ
FtaW/pXQWG3/pWCgDN13PvvHE/9IkQtA40Xw+TEw47fK3enOCms+ohCeR/hJVryXFiEuVo4CqQEO
Y+CZBeCd4mPQbKoKmaVhZSiCbsQoMNoNntJNll9tA5Xg5MNObcGDfNQ38DW09DBKNMxJqjvvtK7x
bmRN9c1UW9iQ5hrhAIBjp02hTW9zQIMzZAcFJTzL9rLaBoEkHzq60k6D5M85T0LUEfJzHn7460jl
T+2/mHpHSlMYZcMe4GdzSvfMno8YU928sJ0OC2WyyuQrFgpK3GPo0LPA/dWz7PozIdk3BECTRMqm
tqTPPcmSBX64M+O7FWzp/2Pqj7uxXNIz82pR4mFyfnk/Hv9kG+sEt+4xtQTts82fUCNUMMYDWtw6
N+ZTIJ8DzjskhvPuSkxxG4wH7few1V0inhWXpu1d4N6GuVXnPkjwPKjxdQBsTcM5QNxGotwmveZU
3O0zp/nZdnjCBHHC5KnUEI532zS9268LC9RUbGYPFhsqWmm1KLHMve7QKYq5qLsQS9sLPzJoY0oQ
zqusej8mOuI6AwzDFAxE7OlOiXKeOmmstmbOWDed0uqvAsy/8yFijbh8fjtOGCzVQ1zIQgZMKUFt
qnlP/CY03/dBW2porBVLQ7k1Pmk9VW8Xj8TxWiJfjRfScxClGpmCmcd2ElJYKo8BaOLg3xt0pXOQ
Yd7pnhbQy+904JOFwIztEi8/MSOS7qxBx4ZsbiojuuOFOCbxHqHk/zONoB3WwATWOXWjUjT1ttWK
fBR5Yd430BDMnaFmILn3IU5o9LxXxo5aQsv9ROBQnAmLQCTUNyvcGiQB8MpeebNpaygJjfDsm3e1
CbhxGz97LhyN04Lr4ChD2W/WM/BzpTp8k7LWskJUssADz3Q/QYawx234dBvHKV8nODFUtHJNKYIi
fyG5rfVGG1wkWiaJnTsmtkaWrjDA+PxPHT/H5x3CNg4ryooRWCT3hnWAj8tT+ftGxD1aDbUsohbI
qyjuK+fuXZWE6OiBsKT10Hk+drr1e60K6poly1omCC3EGJcLB57wO0eIyfjzZKkVpNimD0fIYyS6
cLcPSnoJ04YkUJ/JGa/pRi22o2ViAYwxNE+y9TaWBZ964LdznByQEVj8dQckjlbwuzQw0XA4EV8H
sMOFKAf9sH06Z3j3ng18ytcBc2LhGSmg+1SETX/cul5YqrIkXozOkoA+WvTYZhqxf320GRAQNpuP
t9YgSNHsseyiiaCZ8XvmC7nsYPw+4rt8NLiBdoNKceQv4QDQMWwEFZjSqxdQ/LIdGpyCszfM0UxK
zy40cEMS4v081J/eWitd1P5ESvIqxlDMfynSRpVaauraDemCAMQA0/dFxK8yY8o/qWziHCtRxFEO
3eLSYuQOwMEbJV75YVnu7+C5Dkj5CKp6Md+uoAnpNGdwWda+V1fc2bPbbbAOPTsudtpGMpYlCxkv
hf5oWvdK52QEKabZJoyNmeXDWBD1nKcUbHFdZ38DKjJ/XDLia6OFrifm7v8My3n2Z4QYM52ekPOU
EUPSbEvPls4F38tV1Nn0rVBh6zvsykDvx6oc0HTmnZcbL1ON5uBeOVk6NA6rKM0y5hjcbHx5gmH/
YDNB3d6Pp4UDdaUZdTgQKWIJ58ZVBQPEeDXEkfdVcI0fswDTWZYK3aYOT3jua/9tYhOm3f3lZu4L
sXPHBTNKYvmYqC/+WsCAZDyv0sAtgVkC1Vy6lb2XP5vgYy+nNfFHAFHKQMTvw3ri+mUQHYiq30KE
ptODNK7RRNq/3U+X+PfGHOCWEj6/3ahdaB/4cXusBn8lny7FVO8Lz3Jo9WZIX6bGOD3emmxPyQR/
blHPrnMLCOCdYoXLXF9gEZIj+CAO2ye95PbU3Xbi33rnzOmOQQvgQ6KitiWcfvOACr+sd5EjP0WY
NhtJeEcuguWNMKNDjaph+cZabtn/Sp6h2eMOveAvlv69320IyHNhNvDVn8ntV1upaTs+lTHPzE+U
hEyE+KVr5Kvpn71mcrrDOd/aMB2E7lVpUXLwPSb6h5Dz3yq1wGyC4SOj020yNn2GGdpOEVdimf88
UM/3ucXwb9fpBVIbxorWCr2fEMMaPVe4aWwFCsVVV3+Y+WxAH/6C6YZc47gBMMOs5z5Y8gDm4fxJ
7CkOdIyHMRuM2HEpFolPkzfJ+MHqYA/Vauz3REpaxsr1jRMN7xB7MPhQK0jjdW7bG63ydhWzQo1T
dAxdj7e5LjCeUaZ/vbi+QhR7EaQExQjzvd1Tsu3x4+isd5h1G+Cux+DrE//8/XN7N/+Jo8kbHoZI
ryQbFnjunicBALAlP1sPVJrT2fyoUMN4p1x8Tly6MEgIC3IV/IHUG/BlerQ/PipQB+w1YLnVHyLj
XOPL8pT+NvZOS70130/NB8xJYovgOG4jQKWYw9liQHVrG5rHSFNmZlFKEdcAMjkIrjnJDOjml6PH
iSivfY8EvWfJn8Wbb2SP+5w107dgsT35OmQU+Rl9Nq+cEKODGIfkjFDhdHz5Fg5KkRO4BMZqwTMB
ebHTki34HgGoL7mipCvOG75dwLqIEds6QjDM7U+zdUp0y7nUWlqbfD/XQyRhwxMNBP+NqG5SX6BB
DF1TmTjNuLu51Kv2mcwlRU80n1nQF3B7vqKmnkFHeX0RuN/G1WKyWu2fy2+BokXH2MS7jRAfm4An
ZzBgPxzsu3jQfbhvZ9EMydZTC84NeDSckrzwHqqzMuuIkE9yMxCtoUUWxQMCO1jf0Bqmi34W70ZF
J0/cS7JcNo16PY8kZM80e+T9M+a/xtt9e9t/sAn8mzsQkyf6cmucr6JtmiGDKtRLvXQ7qI3TwAdL
LmV3doPSvS7loWZhKlss6FLqQxej0nPSc9XR+TEB4hP/MnoLav3eNBqSquPDAu+pw/V2Fp4JonwC
esCILqz62YgftrVTvaSWEhZ0KCV7G+JDQIxexST2BQsIwfBTdpAjpe+AzPFtq0DdU01Wy7Mt1MXr
YPRIgn2v4zOu+Nw+OdV9VvKmmmiFvEjZR/Op6GyXc9LZdm6n9XWHoUlVys4rn5oOGMpQm1V4lYxv
u/Hw1tE7PwqvE9RpuFnn6gLp3iJP1rEwoaQQ2SLO0bsXNe9xXEZaGWMi/70iwbLWKQHDMPB0b/hH
x4jx7UTxEkd6lK3QObow36GhmG5Ygsr82viKsCBObU9Qt4fN97+KlxB3th/0yjkh+TJHJxZrYkYn
QBAvftXRbZPp8+Zqyoz7dTYAkTDvMO4sBqrYDI493S1SQ7EqXZfoX+utV8NY4uzTVoFs4VOi4UJD
h//iG9mw8/TVVQXk/GqdL6GDby85/umVzajzuXn+BaWC4JV6JA7KI2qQwLL1uCL585kvEyOCeGPl
vvHUwypMtYdPIGqscTZ9RsxfgGimggU1bhNaViV348WI6obTipIMB/PApfjgLSeYr05NO5+U0rcC
AIsjW+iALWHzm6qp/SD6XRYKICTIO+cooWPAuUsDPmzpOGRvyhq4mL+TKMWfFqFLCuI+PNTrSEbH
ph1qhtQt28MSdfL8xmOpJqbcTKdiyxLJQzU4cuEfuej4F2PgMUhb/4FmA/f9v/jnsR7DLWaQR+s/
YG3xfgnRlyHtNhvArzsKcgB4aSVjIji6BakLZRdD2zV9sZUCnwjtHOmamTcayZymFHp07PtAaVSD
/AuK4uD4/8FT2RcoaBqWCSXuy5X1PVXsQKA1UexzoKKt9AhkE2oeni+DKXxqArpTzlmCdgBInDMA
6dzFpg7XmuMxdNFBzt1OuPhsAmYkT7sSw3YZtv/eO7yay/uJ8wEkxJ3nNaqaaqXSjWKNiHMawkY3
52u5R3oX8grsHTuCb/5isc8vtcYRbgAthheywjBd0isnqIiHx+1INgAwUhOgpF3QfM0xVw1BSNGD
xwW3TBtccYPqgSZJG6qclgfjfd74bOdSTy1UJCuc82jgk4y1/pJiZW1KHRbrzNgr1+ghv6qIfx0n
lz6OgwjcTJz5JXfN9DAYz9RCtgZdNRNxqradcDMBu82ut6w0pCj4CjUdZ/uN1abIAa/y4mJLDHzY
9xzrf2RyjwDclexiBXptNdNeO62xRHZEBjKWKpMG12+b+7sb3Jp487TnB84hgouzxQEzW2EPHQ7j
6StouuVMir/1LyQVrGi4j702xXAlo5wV7PMy/ye00idjmznqUY8Ty+eHuIoxGKRGVb/K6mU0VdFy
HTZRNomFlZbGblVXowSz2QQLBFbNZCAaaRiXC1cTkPKM5sV73In9D76ZWAsDtgQJ9i7j/35oI7KQ
oC68geclNzCfup2DXJ3MeP0gxsMIlAU4MzQmWddiPqSmYnHJ2wSH2oAwopSz6gLs5GOoKqeEGZe8
pVVCXUOjt1UCAP9a9Fi1BfMw7NsFQ32G3gMRFHd/6YDVFk4d9e1EOzx+++fjU+ASfnfa4YMFi3r8
dEqugbdvwEOLexKn+d9hwkR4BTGrtdlsXO6amcvKraGYScgq2/XWen/N+7JgAVpkRptcgJ2XYhCl
E9VUR59EPGNrYt0VPrrJj+mS++I8ZSiop9RauGEjzWQxm3BcYSfrtjiw1m0MTwrSLPmw+SQVqPE0
XdnnTuCvII9M60iVqznJKFc3TXU2wxTOABpIAitj4BTYW0RNxTjXAF450qyZbvu4+ShcGbGCu0q1
6hDwGCpeQU2R9RFUTL87FEgS4W2c9mnDWklLax54BNP4WaZb+5OIDfGuluD07eLjrhU7YKGe1Cfy
HQH9LYI0dYVoH4/P1aO93CbNKMZ3mgUgdg04DvKquk8VH/Mgi0MRGYbJuYeVc5I2JaYugDpTW3oL
1lfO7tDiGZSZsOcLSO2PtugZQRYjRHuEIrUA8wCGx6ePQ4+HTgatRCp1B4HsONKxu8ZtQGbSGl1/
xPLBiV6FYhzdpvDqxhcIr+6+ONI3hSWezNQ+2njxJfntxJOtDbhs+k4cmRQmoOTlYd2nXP4tV1dR
4mOW/NVn92NxX7ghh5Ojw/G6QzUtcxUrUaEle5W343LBY5Jhh8f5ELWhOEhsF20dFvpJ4B3VJnPn
eLmKF5RzWxnh2MYPRWpa09VzqeEZw2+7j2K67gdLuwRXVfJNCQ6sncvsp3rWGCCizFuPuMTlgbWd
Zms/BGyqXclMnzdA7qjuZ2LqPpm8ZOvSgKSLOMuscPjiVxS90u8MMJMVdGjMuWcK0ymibtekh2Qp
BUBP47olC0zldWqD+9GtRZMqZG9LT0v5YFHYq5PZLPtoMDB4nNKtwGLIx0IxursWbzq+VTYeKMly
L+qw3gkeZjNRkPsCGcAqUiap33sKAzL1Rwi/Z77dAp5AUAD2vC9Og0L3enQTrHmEPgbKVWTuOdpv
uQ9CoJ/3f2xGHmxjGUzd7GD381jRZb1t7n+6izsqerE1lqv9gNCCjUgtF+24+lkW5I4VjkJDwnpM
XN8xLdleawxEERBCWzIV5KAxqZanPaOXqChysxhpdG16ZyOQ1X+R8fLARqXGSz4DR6pMseLI0wYF
PeKzGJqMG3kxSn8koBPMbaFg4q5ZOc0bge2hWnQq9mGOVz8Rp5qBHUv2QeHXIvdCxZEyUrlh4VEe
rMTt1/BgoUqlseDbaefURDnKodwAEWEDGhST5z1ngyBPFVgj1UpprpqioDA5nrJO87wnTj8eDmU6
zQAbXzJ7auYwgZ6thckDYxv2ta5Msj3K7nSIzARdhzBZfERG+i93lOifjqEHdDF0a1UESTM36BEH
E2TdVegOq0vRo+KViRWSFAQJSM2x/ghLUEZiT/5/3uCUKLSmOMqZ6/Z/MiWWPxM6jDkgi3ePfSPI
TxoKIcD/g5J2N+dY1N4BPpftJ0Z2cWpzeu3g8n9KnFcbcw6cN5siSKIPBS6w6YRsbsIXFEimOo1o
9JJHBRpctI++HiWwQv2AKG0drzu/2vC83nIfyhMpBfgAwc1W5KNFPr+dYW6Pyis7GoiCPQs98TB4
HfAdy3Gc+u/3pWQHyflb8C+YjoSW/33kz7zfGLflE1XQn11ft9+F903eeV7C+MGJ1JMmSbZdTdHk
5KyuTQWBT3aBJk7kglZkoqimjIcHFQgoSVQiHIIxxVE5wzxVdO1urKnAPTwCPAN6qJlkBL40u5kH
xMemeddgNMn0WnTCQC2JPBoXEy0u9jON48d8UFYhWNNyvBEGmF63I5/aAXl3nwSxmrG/Qu/wqloD
VQOZoAsQqYujCb4+0YIJneQf0kRT4SytSn+TX7yvSPAsItvbC8HG2LKxpWsqijCws4nCvo9f5uJU
ZdRugcdxqm4DGCiq6aF8+10B3oGsGka0QMf7pYMHKPnPkUy+O2ll1UURnMKd+ZaAFUhS90yLTUQk
tNOM8XuQh+KGTIXuSS8YN6BED+fBVQ00Y9ZgZrZRhoUclhnZtLzR7N0K/wdM0sr8oBysJ+KTUFKT
bztvYhDsQ3cF9dV0Cd207IMcshAbSR/6oo4O832v32Il2pkzUmJdcj4Dt83YVGAjasxf2puP54Qh
nXrqnZV7mxU99hcuhtuDAzNKTT+d+2Ec4z7r8P33NWWNV8SDPd8RNi8f7JIHSHHwwSxrmyA504Lr
BSucETz0Mosa6VCD4rX0KSC3xAJQsbKuP2f6rTQcxULkZx9uVpReOqF/BQJ0EdrK+ugZwXqrgoDN
EW6QxwsMXuGYz72bZ3QjQGNdCBImH55YO2w3G3u6J6/5twImLUaHvf0E+J5PvaFJL8mL6EaF/Vai
Op8ahDY4yXjnpNBy8wXW0fdmXQS00P/JRrifJtoglxjxqzoX/4hLON1NvuWLfrbuPhqpdwAGEshF
/Nc2lrsaxnLp4jWKkGXjyjcCr9/pi4cggJoplL4EiIu45wkE1AMEBcLRCNp9NmnsyajJguipABqJ
zZ5jJfpA+GTXtrVCf54+RngHuiFHE+lSC45NSSoe4/l1WpSdPfDk083E5/DJ6vfUkgo07yxWS1qt
sTv3FSH2KTnrDwlXtJ5UmdySfhgQNorU2maUNJComYi2LwEo+qKAk6HXiTqV0QZMsL4JuNw6Bm9X
TDHsvC6IyIL7I54QXn6p2xPbuUAo7yKZ8OOCQd6uCvQCuVPSbIuDuEE/rNrAJGnG/GbB4hX7oeDM
3SwTJcK8YXjsVSlvKJwIkjixHLW+TbIQpZbe0WUyJWkZgnSVyyrnd5G6Uw1gNWU7l9Zb0R8ouEic
2VJ2o9R7uCKjl9k3ePyVzm24pnM4I69mEGHJ/J89PfGCjwC+k5T4/RvI6H36Yxav0jt72WpZiMX8
EZ0PISIfMB9RHGoNibSTxUGW1nU+67gDn9LIVMlNXwk8EfrSvWGmNHD40qqOLrjsJ/zOOSXr40Zh
ov8i3tiYDvydeRoAqPXVzxGgCx7pq29NDaxmJ5vRxxHzMbQPyCd/g5UrT6enGuV9GKp2dlvUzTTq
wLBhUANbzyG/Ohtgid5clxvVQiO4df9EDfUQA6xewmDIyEA7s7TKQTJkRJju401CuzmVaHAM8tNM
meCRlZzObi+O+CHezS6PcA6xVLEzb3s5O+YRX2ifq4fnGHQ/wNzl+Eq57d6LNFv//BoAWUrn8xqr
edYX744zsWQUmuyNDi5R7CHiCtbjip/KWAtzoW2P6nVlpwhm1VEC3kK/Zy5HGyArhbidZA2cve57
ndGBqK+9Z0F6JcLvGl46tvKpvPCmUEIW7oluryUhct11r2VC+kqKlo5z7RyW3HvQFigpFH0yq7KB
+aFY4RfpymKE6/U2ZGlf6gE/O4CRKV4eXhc8HSrW1V5u6AjFhd5HhEDkxFaiKBykFZdbSQW9pvGb
8/wbhiP2cv6rb04DWh/XVDY6gHxzJPxbGxfNEe7I20eIWxwMojgJKyMrR660iO0xJcqGXN7+FEOI
+/YdFkFn++aG9Y362y1PPLzik9vRAN1i4mnvX7ixpdAyj2oU7qb0Du5ihyF1ne0LisdE37WHVNcW
rgtYpyCBOtbR/LeUgypwK4978XO9zZ0+ACMQZK83csXiMyDVbx1za6IcAJKk2suOhyuF/KKVayrA
KP4Y9PSTUmEazI7RvsEskp9iHrFOs0chiMZXD3oZZ3Y2Datj7QTo2qiUeTZ0BvyEIrfAirVyjfMD
WrX1Lwx4MkfMdx+TQgNSPuGaFRv4vyErtL4k6BdctA60104Bxhe4PiwHvXGybkLyHvL7emolQMwk
Kjr4G3pJ77+h5m/cKcqkNhNdXZqVuIvW2qWcZmsbHzhKZ7eL7tIZded8bdS5v8IUEfLRNve/pmil
CHUTgNjD4JWv6aUfC+DQEt1mkbGtSMY2y66gcj/OG3CxMAELw3rZ/sELBDW8NqDVJ+2aBjgrGAvu
DBBOwLBA1bwGVLLgs+C+QN8zmq9LFngDux7SyvYRJlNlOIdV6g2QXKY1LbEd277ceqCSEpWobVUn
XsWAvpVS31clJILpLvpci031CGELYg5Nd26FVZY5dn2AMPEOBai37fA0jbArnL3ROLoLWRGM+R1F
JeORz4Gt+Li85eQYxTK/8kVpxlLmZ47nzg9/9E/yWl2+9yjIHH35+N/PM6vuCF1ad9LB8sJ5PUps
DjQJV6nA16jGmGFLBu4Ul8wSEgFTMfyhBh9DSWz18hwzeb5mTmfLOMpDL1yvA7tV9zvDlQ1d+i4F
NyraR7hH0l7c4gFomWDQKhG00tUjX18gk0cOHp6j91iXv8sl87dvwZpP/Wv/HG/xWcm69ZfraXWg
ErYvbsV0MSE22ugix2mLNboYvzLFc2ng20TYGJL0Yk5GZXIc1lU3x0jJE/tqeubtr7krhl2zIPFW
v0dpNlyNe8gKVye/Kg8xhWEBQLtUc7tEsC/2s4nSoGFeA4Zhgm1znh6MLFaEvVbwsYhXcUPlcdTk
xOd3R/9ptGwdajwEzvQzyZpTNpdsghAdx51nYfA5MRGNK/m6dNQek61ZnVH6OUCvTdg+H0s81QpX
zJEkO5nfOwZb4bLK8eD7y61h51NJdLLa2wM3S6xTeeFoQHU1FdtTduRfoVFlNe+YXb4TQPwtC8N3
tJeBKayQzYBD1tuvnQ7fl0XJBgTAWt3VF9WQE2I1T09UKk2tkfin4VSYosJojdrs9p8ZkwTJT+yr
JOsntelCtAeaTbs035ANdFRqQs4UQ3RwHHEuvZY/2lND4fJZ6yz9QI3GvJ6jNYuAKtGqoKUOj89V
vIUWAbyRKC3gFg25rS6FLP2uYGYY7WlLbhlfpe9KkpsHabl9DbbzGlFXinCZVb7AR6qrmYDCqPy4
g4OFhMEI2UkoUaBDXPu0Je1xnqiPX1BuG22tVz+E3oTXlyLRQ9wHRDUv7wZ5FJzadXADU2phtt0O
RTiWV8yqXnO4fkvjS3C9uV+r1yAKyaybDdn+O1Ffu1btnFSVfYELlEFSIinpOyqKdte9AIg6qiiI
/XsZveLTX1KTR0BM1HYb4Hcnm9eQwkbm7iiHUuD8SsAomCpW2ny5zSH+dgB3dE8PEjZINS2jAJGC
oWCTb3v5YlmF1uLJOm0212H3LauD/EZ0E+s5WT3PoGEtpZ5rXfViqJdQ4Dh36omzL27JMASpOjwr
iHZyCPcCFHaHDctyMnRctze+X6i3vMLi3J3jz09JgFmFjwnnBpRQzJRUtbRzIOSXKvYHX7mfbTUn
0CgrGAoHRWGg/Jm0P0XlqJTKiEAyt7f8eJkDOIK+n7cS38LXP4MElApIMdkumZZ58C9Q6PBACaFf
w/bNjJciKq19hv0Ab0IPa2LKg2T68R9KaN1fX+iK2ESbJmv5WAVa5xoBe/hxHP4FWGHrY07MLFW2
N2FIof/Hbw+g5cNxeJymHIKMaQc7TH6yLBNT9xgooSdCVhh5nWV1i0E1hIz8Z+ZbuG6rIS+Q0bn9
cAczeJZd2U/S02EFVaz+sZPUrpmfWxg9gro7JUSSt1to0LnqjHMfDx5QhrR128mF2hsPd4t6C9SP
O7/LjKJrlA4qSRZDVOu6ECr8CgUoo185Dwe/Pc3bP52m4heOQUMPo7NUHpcEUfPiChNkvF7jsEH1
vCQ1DscN/02LcWk+H6FaPPz1JQV8kUpaGxcDAMp/vRurgytNUXUZxufXZvqYlBAr2Bqw1LmVEbpe
0nZUtcvRsfTJlIJKKxxRYl1kZriqxqM6ondWl/qbRwtX2lRXSmVFfVvkG5cnkCSXHwu1DdI8VDoN
lrf9stNp2ieDoUqBgzLM2T+JZXjXqhOsJDniGHNkk9ukX116JDKrt0IbWCC0T86ZBIXGP1QZ3YEo
f2O3Tox2YZuVIbqsIRicBEgAJwdWXhvtJIdkQVHUflsVQ391DyJrdm8BFMEhRB1W2kl1o9eY6YXI
G9L1WtriyCE3+AMqNcSnbHe7eozaDyNH0s/8IfeUqGZj0El9gG/6NorCqGROz2K1xWm6pmekEnGP
A7ZYRW9WBUXnZrL/mwBmDRv5qNBO63sG1Bu1Zhabrie+5BHxtUIM/NptG8BImYMyLEBnmNXS7+MS
C2j9UH25Mu/BpaonYW6X30v2gnSbqjSIr3GtW3Zl/TJFhoeR+swmhU/6qW1/v0w1ojn8aVcXdy2L
w+0g2aFToPzlMHoeVAUL2lM0aatp8iNUkVDnAA21/fYI0dzOT7GekMQOHNhzZo4aMIlwczE/g3Km
sGn+JJPVP6mwVDdzkaAI+X9tloSn4ejPVq3OijVMPJskLZ/cwP4U/XSSjUr62mZSOm9SHNU/hD0E
v+FFxzY9nCt9hTq6x6T3saXaRSsykhkfliZjQdZyBhHu6BNKL+p18PTYeUKvOpfFgAZ2TezwOxWV
LVAkVuVWoEa3cju6z+fpw3XCnMI05hfreF1HS3R8nw6QJOIeI2Nx3MhgDkHhIHS2sSHzoOXnVSDe
sQeVYPPEUiM2wX76HjXTF0AXYPZ7Xtfdgg+9wpG+qruF0bUDmnuLfMKvnFCle0kOkZ3J2LxRQ9yu
EDy6E/GXE2IHa4xa26E2ikWsovdr24jXXF5N+xvQhvuPNszJBO/Hgg3Uq/nMwMJA86jnMskqfAsp
cYWVVGE0hd8w1HzThHx78eCYmo+otL84PhwMEbAaKJa4ZZ8cItled/FlN0BNScea1C779ogzMX3S
DPof98UJUncG4WFaDX5INTqmJcvXK+pJGd9YW3TvlDOKFIVF73vqWCgIx0J+xK+ch8UAarUuJiH4
8yS5jTFSqcffA8+wzDHsFmvA7FNzs1mx5fxKhqc5QxnG68xcyGwBecNe9y5RFElt7DU8WJyoZ8qS
alMDZQ1jV6gPCctrUpEhd6YZMvSLhUeZ/BB3hR7jCGqkl/GBmimDF+7kZSApFwG4iWj9OeDBFDge
X5le5L8kIV2e58Ugb9zgk/VxTdqTFJBQBGsfVzoO322wkfeuJERI8kL7ETcDFSj7kQkRdcw2Xnwt
GDBzSL6MKkrnRCE7oY13qIp7GPG6EbKpQPnBboSKLa62QEYKwZHtPdrYBKQb7nOGHskUUZyLW7ID
au278Kz9bmRYv7RhfqBXzGjQ2MJb4cn7Vc+6jMA7CmQACOklJX7utRPBefx5xYyAj2QooAtjkuJS
2s8l0+ndj7SKEoP5Ox/B7oZ9XLjsTFWgGDeVo/mEmuX45FizB7+74tFxRN1dMmHh0TJaMgcmTpiO
njnMH79exsTN9WqiG3Ch7/tUS5YuVjeFLIMVXtnaT4pH3eqGjqhdg3WKKiJ68rdMYBt8Yl/lSGmK
ZQB078Hw/LoisxiMLTIPAQCcCXnUgC2M32vBmzJphMzB+FwF32LiQh7/lhkniKgxDVHBys6nW3n3
K3AthRCFcDRqHnqBK/vQhWYQlLXxnrz55Bm0XR1QKsanaMnTTKTrlE4xfx19A2Z3uP+bMTQJTDbg
xktuGAV9SlIkmsYoTSZf8HLNE6cCkob48IjoyIq2/AHck1yqAI+yWXFr+H0RsIK8BrZW5gFA+Fwm
CBwlS1uNoCrTEwRW9BQpC2eQdcIRixjWnUwhcU9OfhY2sEkVyKSz69e/adzpp3BCEcjWiK2sMdBu
luyIiEyDsgISxOpmAAvKAkmcL4WI9DnyA/b8EZi1gOWM9WKRZDMcfZDhBjnoRQmRo97v/SxbQgCx
QSlRLH5MqKji4S9gOMZLVGGgOFoqoNVpAIX9+HRcKsju1lMyv3qDtZ3uQmNH0OVK4VfShp6k+wqE
c8c4OuTztHEKPBleEo3Xc8J/Pd7D7HnaEWP/LEQ2JZpeXfWpvSLDY3hXQvxHXsxfeHq1JOgCF4QQ
Jn/aKdRU1zbDO+AJ/+5VuMHCQB8zF1tFGCCWj81COdEWOeUm4FgNMhH2ODjvVuAbTOnaSXk34Jne
JRNNWNlQJezg5gCGzZ+zxmJUtSuWFUCabsg6djEGNkeK6IHAwETdjG2AQ6e7eWB2gkY3z5etSLJE
iz1Fx0HUrPvIH3n52Vj7jHBhNiEL6ZRcAA0qMMUqg9ZnW99N7wS35gwWHgdSnwKK6p1flFmTx4K0
UhE6Q5/Ee/w6egiG/FTvMbqYs5/h/f14nZ43RzwAmP4SP5D+Z9A2yWnlPFfYTQWp7YI6+g5aZSYl
iD1vN5oga0/i9DupLqae8WPh8ORhPmn2ENqpN1DSzw3kj3XxgUTI1aZTJfwcmNERA+FudB50vCtb
tet8mMbzipP+Whj7zhX19vpEvkLV150iBu/duyUpgqj5c7QN2rB8d/PLEUh7QoB6gGjUSdAxddy1
dTvL/cVUy5Kx7whF9xCQ1rRM/CMoRY+7pyV5LLmiQxGSgv+pjr4Irveu/2Yud9+BdhGFUfXFhdxB
y5OeaaY34IBXG7ZsZTsOBwqJAjzftrpmragEh1Fg9NO+H1G9B2rKCzZbbymbio3BKLlr1rLEomv7
2x2IaY1tgoud2QuHKn8fk+j13hdcOTkEeihfNaO0y99aMAn9X59nHAFqt5Ts0ooq29rsunnm8atl
yyGfwo9TswpI3qEby0WtjWxNieXg/h+T69DFv4iwR9tiK7BUEXkpYylu/KRWb6SyYMSzhz3mnKEm
8yuxjGJMVDFq6Iddnhqt4MxX6WRlhk5mc83n94V7XgAd/LkQ8dJICW0NcYf2N6br5/YihDu6CFH+
Fcx/ExQHS5h59jyu0FGq64TmqD6a7n0Gxc1pFcqLCQwbf5gVzx3M2vcPJ9l6yG5Suw+ix5++/K5O
lxvdTdO44SMfIIfvr0ZeP+1+8D5sk/CbHuyCp7WeACA9qg7ujyji8h1+LSz0A6QPSM5Nf9niOOhQ
iqa0dAhXWxYktk4TCxjwfhavwq2kMVVRSGwtHugCVrzW65x8TJnWVfQ8j07qP5rWd1PvnsGCB5UY
Nw4NPDTSJv6MF07SY99vCizqrD3HHKGrMlCj2g4+U5qvdAQxE7hF7C0kO9oEoUjzcpJbKv5fRZAc
0GQxj+OfBpACnXbetEs1MGeSKN8KrhdrXc6NfqGflTmqH9h8Cxzv4baQKDq+RactSXFhfVdXRGDo
FUHXbmbgscCVA/RNwGzYAnYTERq5vExw7mJinWCSfc4CHTxdmPuz9KpdZz/8k/cX9cYYM84Jxg4i
oZ1fOLf8fgmrAMo/WeMU71ZfV1tCxEPVUlWQ8NG6r4UpDGc1vrYM9BEYYikh07X3cmzBOjIoQshO
Af5DiL9WEqPf22qJerhUoNThm2sEmbBQonXItDo0+zrDlSOB9oqnM1BqsG+5luTNcg9I9ahe1cD/
T87iTtvvHQIEQ8j10cTCYgHwS9d3mW5RNrs/nhdr8+nYSb5Y8UZzxJ88hvqJF+AsHUgU0oHl6pQE
KYGLrmxr0TSUE2LtF5UzUGtSY0NiLSCtA/zFB+Ua6QV60rpyI+xL1LNURgo2UxwfKU+PZIEnVWvY
J4REGW6B0eXYLE6yrdJacmXaOsWD9QFr/zFZV7T+1ifbP95nXq/r3lI7TbdbveKGROScZ/Q2UtPm
4h0UDbGUXuNidhAHM/eqfGiXUyd2f/hXSLmMoGJl7fIZB0HIWmO6Z9I6dlnSzHwe0ERyfIxB7cfC
ZlUh9OguZvP/MDR96odDyytgQKwCjcA3T+NZi/EascNYHMCkCO91Pvc//1kugX6lhBptJv3LLuLz
X84LOch6rLlC/QoHrY8WXQ5CpevJWK2Xv/tFTHdqZourRL2nGved+k5Ro0X82Hev2JmptDsh4usS
y8c6k1tGFbmhGLcYg2BlpGi/ODIkudvNpZSePr85MViS2pqO3LNb/zT0zZ1DC4U3K5c8C8MjJhNg
MWf/U1z7PT7XObEMCaEPl3cEF1FcYPvPqH3/OpglQ4fvF5rpK3XM8iP85VU9eEpiCOStsMiF8cr5
+tJbgnLilyaUXiVLJRmuSrY4XqHlpIgHQ/APLL2yZBgmxnycnNnypUYFxr22fzoFN9BBpRqqS+Cj
CMABciIqBM8kO2b6sj92txctvClPcyTWH5a2f+B226EQdokyGi5k521BssIwnxL0YJbg5TB0tFDb
V1s/3JdtzH+mBX/AAp4X4O1M3ScWaIVW/7pehQOTVEcgiXoSYQ2RweVJM1cSIHLu+fRVPcaE6F1I
RInR07fcK7TPrv5A7vhCDcw4w2G7OIVP6UsPHny1498t9hVM/AJJm4vAiD3ZQC1f0QG30/u51GuN
QGe2Fi3DtaonNemT0ynPHrFN6id/nrbK8KQa2dHFek5Ouh/7EcsUNN/SuHWF9a59yPExm8hqsEgi
ASnCddmWGtT/G8LTxynn+pKNTmeDxITEglTaWD/Iw4NpY0KaqNaaqH+brIvuK9+0qc9R66oZnLdH
CWacy0GgbEgSagepinMHXIAEosqQnQ0amb9LrvX4UpW/OenyWl/rUo+S79DHnsNaDxzCKNV1L04N
IA6cnvQ9KxwfWqPjpv64N3RkVMhtb8rz3Hv3IU7mBncdfHvwEqItfg68e3UDKByqKMl+zDHWBmG1
aKzaOcqvLfjQIWd7aBGBqNE9XnoBXsWhxgNTRVZHJb+Bqu0BzzDmfqo6hV2mFcWEIHAEAnupJcFO
jtPMDNd9KIoAKBH4eDr/brJya24AHD5ACIGhHC6f3Mw2pi9I6tSbZ4rYDFOf+J+Lkg6ckp1s5X4o
a2DkbV8oirc3ahTbE2L0AopSyHLpYy59XenGZYwi2juhv093Hc+tyu7rYKt/cjmtLe3rIlgkp34r
3xelPNhTCmKo8JOX/TJRjoybYAf37Ywb+SEyzXqKYHx1827FpCLr/O+dLNa2ZSnsDCoBAH7lXOwW
EFlTKUOqwSMJrPiFnCd/7Aoy3VTB/toNnAUTv73CZpdJE94vwLh1VUepRNFTINv6syei+o/cWkFg
/aiWSO+Aa6hpFh/NnQGul3MEUhvnNczu66mZOwpDmmzGhTvGdj/eWZc2IXadYkNADB3X2/9x15eR
uafsxio5m137nEXSMXMWovpQ0OazZnwQr+OcV2qfTtZYKhlQjm3Xct+gEdWpaFfdpb2ui0nILVSa
olawIwV7e6FLKlt/6qRCQAloeA7Q4KtyByeB3BfsKCfL7u7KvU1y1sYFYG/h6GgEBlj7+FnMdpLq
Z0pjCUXYuA6l5ve40aVmJsUmgdECHOSHeGIxx1ISMYuOHpHiY89TPQbnrLPrGvEzZ42vkSE5D5Pa
18aVBfJnzcJDKqbcQFUQkVe9lwIqoPn5mmhdoM/skz6ri6uMZY1ogtUejQN5sVigf7EI9XVG6tSg
YoswiddulA+0tcrauDeIoPRTNXBf3BS/Zp+hvB2C4bImZ10+BkODhoK5hIrYs4xddwad7duB7ZZP
CQjkW7LWYV6WT5VNb1a1Ja83WxMmQLftmsSMK2yTSCXcVTyA2tBtVYSVDwFpnc4W7NdARk9hoKEA
9WMKxAi8wfRiz5uqGqmN3536auPPgjmkhtqnrIEzPfTPu/EVLia06iTH0m72KVQL+gxNEOIfabIm
7e5WnHTZHvFpLiTETKxTsRsk77FIlm2EHbKLXtgwGD9oPNLymVbm9Fw2cwiXRNNTs8Bpz/XH0b0t
rHPn+JpmwWIVU8+Q3+84DNatEG3TAsDr1RWt23hvbEIGeQLqHG+1Pgk+JjOgEIk39czwCIYA5AY4
XCEuVFBVdeGF/exxDyh8dhnxRCtUriD8HiRpXF/rbLLAXp89uGjiXi1OGCV2w9b2hT3aSlxs+bzb
mURnQaCOIuUOB27yrm/ZoiyFeYHRDaVW9VSXYAbhaJbss7YLdhroXiMJ25/G3a9NYSxPj8usexd3
ZtnhRQ4XUy89qwR4YrF3V+febvObrE+wm6eu1edV4vf76QgxPzgRRhbbobvWzBLu20M4Qeukfmip
+PODcYWAHY7aBwAuCvZXbPg94gikgFbZGy0Y4G+ahq/jl8b0+IDM9WHyaxjfjNGl042ilZqbCa/0
eU5uUasrAAJW7HMfjcq3OmGSkc8bC5j4jwg0r7wI8L+eGJndm2RXtLScNmmM3tnfw4Lb61lN/uEv
Zf9z7wL7qlTKegCtz/7wx9f23REvet2Qzy7My1OAFknFH4b3qCgrkeu9YnWL0AXngsM77UG0tHFY
kfXXOpe7uYoECwoPLQRJoH16sPy/RGdQFi6QWL+dxvDZVhFLPIjEIp7CsQma/JswTtgq2sCgMEuI
aF4N+UXwClpHZhwhN3OajkPYrF9rSaSAFXsMPTo6qGTXsC8DZ+OGabLDV6T+Ipe7uY3pFZGsv2eJ
5oh5gctqipspRBxgU8kcTxsVt2c9dp0FEst6LWIuGBEJpI60UAv91W5Yh/zjmWdceApD0LXKxGLe
i20ehdsTJNDZxTH7VvTaQwbwI6JeK7TLU0kmhTx6/VeuXQnbcKCYmjtQWhdKcUc0fj3bQKHoYi4C
FO7ymtdg5Hb7VdBonao9/AtXaPFEmSChxoZGmXSoKM3a+JCJo/WWNghfxcDLc2C4xCnxVOM7Tr7y
/FtEoi7IlJtrvPeLBBBqZRp8Gwmta4zAn1VCi8gdomj22gui44WYJNu329pIWV05ksFQDiuDYzki
8KTMNqJ3/N4ekY8FvdiddQKj2lNQJqhwpLqZBwwpn2oEF4zlQSaKEUrh8sJ/Id/wq9ZcWWIFrGxP
9rN0V2tDZyH8eB7C76lUBmwk+NhXciQTTuliM4eHmzzJRL70AQ58QI3OEPbg9Afmut4UjiBH2LBc
fKs/X62yhmhmJtC21DHQbbDn2Pbe/+nY0rXT0pkSRL9Xo5kmr+A4ZHRy2ju2KyQscXmDGa14eJ+n
pMN6/kz4mDU2o6icHqn4iGZerhMY1oyJIIs41IdOxh0HYdXg7i6tX1TIotRY4YaLySHZPAP810v/
cPgEU4OWC7xe1mFRd8KNHht6fQKHm0fwbWY7X5MsQOQLu2sLSa9kb2h89gHCD+gyMIxL58dBDGrm
CeQnQg4Z1OsuL38W9XupxZhWXbx83nSf9tebov8iOcVIr0OO9MM/5f6h+TTm5bxlvY+y78BLs5aG
wFM00HuubL4/CFEdVFrll1yH/rSxkQpYcxbk0vCslYhznJFz5gd5mPHy99Kn2bbycSJR2MEuhO3A
LI6SMNDggkE5thCUIqmC6RIa0Qdg0ibdxaY4lgPGKEgVmFjZf1kift8TDt10Pg1t+XTiLWzoxCzs
U76emH0/L78QhpAAHD7+hqO7qQLhWAVoqmC7k8wmG9mGDdeMzTQWCS/mv2s5f8av5+7txgpF82+0
5PQ7H0JlgGSizf4AKW38RXnKU2LN6Y/GYW4I4fFR4pgDafhb2OSCJQZA7hY0wXwwvS7Eu8lb+P7j
LCUybY4Or56sR/5vJWPeBjo8+OysuS2C1CbtaZ2Tvli2WcGLcdg3K61dOthcEruwVD2aBJmUB0pi
6ijAYdaYNdPml3viso6zt6m/qDfF/MX6II72uhnn/cou0RYhbmysZU3LYgD8iKRose9iZVStjvP6
WEBCzvg+U7yzeqcTHUNw3qBNCGn1qV/DQDjYEt+wJZvGrQz5e4FMNaphKRWPUwhHqxRiNQDD0680
xgzQi1Uf6KIWl3kypshTURDgsgzcJfu+koAiqVFSjdShG6ny09epHluI8VOzKiAGkwtGhf04xIIQ
77fHjzep2GfqUMAq/Tww9+sar9AQ/pOZkPYd5i2eU37JVr4zqSp2ckeVZhsnGVoamCDAvw8zT6OZ
1s/c1xFSYMhxb1vL+StBGHzo9uPrqvYMSBpUJquKBqRNlirZUUlasADWaC1dorbT9Ohgdlr0LaW4
Qao73rokznmjqRBA7FvQwew0NKcImueQcNgTF535FQzkIKLLmrOGvRNiy22QmX6nYCIz6Cpb5WlY
xeNlSIrm3pv1yLif+yKRIcO9XDBfMRu6q6YdOM7JaBxtk4G02eBFrRzmDbdUYAshVQuu/5/bIoXY
pr9GSs4Hy0V7MRM8ETyGNn0Fsca4sROI03lv4W0LFJplTbKlL3chMqaNaMVRpL215pDtJ31rxob6
1N3eTEdwA8yHtA2oPQAXc9+iKwfy8nEO1Cqm9huBrq35LgRdeJWOE7KOZlL2t52HhnvgBXqMAiXw
P92LfhIEtqWJ9Z5oNVVSalbBBeA0lgOJ8dSUj5VxNpfhijcZrg13HaEZ4nOsbHXuHowzYefY5Ctj
UFHQ5mqqUeCtA/OqbCtuPxwGAEVzoputfcmtH8SVCWznt8vTjxvKBKfx0jgaDE5PeY2AwlsZd/pN
64anUeZUPdfczXk49FPsgFsq5HVtRlXATb9ySMScRraSHxV3/Ktd7aWSw014uxmKcQwG0sfB4E8Y
/ozZcX4vM4ZkEwO6TUwdXD3PvPv6YjS5vOshs5FdggvE49iq3THcf84hlZPYd1dZJ24rWBvvGfAv
d+jcA7bq2ZuYWn9MC1TGxBzpL2OZVe0XB+dWCNHvflSqrmKtWnhK8CsuqRW7085ljY21PJaiMc7U
k2TvGFnB001mAmGSGnFn7fLEU9aNz/yoJ9PGsH/MSC4h+/jt8lBIN/D9LN3/kEf1xFJMmyW2pIj+
WOuI4McZWYBwkZIaG8Lh7fd3urxOghNYPVt6FCBbzlQNhXV9EDijBq4SY5AKVmx7iLP23pGEkEJ6
a/UOI0UQ2f2TWKvdSpLIM1snHso/APBXxup8gArqO+sODLJk2Ggxiyv3ZQpq2OUCOIwcHahQq+ra
uKgZZqGnnqG4VnsZTH67r6cES6us9zel5Uv4f5XIhDuhOE6VpjZEbJuZVTIt+iK4hEcoRGA/ftYM
RapGgT9XMKGSA0+jQ0efA9HE/GLoGQyQWzbGmDqaLYIVGOPdDMqwioAv/KB1sVVr23Rb/SY1PG6S
Sp6s+pAe90raRuX+RF+3aEnMXr1vMzbT577PZWivZK3h0t0Ks/Z+4S5FktZn44kXc7PWZr0Xi5IL
odo39sK9BiqWT4+3/nSAimPWYMeJxj8+cNiFBQXWIMW9QqQIE5ozOVXugqnbceRsxs6ACwLPCmS4
zYgt7lMmiqJZhWc74GjQXj5Hjn4SOCT3Uqgtzl8KdG22Ew4EI7LAZq9NiiM7y4RcMU5W8+Y8q7Sd
frmzRv4DnjNSZaWNIZzruvIiBAX9ioti0sn9MY53hbSRYwRBULJJPmOQ4l5qLWsHU5dj6HQyjX+B
Rd2zSezFchqYslpCFXeKfaczBYfEfekkC2OTQq9UfXK62XVw66VYj6Ur55g4f+0D85GQLQ0aYMTP
Q0qSGOjGc9iEOM8C2D15O9RqXb6uOFiPvW7AVLjOFnqWsrlh8j7gPT2aUoaBwRRk0Dnv/kpmRAaS
7ZIiY03HeEkp+R5vFMZM9rcZwVEc9E4JDPBbhgT2DVCLQvIfsm15YOLElXBdMDDBhsE7FuhnPq59
Tp6ISfheTgaqP+M/PaYlChClOvecAieX6RIPSa8q4/ZI2Nf+YuUgtWe7uGBf0/uIEMRSnc1HY8tq
s6dDsBGXVk5AoD4yBAISgicvbQNUUNJc4op6taGTcY7RPP3JRAVh6kqpipXHJnMFKuG5y/II6KSP
m4pVT1Ae4Arv4MfjVzrWnV01W7TMKItiTeXOCbPHu9P4G+f1nbJA7SN+WYzoQZneE+EWAV2+84cc
Japb75pzhqTvo9KcHPqVBTqlnVMmrTlc4qw2S6PNN8XmDJ0ReB//g6vy3Ai07kc1dvRgSW/bqN0g
j/zyOXxu8xFqBmslz9/qUTUFbU4Ngdoa7oAy5BIgvSGj1ziUPjZSIdCUlKlF/wn6sMmONb5UP85h
iTJYM6+dvIeG81US3AmHPoRhvkjwP3jsmQq3XBaThiowvFdEfYM6BM4lY2z/PtFzr+W1gvqMpUyK
w/akRwKQHWcKjymt66+5P1uoGwzr+fYQhohZnd3yGpbYJOK93Yy42yGUhDMx5zm6y9CsAL3ISS0G
DnlSoaWR53/F5RqWfaHUGmTuINEY6Ti2ADBgeD0kzw2/kflFwwCNzirTfKtB0wDRProJMKmRtJ6f
G9KSC/IjtBRWw9OozVROxWu/a4Mb4Scr/qIG8G1AEWrtFW7bY4HsZbBARj0C0OeyIS08f0QrSEGm
C6Dgp2GjTUpD5GR0sTW067/NiBrQlLfZ2k7cJ8etOF5s8fnhyAEiU7RSCqtBn6SAc1CB4xryQCuT
sfetzjfvsTowtmgdqhqUiiKR7AgJUZB8qIPaIANFjXKVKgGEv3qaahJkgo3Qhgrz0nrsMHv/otUR
2CItgakawHq9OjV1Gjze4i++3a6baWsbT39O+AgnoZ08oIL037LXxUJgK+YhJl73F6i9bMliK2Ah
LiyIIkyKEtPCtcwRw44rZWdsj/gpbRYoTaUWDSK/rAnc57rD3yb/+j0VClRYAP5RyI96BxIojCma
j1xntH2w8x5jXzwqy/ep7Xx7VTdJQ4RG3P3c1rtlxIfMUuhiytFb/mMGiArJAeGw0Js0hwgiCqbP
lBG096kcr9MjXGn1oKlwhCokZhr2SDh0OgvqiPHi2H8z8iNGCNb4FfUF7A+sBhhgj+vlXjzvqk4Y
ypjZVT0NFXDKOQShaFltp3CwSPaa9wtWfGjDEDkW5clYg3o6M/p/eyYhIYm+OK/LEiuXl1RzdIpg
vG3tzdpXHKtSWBOjtdoKmiEI1edwEad6lBSQ+ao9nFScD2ttlLVFJzItTeThrae3IeFqSJ8WdLWj
aL9JsmAkC+lz2ePFZSbEfvBWgvSDwFKQQhQPXiG7gL+t6sfExx0X3JYYfzc3mt0IYZ0uU1F/9zmL
tpGN8E+dNdFEYZOgSNA50UtK3hCqdc4gKgeMSH/TLG8Yl79MCJeR4X48ysgSdH5asLSjuhWlPrqE
RHwWnZMpRmlWUSUT0DYO/tyGN2a9y+stBEbyntLRD9XQoxNCA0lTe5GgTQXRE/vCCfNGzZxRBmOP
1qYu9iPQ9dnhwrNcztLOAbFfrArP67ZEX+aTG6vtrGEmgfksZU7CPvbZJq4NR76ZYXHXrhvYgNm4
QohMipatkoku8J2C8PdIv5QfLORecFPmITXfZ0cHI/hVbP3ML2cAuQpK7GGp4JxZMWQqdSo8+vgB
yjQtfU0uJTe7Czq5jjcZrmYlnsCNhONLPGnw4Ijxw1J6sumQomKqC1vD6a638CFbF6q4CicNPZ96
U/wfeq7gdd5DQmbn+6sOyhb5BjtEzm9pHnbR7gUpKwSkG99gauZK3k17OCGSOdTnHwxHchKWC38p
1jb2YkNo2GGKAQTNvb5de5yneE7IgdK786KXmiWWCmXelx/Ay9GWvxqschsVcOLEBovgi9o/aJzf
M0V/hBwVxDT6JqfvzOVJI4eswx1o/qXtmJolbrG7x8ZMz3mmkqW7rDrOEbPf0lx7tgM82QdQ8JI3
qkasp229rv2TOOQQTac6E8TQGNzipIkeupPMDRJ2tSkYWkRvqawRakUJxkQjkuvIakPpCgxXphuy
lEHVSkQD10S7B7VMBIw8ZK/nZxwUnyEtQDnxTyUQtGfvmQJNM8wTwUIMpjhYehgc1WvDQwrOE1vN
QHPPn9G5V/TFCxcgEiBa0xXf4G4o2PZIaJ6unXPmvEJc1avs2LhSs+y6O6yMhpeNJkNt9YF4+q9+
RA5gExY3pgy8OMeJJ+cm6uAMeYEti1wu3uVE+sYoA6dgDOdKP21HU7/zdJegkv1yrb1C3gbhylcZ
tk8fqE1F0fOoVNbjKeHee5fXLCXRLR3q8Ur8ZlGLHguKK+emLKRUzSZsrrrfh6ull0MGRipRAW5h
uwwDWSjanjvv/e4/PTEucrL3OCfeOuSplvBPZSIW/PHL+vvoMXLxKunIF9V12u7YTUCMFSXdNVgM
QfqfKf+Le/2alDMmYvXzAQBcrbraUTjbiBz6wlY8Mozc2+AbAfdecFPN8Br1WYnYtkPMiCZ2nfmo
abYFcn0unAmPmUo2UGUVarpOHxzt57kAXLtuN4SkEaiR7QLzHsJ9YsN/Wd8+DeT5LI5ewU21v3O+
mseErjOicU2IudO1cNq/fjyxTUTzKg123YoJD29bo+xVWI0ekM0Ur+bz1/BsXS1PMgu/8rzTQWM5
k6uhqNMmrqYczpZ0/hj4uNkXgV1xUlrQDh8c9voatdnG0+05LDA9jt+xmIOSiNdvP6G2s2RIXGfM
I130dDLMY3qlkCKQz5gQdysNrrt0L3GGzQHNMIod8uHdgGxSZjRBPRgWC6QHSZ5924gDn2ufA5Sc
RYKkssKZi1k2dH3Kh+idREHYQ6otR2LA1VlkoYYHqLkuOlDEqy8LWvGKtEnDzwex0ag9WTPUmj6M
Ef8p9KMfcupnJLr3XcqZLgTzJiI7l9zgp5xNxm6fgcHFy2tPijaOO1+n/ElCDVTRXUZjo89LJ6J5
zW9ETOhqlCi1dGsbo9lOw07Hay5ee0ykIh85ykP+89KXtcp/IJqismc7SWZGCNUtRUW91/gu9unP
yC6F66glxglOfVj2t4apS/zG983aTgE2TZ+g7UxugJzyQJePzb+4CZ+Q3x91qFBlZbDJTQfxQJiZ
FsfTOhTSx5PMbyDNBl9pGL3doRvZs9jqum25ttvEIEFg+JIod3K5kukGvucU4aZf25wUr9T9V8+q
A5OAZ0PYsazUI2ETSqhXz8/XCMenAjcsplg5YAo99+hnpL6YrUSUGXxq3mnHchlAMaQwp+x11Lc2
W1mKPcOSI/F5cA0Rxvh4mM4a8OpewMeoKzxj/50crzmoVN3FotlxGBEKHf7F6CI7qmD02O/Y2z9f
l/i5HcYXBGu0eN9ByI02ZxCuqYOXtlta3vH8cn6y0z+6K65IdCVDkiDP75ZyDlb3IUqBjT1tJaxn
F8aJQG3DHHln4bleHjI9ELkX1INjSLa1RV7YOZ79XO07iVtkMFWHxkyp1g4G0mzjOnsQCz3tgfcZ
NOxNRhqAc2evNlPSnZi6kfIYQJk6tzvtrvUqqr0YmErcOok1UBhx8lgrlQNkHVy8Bz2VDpGMKtjE
YN7fsC/90VtG2bbFAkM0G3t8eZmlpUMZEjyuq2Z5ry6lf9JaSDRXLrUCmVdRQHlpAaoBrxmo4chl
lnOzfPNJRTTE2uCSFWnAy1x6zxYHemdMtOjfvFS6tUlVSm2ykzpEKBC5swXHnQK5jUKQV6p9M8no
LymZFUOlUTk+o8BZYmzb96QP7Df9wYSCJsVh+iq5ZhoAfQI0JzMQtVPGtSOCfwnPYkgvofSaoC0k
vv7MfJsEROcOfTT2UT31Oae+B1Hq95MhBZhGWS++dBSMX9NdRJaqAO47JxJeHbrxqFAjXES1awfx
m3BPCGGUUw1/sID9gK9Uj8y0jmKTTs1Lu8GDrlZSM5pYGXxqjPZxi/wVzBTw/YFop1s4PNWsUemW
ojNP7twy65Fw3i9x2Q84ybTFNjWqG3FGXK5jb9NWWmVRQs6nzaA4oIpme02VMyr50kzkc+1ks0FG
UM4MVQ7Oo68PX/NSy/cW/oyq6wnLwClKcV7mIniKKead4AwWIYiRbHblXQgdku7ZL5Oeph4cBctA
uQl0N7/vjMScay55Bf5BlSJqNWB3wXijTxjXHzZ6TDcaRaeREZdTmAXCnE8EbKDRObh6wEi3mite
URoKC16jx6UeTWOe/KwfF3ua/7mepAsSFaFCcvzuNeNlsbGu7c4TAGPrvmaJ5sgObFfE7OP/aIeE
Ar2dHk4F3D4a87dVnNxIloSnO0YioBNQnALtOxeUzPmIjbtNKzgzcofWMAxEcP7c8k07A/7S6Orx
O2Hgk9n0tnf5JPmYt2M9V/5HzV98o4Ier2qWDAWdciXQuL27/afq1a+q52llmmdnHc4WTZ3Fqc4m
TsJOyVuh3ToH+EbpQRuxDjtvJkM7wTePWv/X3vp/pOm730tVXK1Vv4ROfSy7LSUUOHHnbAPDFHsX
2OObO9kuvw8HCgSQWI7mkS9GFnj3TJh+8qW5BQuxSlsM2Z+ASuyKh9VAwHPtsK1RCRcV5AsPrZT2
SZtSV+l7d7lNEAVYW8ycX9+W/6VIcrRwCimLjoKPiHMMLoj2iklS1OrcBrDJdVba1eJ2/Qc6plxe
2zWW1yi7WLtc/umdQKLG0LbrsGQP8ckWg2TNopZk2AF0YwhruNG57WBNjt190QWIj0FkO5ZJOlVy
1EkINJRCAjlh3ByDdfL8jKdb34Y3+bNWjldWRGnTcei3MhwfMXIrpVitVWKOFqcFv24T3XKzSJRb
gayCiXGZu84WEKZH8cLRW40aIwjcohjxd3dmV8lAtO8ufa36PB5vMBvAutmc3I2Im6lP0gNikaz+
osXjKHnBsBnHjbI6OjiZd+Ki97/EzUjdZyaaXeSGNtdia4UM1TLVWQeZBm3gQ2xulDfSZoNcRHn8
/uHs62P1XPAjJQ9nXCbWGBz0389PwOWQeHm98ZusMbA0KSQEDVDyGxvDbPEfcCONHw2NF4Xmw6N8
LdK7l0oC9WnUJkxVOitKUQ0h6evauU6huM/QtflPappcE2Z6XFGW9C8xPYOHguD0LTT+hLrd+sa5
iGd35YWHC5qDH5PYJhDoS6GxeMZXymqOs6O+t0oai9/5aWx7s+9vgnIgfDRv+dXtXZxIn6ZR/6ok
RJpUAyPgjA3AQvzBBp5v4BY8piKtwSoqIwLoWLH37bCVYJtZWl5icncXqVQjq+VQZ3oBCBGziK1s
wOjd3ZZ19rix6y5tVPi0JfO+Pt2+v961KLDLiMhFneNNq+tN9+afYAKnturjuzhHcjsjV3II1xct
hc2gMrQflhprJzj35oxF0sr6Prp1hR5cfMWqAoNqNNEpumVdqCLMcCwmqBwH0IO64rOEdO3XyK9I
uesDuxT0tGS7ZZfp4oekOq7bfnZLDU7WqVPOOR9P63CwLy4LCJ3dTcqmjns5oMxsEm5QqM5869Es
mu9B/2oek+cLuRkA/xEV96jDKc/qaSTxVhMGFKAAeGqtnjkV3mvC0vrJON7kP55iY0QBdj8hgfEI
410JWRR6T/FWwZIb+q87wqiFxNXZVDMyc2aXONsd71LFOO1oIBDmfSHbZs/yjtlqFp+ZhdXdjDk+
yX9j8Ns/V8IRQqe/BbAdEyjaj9IHzEV07Zk4DQTriy30+9SOcPXYzf96xzxrr4HmD49tOg8weuNd
Oy8d5Oh/HFe1E1ewAa27zJupgaT2xA80S4FNOPKZR9VmwDC4vvyJLhta1y409Yvmwuiio7BuzfV9
sCS+FSAb5FTWEwxzW9z1Nf86eaP0cpP+cLc3s6Yi0gve3khAIuxvEhKEGABSXjwZiU5HjYqqPl4w
akVpZUfuxiaUY1fyAoFh8yuOxSl+tlpmwpFEOVRPRD+rVP5yNgXs+pEuQ4La+qbrktyPd5lQ5gqq
p7yDv08UKgeDGihh4T3xjHwhMpbQlqjakt7SbVc2II89hoTMWmZ4j8VgWAVL4IirCfsZpt5oNIN5
7u6H7uelp/ptn+jW+28t1MjBNe8wyaFsUUu4/BYEv6hHJCuv9FMUL6dPxGewLmUHhRL4OvhCJSM/
kI3v0Udq3Xpswli4hbcnHtAkdErOHSI08lAnThFouZYwNNVE/QRP5sskCe/xZncoj7w/TnIZEMfA
hfjNYWp2BmWSFXxfHwlo5MQJw7YZF8+gYLBkAm6qwK3VXnkzVBU1HKBOnfZng0umztSH5CfzyQgq
Q0buawFKrrjtD7e1en+DBjVN5Ut7z57bNKpZIVMMAxbHbk1fSA9v78jqcr0gzj6DSmdoDkhe8euT
puvt2D6e1gqxHuT5zHJJ5LZQVCd7ewNiy+a82PWQerDdzC+1Yk+VLFVXRD3oblL6qCT1R76IBgx5
WTDlDs5FNyDoUYHBLr5eXhLz8J4YxRw3RUGe1Gc8PVTEt+EU59a1QfSWAGfpBDWZ7TLR+uv3HP/0
ycDic0PDqXeNV9YAtDvMV8RHxmvMFK3XK8yIafghJpRFI/sOMfJeD190QpBaEw5l80j5wkLlaXQu
YdNDcY48ZQ35auiJOmSx3m0hkL9LuAtafi82sy8efzJmID8j9Br+2BORaS9X9tSeOmrQxwf0wWzb
oy1iYtWl3hsX33kK7N81x0CJ0ebkOzzT19ENSf2AbsiQYlLdZba+JgypTcu8wUCpPdWMekpQARSZ
GEy4jyicYUQ+UjXwNjZN9Jj4u8/5IDEkNnQ8MM51OKn4mwDFRYztDILOhFB8c50LYyemTgm7477s
3QXFAKR3djy8vVxo5WBUzziiQyocbpa8k6A+K07b6ONYwuo3G+I4DDrlYuhKPjgSaNIIVsEY4wDU
EAIFnDzrrG9TBzD5ai7BpizOuEr1864Y3FIEZqnFI/p3MF/m4jsOqFCg91vViOWl+vZMQpcJNUAA
cirPiCJj2yEkobtQFlO+E/I7YFURpS+oKDwQBBRKnGtnyvGl2yuSCFjmXGILlJL5pyhOeT5n9eoJ
gsGRozIeMrfJlgLkA+e20avCxYSvDmPvSWbmEuD6tS8oJNhMgVYqwWjzjGci+FGnD2y/f1RJwLXn
7kgY5xYH8jXkgF02KJG1Yvb38MyUuga8eW98ia18910rd01fgy2kH78J8OTcB5HgvaSG6BdC3krN
6w03nNAg+Qgf0SAkzIMugOhZYJX6RqR0nAb41NUzvrIgACLfpge+kVnjjv7FnbFu8ahWl74laIVm
kdR/OUZCAqZ9gXCd8Xk3JTXqOQSQn+MTWa1v+pF+6u4RvNm25NNx8AeWV91PXeQZkTqYS1LJQEUX
RO7szwG2i5H3uIa9e/6dSpLoj59oqCkCpMlcXvXer27wZe0sJSHITKrOnORvMsmE6gILKb3Gs/59
eK5gxIVqhQ2Sy5qEabNwBbDPOr2/I/PttA3ZbZkf46J2xlv0XgtHdANPyivcmxIJzywoNpQ/nvNe
WfXphl9M/vAKP7Lghx3jAds3xyOyTILbvWA5dXFueRQ550LpsqU89RkwY91zzt/h5YLUgmDcncel
VwJ8RCIhV/iaJBVRGyuXutuXvDGtcQ9P7LGqe6+DpMKiZSfh/m+kzSHlgQoHwdJItzWyKRggQgF2
Jmc0m70Pd5jRGgBAGDCPVHs+Q05odFhZW4L9PxWBhcGx/KotraCPj6gd/yk/KhLhB7SDbf2TYBL4
pf8ZBtZeZ3dvYP8ieIge9THte0nZxd1Xep4yDixn7yBR21Q7bGTiuql6J0biR6kbyd4UsBSbq4/G
a3IQC9RYzf9FMfA0YlU+OXBkAauJibd7igRzZ0eNvZ2wpYQT+/pwCCsX97s6Dj1dCpp9TDclXWEg
uiox0dJXObfxrVn2hY+ssjNFUDSYGWZ+RLpMKMtES1wDCbh8euZzR0ElDYOpYBaxIQ8RmFdGzA2b
tazRWCpGyFSVUuAmc/VmMTurNjcaGNK01ZwXNz+ViWmiDMjzmEwOGGoAbsDULj3vA379hfJ4X4ab
WXXdbTlv0BmIRkvA/iiUneXbtG9+EFfGJMnuwRhDqaoh1Wm1tY4qIlHrdtNepMYSgHjEP19IKQ0v
tO56I5geak0CkVKssBAe2lz4PvzmIidpaijEaLTlkCE6fz82Nl7/z7Hg8nsLA0PFSwvlzcmVQcLF
Xrq+EqVnu8Ppxm9V74yDTevR9v0YV2oobtU3RsqYE50vKdd1KKpCf7X1wwKaFyYqcf5O2FPtSOnN
kC6vd33jVr52g2CfirkiLW62bfUIccKue2SsYHJlEmcm5+8/uQRF2rulfwQZ8IRR+vC2tRmbP9oF
Ver2BYqW4HxuD3sj6C5RyTo29cPgpdBBo4vIWxdDnyVmiJUmjkO7Bm7SkYq6hs9th6yqJm9Q9dBP
0xVUHg6GcdX8deP51rHURa/EcYfPSWod4qsQ4d2sX/+k2ZYpCOXvrdLVAiKSertQKX7NUnoorzxq
bglN8zr/y4I7zmLbtbBKO6sBk9zcmeRRAgiiuCROCxSqHPr9LPK52WqSyA+DVI+RvRbZhkqHu1Nd
Wyi7xkvXM8fkghNJhao9Dztx6mYCXt0Kjfs+1O5bzKK/bkZO0753WRQfjrq9fAM8GLWQRgUhoe4s
24i3eiY+Bzn0vcDmA1AErcEAW+D5pqP6j89tg2RaUJEi8a0TZnMX1LPl8Au2jwR5Bn85zk0idfIJ
4OCti1SjKvaGUi/cUueHt8iKT70IYSoQOOSp23mcK07+A41Q6Uc+8heoOOwju+i6cpSpjH39UGM+
J8yl68Ma0zfFsq3g7aPBrS/jI2VjwpPkwM4aI5fMyvs1alInMgApOGRwvO+HOOvBkJcm+SWCWSuG
vUCPu/C/mRAx4N/mdnQ90H2bysCfwiVsDgqaREXm9Hv4652MuYjK0iWSJWQh2QKo0YK4eEudRFNW
CNV5Ylg4jiGAhnph3Zm2f2rjy8ZUHiwEpVGzePfYTwth++1kB5Vhmap4Z4TVWI6M9i7dDa5q98eo
e8FtZbL2RpZAsRQFz/UdC1VxEVEEM3cDkMMIADaqN6FRUySez6J0CkqaKFoxmBeIToewYyOiK1BG
Eym8m7etet10vvFjUaooGq9f7lWgzGItPGAIRg6eKGHya73g7Pmd5IWuZDQAYjFU0nXUZwC+txmK
+4drxaV084T95FzXF2leIoxPgVFzgCx+Lwm4pO/RRRKzox0VBfQiAaeN1a6Au3BEkoT4eEn1y4/7
KweFUcYnx4X1ozoIt4FoLZ12BdiCSRFWAQMwtASAYkLfMnTVtSKMQyNYIebxU/RKpgJb7H6TUnbz
PzOYaETKX3jogmZ9Clwiu5moSBc0+dC34/RKW5U92zDbAVTwYWhBZeWXpUxrEIyrpBSjqxNuXt9z
R/ibh5h+TnrEJRL7uOdZkAWoZt6JGTC3uEfAm2yC0fWvaL2mI2cmXBQaeWbQjzMDR2oS7mo3NFhj
3NLB4puDKT1FMikesMHDa4k9nepUeTBMMIioeDRyW8v9OkvCSberNRuWXnRODZq5qqsjCPKV+D6p
GQvCnRjILUmDhV+eULw+6A33EYU0p36SCfGWgMLhLNVqsqWgLXQOJiQ9MQ5vlf835Y/8u8Fw4CEg
q0BMVjBdE33MpcJx8gartoe1iRJuIhgp1muLWaD3rQ/qBxEDS7C+FLPTEvCuwZWFiEfne2YIXw0U
njL7HsVKz6Fe67ZVI54gCeeA66q1RE9dgMEbYfDK5rFxkbZbv22wjaa0X0k9UF/kjvnCNbUe4sgj
a5is9zlLZAvrtsNq6Ft2hTKrIpqvTyzapQYd3gMP8WqU1jjxdRhQhSP6VDpTXr9/nkCu2OjBtDes
koTooaju67W3Jw+eEHt4HP0N2vPxFLZB0PjPzlgZwT6IZ112ja3bGrvYXUG+tEMqOF4uRcmIt7h1
MONJTYxWnW0M1X9aNzQSGQi0hIGyq5KeCwUMRK31TcdHos1c48B7KOCVR/I5I7SeK6v2eanXVR20
GwRRucnHd7vYzHjGc9wwAfj6sTmu8pEPWz3vO3p//mSt/+Aalipm2ku8sf3uu47LzkXh6NEQ8Psx
7CX3vnppIg4gv0Fppr98SWDuH4ehe5/Eh6lBsPRJKfGJdmMZTUCyx2SCVBJDSmacCFQKN9xUm19L
Q3MqNYjEU6rxEByS5qha1ow+1Fn8tgCfZHr6L7LxL6ESj++wvkwd8XCaRb9GTmfpVMYfTyIzNhAa
Rm2H2g6a+ml7ajuVwnnPg/jwgLdGwJYRv2j0LC+oIb5QNTt4NPFNuMZ9UxZFnaO3kJI6QCVApV3L
wwb41H8sI2fsbU0vC8GNmisTZrDT3R9V0XuSep/u9wsBizt7Le1eBI3sWaOxR0SZRrxSW8RRujne
cSvatxLSDCGFo4IOMtQ44BfBBDajPXJek5dW3PtgTAEUozfvaIdPByrFRMepTJVXNlN7lrRk5MdR
GyrT50nySKvblLU9Fom6P0wC2PKHFxN2ZayZrnpIeR2lCtU2BDFjAM5EK1CWV4z9GIBV6vg0gbzT
4CzIJt8lb4F53alHLotlBzfnMsX8nD7rJak13QeVyyiX8uBtFF/F9BHoWupYU/2kFLK7knwDlZXv
FnDAvbVbQAr4fo7VFLQ6PglPjtdrufDMSbATrlmRajVeAFzeaNzYoS9q/XwPvqnDZjL9FIt1Rwu2
+XKKq8JtolrdJbj3VCAmiBdHnNC1lGMvX2lClYkM2I9NnOyrH+R3oZgoi6IHt3l2bo2UudWKBIiw
iYQQrUjcNVH2qJnNTD6qBqMZkHzWeiSGGQoQZugmjJXfayCW1g6HaT4sX4ZhsBmZRvWx0PKOUjE4
FdbTlvdfYO25nr2z1/ltw/p+iJd0xnObxokKtf4qUR4WTo+DaClwpu4Xjqf79Bm3L67/HAeUlPIb
PpY+Bu5X38zThhnHQjO+Ld18KmXAPPkpDMoM+Po+vlUyi6T3e+06lwC0vU/SS1lsX78yhBjrxUw5
k/QZ2pLugxIgc9R/6UTPjBimnVl534GYuF6tAe0nMBk5zGz6yAfdIELl8X8lXxL0BH9Hk7xSoCb8
Gfj4Fi9oFAI+4HgcFInnTFdnmzX9IYst44jQq2exT1npBVSNk6YNTQJqBMP2RblbKnsxb5/18RxB
O7AmZW0mOnekL0GvZZ5c98dz0LWX3dJKXR6oqpi8k6u9HyI2nijU64veygeromicNa27OUJq0y/o
tnKDz8jNKC+q+IcAp26TJzZXgTNg7zh6azsbrOmVoN1WTE9PJ1R8tTT74s6EASF3tene8APKGZuf
Jt84uiG9/QypYXjXQwG2Jubjmbe3MI9jakhsRZGsAEuF+0C/nXBuae39YQZcZMNJgap6/rI7ONL/
Npllo1xH0XzoIDszftIa8LRqbDlN3+FaIOvaR2O1NjKVf5MBpmNPElW+px/Nk0Oi7fgUvH+MOjnu
NxvG8Tw0XAx8KjW4fTB8F5jQA2VX8b2Uh2mvNaQZ0lW2y/aXih5lzefB8xOF0fe8B37cAtu7iEF6
da/2AjGYHjRR+hrAydQQTXBFjPoZTCMeOckDkLESdsJzqwqUvUxE2dOY39ekap6y5tbTgi+pywro
l/U5/VMqtDirZbARSDWw/bvJLJbXjQhyPxpOzQr/xUv2KFlu1L9w7sVKr5t6DpwG9wUo/scxUXYH
kxhCBGS5+hn0jMt1lKbNDyzaB+Kp1r90ZfF3I+zN0Xtly9ETQX5tohwXI/VDStL52jYltTb4dN/e
lQQ4aR8j5E66BIPpIiyvQUCCs3/6K4kvQGgrATqQ4ukwa1jOnVIsE1MmJ5zUEbpsGORqMeL/faQO
oMT1XrJfLEIbUoNAp4UZREWUCA565P+J969DL9/srIMm4P2XaQEgfEMkAcxh5aSQMt2cTNxKELnv
GYAFZzUXYJ/KcavQklITzBnDnAoY0fsEfQd4nELvt/AVuVHMi70B3ZMFh2/AzQs+T5GMvU+SdSD7
DF3O2Y6vtaPCdMWA+812aQnteze4WOmIPghLY+BG94Ovw8mDdc7I/dQF0eGiJKA2REuihECVuc7q
EFTWXhaSAflV8hDhBNSjETNyfcSm9mXWyVT4R7uArhtcboBUEeH2HA5MPBnUikqoRY7UqcQunrYZ
bUsvyd9wIb+uDDsr15GegoDHfiTnGfyE5uW6Qn2Maoc+WjmZgxMg+baIPOdCcV3M0VZJkHT7dRGP
edfxUs1GIV/EuoSOoz6UtpMgbhNqUJbGzf1G6PvCz209zP4Md+KZ51awBy/CEydZRsXg9JQ7WeaJ
+NPMKc++DcPuwX0o4+z6EPcvFGuZp3TbIucfBH/7QED6ugw25ln6nYWSeEVY4ED+R0nLItLfGcI/
1RqV8Je4l1kwRRKQEDonte3RBoGtQztIGD10qLmE0fnJUpAnWmFxTFIcgOp7T05Or67tZJ1EkyJE
qdPOTCHX4Gck3CyjKtRucFVa0G0YJST9J4cgz8Ry/3adT1AkuDd62U/zWLIl8EzqQ5Nsmt36CX+u
yKNnQnasS6ftLr2ZO9PAS4/TcZhDmDEY0ST+zvcCr9rbiOzxpWXAgf5/Sqr7f1d9RU1TPjhL7jKT
xnLZvmNLeMv0K3wLI6ddrPhWCtfswAJO5difoIjM7kWI1Vx+T+kgTRr530c2FOi6BuqdxJi3zlwu
5g8v3Iz/GXF9IXDgsZYy3uH8DQxykbW52Z/wrqTAjrwY+LsubXFf/Cs6EYzmCLCSeA7PNVWcQ+oX
Gob0CJhwYM7cqouljTrxYHfIhug8VR+/amv0msNQ+RvncFK1jnGsGGGp6JAHtBvNn+mVhoNoSHWY
WBQtc3MGdAt6fYkswabR1F/RYF7zqyF0lQOh11ejxwiFigt6Emk+pZIJTNOFA8LMtGeDRdkYzG45
WC7HV3OTkQcB7JYTtV3J+WgD17TAgx3skX51Ykq8wLElZ8CBwOT4jFo1fFKfiXwOrYDqZ/NQ+b/C
O902hMbj9kVJ2xzkJjH+PivgKfiXsg/j/kwEIus5jVEY3X0GFQ51GzPA9RYIxzAawD10EqxKLqoq
o2EcD79ngMP3rh39qSj6Usn5Y+8cb2wtQ/krZFFdWA/uMocmORvlXm7yTm/KKsz2Fq2IPIlrC0br
g04Fy4IZGWtZX3og7esGPNbxIZAVpuRM9meU4UbsU1o6JX1WjsroCKCkvNKmFzdoROo3t4M2Vs/a
EM2k9ToBasrU9PrfY0k7HC+KsX+hYVAUmQmOCgX/JTDRC+RciNX467j2+UUb9XXY1ZBOh0r/e9M7
VMyWcICTuELt/QnpvDVxMe4OL06lYMYHxhzDkHhw3AFFsBVQ32rWY9lPFY8N18qw3/YfypxgK1m9
T3nALidXnH1WIlOaGkZmkKYzR8J0LIB8hok+3YV7ivn0ojwBYN89VQzOFES2dZFkbMODosWrxa0X
WERwR3bFEfaLBcxyZIK++D01DYOZubb7G3Ph6I7xeP1Pvf2RqsNY78WeIncMsxoIM8yOOUZzS70G
eA08seWk9nwpENAM6VSAbDaDaMfk6G9u/l4EPgf9nf6ElQuOqyaudEA/0k/okwRE2RYncHivZSou
5siwibKBwhRAelkX2CoReGJjRQ36vIExhSaOa0fqgnogEC2Hn3jJSPSUPRezBLuKKcmRu3hbWw2M
86VYrOJFTLyGtkEPyuURPludJFb9l+wULA1v39XTuS84YOegE4sSqp7t9FKaglD3erJghf6GLZDN
AHpKv3HmRCo5NXlH/P1jb/NTwJa7tRZPTPpYZ6QdFtYReBgb+r8MHBplrv5JCSO0cvycc4AC4jLJ
NqVMStHzxMB+6Tpl9AJmvtVP2aCeBfJr37iWpKw2+2IPUvv4DH76SsuHCeDZZu8ZD9qU7J6jejXx
AiJyGAdgyyzc5qqg84v/QRONYtnCZR4NO1aR9WJmR6JrqIjIK+whe480+KMCqR64iCYonNjkyApk
QZRq/BugfvwmGHNo8ekwuTwpK8DwPdt9mODIfQeuoDyn1cVOko4uU6vD9xP4fCc95gPdfRKKTG7Q
hcvU8YRh+GPpuNFUgi6VqeNcpAUMfz+nKXe2NJpTYeggMmTMvYuuA9j/Xvc31yTSG/q1F/8ZHpwC
C1dGJYP4zJ1WOHCLaVLLmAMdtpLeXfPfUNkg+aHaMrbhgDWCgFMoDuHguepdoATiSqlyrRFElBo3
w++YwqW+22F99JJ+/lWEFEJ5tT4d3OVYsRAp7/qLcxg2YkMPo6nZ0hNGU3VLFy6AAGSjLHZrlDZx
XeJ4kBIU6st7VLx7wtGJejo+KtGp09jv+CdbRTOfRlmDPWX9bVYlKSu8OpkT4Mz3DtBzq6iaXzE/
9+3vS3HnrdvHwlG1UUy38j0hQLR6L85mdGw3h6o3yztRuFTj6MeCCdBgzAHf7xu4DUmo/uAMclPm
wfTDS6qHwflmwR0PMoWo1S80u9KjCUfMeNlaDFPZRUYD5fLuLn1xsWUg6dlLR+AFm1XE+dAwIzSh
KNXe1RiICBIWmIlH9yoH91sYlTNnHq0ZO5HiSEhGuN34YLbNUl2T3JWdIHplcDLPb/+28rjHyWjN
JFyJkYahkGZyDUWYe5PYzvDs1FLJuLq/9K/QSy+bgxqCEpeAbYtcgiP9EdWUieK7G8g+ovVDYAkZ
d3VOl/adMqZmoUt8rxzmkqIHf63JC43nHZl6YUzTTncFYivbIiEbykJpyxJ94hfePy6rgH3fmX5T
jMJLuKQDylpcqwt90VSNzyMmwzRY+ambXFLZ7XFfc+md+6BQGI8Yg1J4Hu/fXtavhLEYBovUpZ2T
SWucG1PORJj3lPhyIdDfsh+xPRhTRh0gFTmayBV00EajNbgaRWNROJUdP5pC4gvEe3YLoAM9zBKr
zclsGkdEaKqjRxUlJcESNkNpkKfLGtt+afWoGnF5B+yvrAKAQevAsvUQWvJ9kv/s9T8VnfMHAvIc
Z7F0K7tNmnA54VcivKsdfx0YLxHJ0MwLSNw4TbMNFb9++Qw/mKyIKEFHpYaBxbGvdS2o7kfSxPm1
G9sYqQfQJszFXwexi1YEROPwFZR+3tk+WyheFYxCbLEszqHq1hbU0x4T9fquSArix84K1UezvTAS
xc/9uaQRkJ6o1sc9V7NlJbtgtjiEnPEGjJEtpLaUEZXTDLtaOGXxwwqU3wiHohYkzIi1E1HJ+50n
/vAXTNx5HB13owe3C/qiMzq9HMjPP0IW3wAIiFZt5w4lWT8U0lH9g0ougfjinpBrpdSZWJ+JFYM5
ON6cFI+m+oLlwfolMILuW/UYBjpokHU0AklL2n//OT87J7N3J9YYEd9X91sSsE9Jk35S05z0AZb/
F+2RJYeCX0nHkbLgK05rNfa7Lf3KzFKaBjNs68FOtpurpZ3Xe09hYipdy/Rv5I4WY7WeCrgYMtSE
oWvGxbSTJCgQpo/HeutZaDU2NtjOg6kZ1lTTS0ruJJdNElF5rKLg9aZbI8FwGlApValcjX6Ms8XA
LcOdnDRzd8EXIRJMw5SI56Z0BcF6JLeOMIu+4oIAnwbCKDV+Wvuw8yejKU3VWyilwCHn6Mggc8Us
60TzoIYKkJzCfDF4+HbbCgs6OkpEcQnR3j1JgRbTMfJNJLBuBnl8FbZA1Gw+gVlMjvmn6n4HBJz7
PrH4FWZaBUfJvyGGb6CnavuZEYf5AafrnoYh/JLH2c/XZbqkg0pssJS/Tmd1gVg8Hzrn+6eHDY7W
cq6XOYFWndt1Y7Tz9c3nWZB1uUq8eFvJKot/wKI/4/sB4qwo5cP4hRdVt6KKWbXKWzlwzEzS4oTS
jjUUX7FsC1WPeU0FPVoqTE2d71AACH+NFgb+O+LrbMD5hALqCZrCyI/FNh6IimnZ8oIvdfANEsLH
QhA0WhV2saA10IzQ8kSJxMLMUAS0zxWhFOtvIJky2oGJ3uTcnHNJQDT3H2phDZrWYhQdK0wEtv2N
M2655vRmaginaQGgZiLm+7AYcc7vm9yhETOx0wqO0Sm1AUSt9XhNZQtZkJ0Gdkpr7SYwMykdgA7O
i8VXPTLP+3m1exZuT4bbF3K9vldJWkK8gUP8/EicZwhUKieqlvXlVg0j3+ruuO3mB0wStA1jdMCh
4LPXbobGhppGW5T6yOl0qUZk39V2Y7P4WjFH8DQ0CrZlFJ6qkcK8u/PGr28DFSiA6uS6GcrInWj2
6Wn4T4J/HmGnqZSKKCNywlLB/9zugDAzomdoOC3tqs4jG9wXJYt2KeQCJ1m0dVP26J+ochpzI9zG
V9bIOOXstM4iQSLqq5J2ybdJWC14q/Zc45C+feHNL2FCfKWyxF9xBjAKc0J5/rPFDAlF2jijshbz
pusabyKTW5ao5uUprsgFgfz3iUzBtrHIkuSauYRH0r+LQRx2Xlig8jLUmagTPxg+PIoD/luhM465
hBh5PlpD0n0g/TP6iRFKUMGGA1qgSoZK1nDE2nciaI8t8h1oCO3FCiBJ7PYbB41BFCxbvGM4I/BY
rWUxGdlofOcGormlpNlEylmtfIneXk92yNBieqI7m+XH4FzScLpwt61lana2EZ2wQ+fll6o38kpc
gwvQc/UmyEQvcgvhuc+/BNG+mVUQz9T8xO7OzPD3FQMSX2wn054AaWoDN0TAO2msZsDHKkiEpqrj
mW+iIczNc/hvVg9yn1bcycD9pTZKSv30JoTJB06pauIFZ+AV97zjIW1Mz217Pb5yxIrqf3Z2fUE/
gP+bkQau+cwarpykKC6pT2R3GAwC79jVg/BigRwoIvtXZD6hxcTLUoyM8WHFQfW4oj0/MkqzYq+S
lRbTN0w8uZQeCLgiugj9rb2BUnuKi4u9Yegk9uVIH7Kfzv+4NYWfG2MMxqyrbhChTuL7F3EzRwm5
X/QGkA5YPxjK9IR9fSdg6XF69jd0Kr6iaNdhqTDZhX7/guXQJBuMvBaua6ch+VaYrr9j2278veVI
nfgfAM4HTzoAiBDVllZ8z8veIiLb3r0wmY3TepY12iDn753l9nFhgWTXmUJUIAR4YwcbFm8zkFAi
Lo0LYKPNNVJIyOs9H9ManpL1i49CzrZdtYgNplUEfQctlcup0wUgbJLR97WEwEXetPDg9xDmUzEo
nlWQTYXc0HCAQtHNq2VVNh/nOzGnBjoiSAG9uBmcjSEQwLclJwcMf+YhyuI6XGwgIB6W9TDIBAoN
lJJX/s0Luax7owTAuPm2sb4f7pbaAnoqVgKDWsFkIuR4itZ/qHySppfyQrxTUFFtYc7bRTKfrlB0
R/A1UyjD9ZNiADan9N2IPgzX01DRCBc+wFxQIFyf8b6NuRlnif4Ye80p/6li9Pef5FLXzFjRkMlO
+s0lN5Tobgp1nNg7FQLWmOUxYnuAJ6uLm54tS3yH1L0KsHXs/tCEWIRPM24NUdEpOvTQ9XYHUipt
Gb7gz5ZU7NyDeqOc0Yd9lgeKaMSbV6kH27f4EGMPi4pSP3kdgbQ7YYWqeo84IibeKj1DYVEw8ZIq
q/84ebsoYrtAx8S1ma9nWXJVkDuD1E4+44u9MfovQpCPKpjuevFtvKFBxLhXKe/vvVZDP38ZgE33
ztLTT8LbLTZyKlbjPJ4jkwSaLUGGlAUrLZA0jvUc++qPNCecv3H4Y22EizRdD9X1Lm1ilOvmHr+E
xDBMydaulWKl3o64ZSMUrbxTQnxJzACXq3H8bhlbkS3/GLwLFP5BBZOdNqeQsAhlUMTjYw4lEd0X
7Lb648iyz+/B4BhPt84SBmK5NOYBIZECeZaA4J2rYYggE1Ymksd+BwfTSp/HMqnZAIq8EoYLdEZV
G3PSeLOaj8CRQF3Z1xJ03fjy6NkBf20rJS9CRSIFcS5IeVApRitvQhAsFJgFnXnY+Qnwi+rC9EXE
Fnt2rw458NoanmbVB6IiLmZX50IVYU6XZjs+12HAob8MHJbyotvyEkDM+v/LAtKIGSAd3YTvNRja
/MFxQ2IbmtcamZ9EpDRx7lWT1ZhgoeC1ZMU1qp/YE3+Xk1LqHxn3xtLm+l6I3bh7sToY6fGia14y
FZISM3qLX32/V7segnPiWwSdnqToD/v95uZGMwE/RuC0vDTq7HXHmBFuyZ0W9rSNB8iqY5gLkJcL
nWTSDaEN6EtH54z+I7VJa+CZMsQIP7fR+MSs83YG25w3fnFkvgKGPa9J25H7Zw/nqy7EtoDwg46y
91jE+I8goncj4fzr+0FIK+g253ww094V2De+b45ByhF+kMWuLM/UxlPxVbv3yi9QnOgY8JNWb6FT
U+Txui6GdRBfhmpvsPzqMF2DlhIxcgo2tAqWI1YwjJZUTtYuxtVFKqjnE/U4rLH04qcnnTAbZxCf
7lQWwmgEDIPrVvHd7F85dJhaUriG0spkcD9YpgWPG/tHkYPAXQO86gNHrwUXdwYRBW2wawyxgwYl
AsK5X34LqtiRc8Lx67wUgCUT/mB16JGsuBp2/mtV0ezVqJaaDkXCzL8hsfzn8Ma5whtSo2LbJryN
mPakd0d0OsZe05U1WuOiodHt2F7+2Y2rE4ZuNTG06Uah+w9FqKhZ9WnkR5Nl5UdmbQKfJHJqeabk
3PKWpK+DZFgp5Z1DcA6OT3FoA0+QAYXgmgrRBJ+3EFaWQ8hvUicSksBzIXRQIvYDjXrYXehsvpqS
YZHA1e3ECiILcfsecuby4n+Gp908XjuminZ1wMbbRjSEEcG/rsQM8ghxXbWNGw/mUXROD0uUer4I
hSlX2XM33mXzfgJi30vPIgfqtagakv7BheWZyM/PZEjUMSAysP1TGEfQKKMT6i/f4osCc1CBjhkm
6Qaj4A2ntVL1s5xJT2ESZg4H/v/TjgidiNnOPzbPgeAcjOL8Fm8Roq1jtyiZuJdocg+myGTAI0jG
/pAVrVgLaggV9ujNGdyog4j8mPgMnsxSmrukjlTM5KZ/2+ZolwgF/N0jihLYGR0Hy/FWzqTyfJAn
8Fx4mkLDQyTCcbwoBRuhK4oXpfkWkhLY3jZF6V9AH4XzQUbtQeURgSF9uvNrZUjdpp7ZvLlVXf+t
dRtkeN4co699aeHlwZImvY+EPAl8OevF/0E2TnJ6mvz3gampE71hTuPlOStBXf1ZZ+QAnnomOTw1
dJx78+Oz8y/7g+gWDwpa3xRJ+BeE8Hcy4CGBDwlrWPwGQ73NXg+1H6dmvPaBjRteUpopCnc3BP50
GpwGem0g4aCz2pcuUZoyamaZ4/6+pbzq7PxA2/WMVM/9eoBBdvxREVBXwiiolgwCDz30UhYCVdW7
xyo8t2cTK6zIBLegq3uJog+YSTcwJU4jfh459mcY/lJJuUDawRnFNcsEFKyH6v7kzNqoUfsbE9IO
kz4TpAzd8xT5X0xvEJTOZ8SwGIq3R+1lgygtulbz/lgNN8hYXDXU7fZxWcW/XbPteJ5BdRMOQGHM
/jcsDoDboJfg0lAGFmgJWaaxLKNkDvHBL8V0WD/zMumJkf3WfbYWUOU1W6Ai4hbr/UIJSvB3j9/g
4jpseWceP+PTnq5aS6hAcDt7gcda3QOGzO+1P78faJvlUNU1Q1IXxvNTiZsUaJ6aJB99lgNWgHxB
OOybziCqWTi82h1D+sR3b3UuAIV8n1FmECfrzkU9pveYpsvA0cncuMiyLhmGlQ4AnqIsxfKYfYu/
kU78KPdslybMWQTOFrutynvRdr7tx/EIhWgXDAQ89TvWsVdR0TOFyaA2lJscaX9dTrhphqi02n9F
P6duq7NHdp7I01oOiKwtgFGxDCuClUBQGvZwdG241jxej4mgzMtLlvuP5VaOoRIS8t0cq6W/kmy3
9aYtvcYA2j6UHPIN4ssHSOCO9eeP8v4jcQyADfPf78iiiuSF5lj0QK5cx+7t3yWDzCOgyKKJ/V3q
lX2GhJvpJo0I/S06SHYaYbc7LAfFdwv1JN6k3kuXwHZStxGJqxl/Q7WwvK1VAnIp07aNpcHoFM8P
79PR3ScKAh3y1wDOib/6r5/77PDfrpRE0BbKvFT6dLK3SVzfhrc/EMpksXD9++jmY+syJUqhCUv7
jurEDwr0oTygeJ5L/Xw1462QGSPrHirD/geerydqou4bmkDNvMaqTvN2sFmyxYbOFXU/XDnwaaOr
CBstf/kicsBNM5BIDAh218+ho2jBqokDLfE9/rf2fJ2xeERw/PZqOGe5RbtyPo0Fx0fxsRiLmNy+
2XldKLdi6g49kuSS1pCbHbpyN4uBuBbu8iI31U9GO+QKIqID+d9Nk6T3foIS1QVHS4uhQuTVxhdx
jCFzFPIK/V5B4IQFaMYFE8LhlzqEgw1FOcnhsDSV3D2R/zypV+VomJMX2seA783/Fw6ZZqd3mWk+
itRuIcg6gWjjwt53bxYveX9dDrvVM57eFsCeI+VcR4ksUh0tzJ/HeRV/PaDu0dOF24IrK3HhD8IU
Lx36EyQ5tT4ffQVwuQxSv+AHMJTUxL85EJ6dOeFgX+8swXlMA4bKzKebmiZSWG58mBdNWjENuu/z
AvPns9fp57W04pwuMFKYjHAFS5vDwBUeAf6gdbRj3q/VevhZg3EXdYklO/DAoQIuSUXMJ5D3sNs6
xHnE2ZyRizZ2znpQ5JTJtfu/AlXbhWhcWUHBEpa71ts237ee7OGbh7JxPVvmxgGrABFJff31d2ZQ
Mp8PXhg93UM6Bads/cmsuOY7DI1WoZnR7S64tdxNDfYZI8vMIZb/M5XdCrMRvs5QAvNYaOyBM4ae
BDJ7ZHvdikQDiU7J7zclr+uukAorNuQS9UQ+jsk0TcsIVgp6tUnwqb8KsXkSgkzCNvcMvdkOsAzC
/AOWrveyeyBTQP/dslIfh2iogqiPkjmNjwRUXGsCIRbDkl/JdBlnMHgw2YqpvRDlYOTcDBFVC7ZZ
9UN68K1WzteZzW64tgGL6KiwhIAER2vbpYRry04Aa4s8ct3c6CcF0JGvDnAJ3qtnehaNHq83uzvO
1fRxQh6tCRB2XOV/uHVV+tOVbYcZtFW+8p4LGcWsEkNEXPUSlF02XS0sDX4NIXXFiJzTclWSbi3o
NnAjYpuV93EDdL3HWrf+3JnCB/TMtaDQNT7tIJVwGt6QxEbD1NJ0CyViqP7Zra69LTvv5ocqqSMG
1jG/wrFq/a5aPnAp0eOXQ8aAIRSugoxYxgxfZeUQfsYV1Fi4UmH0ch7BjwO3Hp/F4hvDpOW9Kw8Q
jHj6T/cciv85YWS3JSXvGWKJ1pzyBxWSHyQe2mgZZHX8rT5dTAIEiwWJJcquneat4xMAKjwWvyNY
ZMNe/q+4g0t3fbCeV8tDSzpSFD79uhO3C4Yin4EInttNlQFz8NLWvv7vFOky8sKqGemAtlWUlFxQ
uii9YauiBgomLCEfNtxecl2NPNwkydpwws4zNl9S5vpG6ZUuPW2hGIuZ830gNobOLp0W6Ql14jiM
GvjNwPWQxpJM3hocNiNQbyATOIBY8t4J2MFW3fQxDFfl05ObvrKsAtI8jaosayKZRUeEawDUXwt3
3Hs7cCdVlcpD5AfRWixcDqWKkrfFFDWIxfKGfITmMbzwe0SVItjdH0CaSb/pmZb+W0v/5T/lBf/f
SP+1tS+HeMeOuFApeP+O15DEX+MsnAijYZx07IRatOtoiOhJdztuo/RRKs3xyp9Caz6ZUidVARpV
EjRSxv25O6PBjcm7i3YXSerl1YDQZaBH3LJ49sWb+z7kBTd5OuNgXCeYKuELkicZiYNR0ZIJORjS
TVzfpH/REBtiQt5E5mYG70O5k6NpdAFkEyQl2qfq0UOUKmynnGPo2qEpCOKNMu94eFrgM87ZiiJi
Q+RJXX1+A5nxAx1cdofG33zZpXw4KTFwIw4Sxsx3OrQ0daltfX1MwSCwMSkWTUEt3N7/v6p+yBKf
VGOk+5im9ZbFMGxW5/dfXZNgbvwnkw4yaXbGdPFtbdFf4LfelaiFPWFgoj1XaImr8XJEC7QkpX+X
Mf1DS+1+Hi+H4RQiqGUrZbDRr8eF7/Kyv60eBF2tTZ2yCvmsl8l/mjOqGKMhswwHc3SBUg2Bq5Ir
tFrHY9RyxUIACamw6IA2zc8cA7T443i5jaNH0SI3Rg9BDlkjDTkbjA1qTDqgNqqTX2ymaJM5EAXI
/f7Y4nPEFqtp24Ru172fyhNuBxnVJV0rh8u9kT8zgKCwshvDtP7tIBZmaV/oT6hDnQdnGQZCOvuX
WsNAZ6TdJE+Q7MDgYUtlPBpSVE5YFRWHb4DmxnhbWLMTHQiIDzPR6qsn0+7FgdokfLkM1BfTMv3x
FHdmiMHpMDvR4xQJeQvvx5Q1TtpCUnOYeqN7+JgI88wLcwk6kImZuGXQ4p/RmBPfXOr1Puoz6vwa
6s6zkNT7sRIpr7J8LwU0BDvrpNuHDSGll38UkMiCx4sZ8eqsWxTpL+ZOnjLiub2+VOh4MvwGS+mY
6aIcWKH0BnVUM92Gyo/3ts3PFmKtO8t8pX5FeX7T23JE66T0nt2IBdjBLKQop/WM16WC2+AzJ8mW
csTu3i91bBc58jC2INtnhucmWeMtU7Upb7ZCUziZu+tcy2FG0P4cRyWpApkzLpA7VQHOB9U83z8t
4y/xIqk6DDY6JmFBJEw4fiHmpzfot3+pIjJaN4kEKbpcUxlYFVpsH032vmNKPzuEzD1YhqWgtm1q
4t5RM748xBb6xEWbwTI6Z5szFR1E0+hRNWrQuStiDP7aQqJIaBSq1oMC1len9b0o4RdKQqDfiDAw
DQdXUQWz8eCrNE0DUJPE5W9BlWIDCNY4fufseY0kova24XoLl2UMvrnips1eD/UPmDiz5uR82ipT
Gy1x5/Rsmu2DJ5EWYdTNpo6Y7uhunPpXuTl5vkdfem0fB71rW+S2qdDsixTnh0MTdPahQX5ajWvT
Gk84fBsDrijDsAZ8KjRLQfQRUi3RmTS1uOQEYXijP8F4qYo3mn2mRXUj5iyBdxJsqlt6TKZeR9su
Li/voANdRGkcbr1DVNv3dS7l+Fq85/pcDLhu7wbD+ZrXGFHNGOVN/5VnuSPA7o3nmNLVyp256dCS
m+tVnwQBAsbFZQrSJ1xYLKX46xpB1ez846+hJkPtnNkCTMFIw6l4dQ1jt0cn8+01Sbfk8je2RmhZ
L7OyzMngomgESL/rwNEtAkVR3yBDLAqSo8koEjGp1QrBFqFPSWqL+k4IYHIwISObLrFLIYYUrBRE
c0Hr6sPr+v4bWbKt7Fp3uTaOI0Sh919gesXaRhfgSgXVUvudQ3zGdhOKKXoLvq3mCfXVHu3FKnTE
/1/8nThUQXqt5EZ7osic8uKKP7IggzkDitucApHE/Baf2BW01xQ9ftm+LDnxUHNGc7qSHC7gbznN
ld0SlPbYFTZvBiApFJe7QUoZNKQIdsmSqCNW+EZBZKlJVIoGujADMHk4HdgC1RVM7aer2oTeKwtv
8k0C1UQFczsKx5CbeXLPTF+d6XlM+ODcMjTsIw+/otDDuZPeNIrDFTV/zGksZMMs+y2XMp7GCmjh
PAdEeMnEF1YlRdtfEW+tOKKYBlm2hQ098w1C5Ph9FcpZkxCe9cZKscqxlrpKbFJ+pGi9i4uHXhxK
61EfvnhP3cokWBFTpZgPC2Js6OA05TmWbXUsEYsBPO5uQaQ4dQOh+DFxpfeQs5bKZgh/9ksZthO7
geXydSHccLPyonA0F2wiodVmsLZixiACiGpfUzr2PMV5Jb6U/3dQ6/KVyDytg05d+ppp/e9gFfNY
/D684PhVQZ1GH/Vjfniq0NnHnnK3Rt4p4op4oy5DdAzobE+vGiDDVbn3VWfywfL0u8RQirrFrVko
liiZhCYJjNfUHcAGepqYh5sAocUbRzu+lTxvPYdrzbq71sEMFJJJIK5WCotbRDnKFYCo4C3wMwQH
9BWcgZoDUKfq47efwfDykduIUm1lUwAktjDVIPIX3FbxOuHIYzXY1UvBOfTk0oTs0mNg4Fdkomni
8o7Q8pCzU8XHTtEf3ztRADz3G5vU6f5W8d8022mTVRYUpLjCKderoQ84VrgZzwCCpfVSh5J2716+
fhEOnFKw675ZAUwg7hbXmjAdilUxYTQGjskj6lJb39iRez7lYMSesQKh5Y4WSKK+16wsEoYCdjAQ
aJ0s3fZvF0Zs38yx9QYriR0xTFP1J3bDZktbI68Mi+bYs1R1oqu00j0tUrIw3nDAlbYhqyth2oql
qQ8RrJqGTNQILGRId4fAktcplgGpc1B9SwPcDt4BfAg+WeNie5V3ctHd5tBN2il7eJvjM3mxD+lD
kWp59p1N65J6S+IQAtg3CbTPXfYNvtzcfC3mhjd9sPIzMU/SA2Ed2RSG2D1Su2gxr0MMoxNh6jSv
me2/BV6v6q9gyNAZR70rGNI6GKaK+B07RL43zmiKNCHjeUNoKUvN7fPkesnya9bTo6JcRjpVrIZe
lo5hSwfN03GZ/H0gF45JmjqLTI/aHHUKp6lFpdE1UE2FYNYxLCfVPFYusAE4b2UIh9H+940LO+Tv
k01UBs9Kc6v9+zpMrmtLf6nGLgEWA0bZfD3XRBhVUhXCNIkWStXCx/kQY5KxMqtSX+RmgaBrykNT
n0gzEqnSgILJ3TWpAZirtNaVyzPjVtQ2gF9hKJLBjpYgXWacPYnVszrV64ia4SU2Wt2XYKsGh+Rw
BukH46LF+zMe3z2IH+ismTJtFxjeANdBFQ2w/+ZnXxQf8wsQUpMyko11NoXkintrRffTpfj/Y/zJ
S02ftB+gsqpVi2HUWi/AzO8BFWTpHeWur/pjx39Jcs2epGDynGpbMWDSWYgvqvK8QA8hlOFgPS8j
0sl5rAsc481b2pRs0bxDyKhf7yGJBWuaXZEExNn+Ze01FmIIkxRMSTjjYgl1lA4jUxCAgmni7zjq
819TshYf/bpRgJKCSaMvIg169FJiitABYvmncitrhMX4721yo/mwVuLsgMGA9o32J1pfXqGtjVmQ
1X01y8hSQQrIrMsMN2gcRVdubh1elHfuC4jmN/Z+NJiryrXagQtIDu7hgYHFduEWxlgYi++DR1QT
j027uk6yyLhmyAyMRb3kWhk1427sSzTBcTmcm1/leL4mB1/YB9+X8ZD/q+UPJyBUV2Mg0zRTRDjw
cmHeLNzsGgfNT7EHfRR2G8Lxtu22eUFdzUcYW7Reun516JjPq7qwNSdMb9keAnjvh3wJMYk3VbO3
O96jtNMW0r0YVKUIb1anO7UxS03rCs3kfEUwvIClEO5OeWN4zhyNqTGdYqKgxZkm9KRHUnjsetQl
gOZOLBC4QvY2MjJOwG7uaqK47Lw+6d0G/nB7Wte9moQZB5B1ERnwSh8t11nsrYzRkqScUbbdLFNE
Bz8BlOhLmZ/aUXk6zUMFN1lAI9yiELRKk+y89QNF3btk85irpBzhl0M0qCAetOKKkYHynOWVDVgn
RS6DYZ/4SZGWkX2P2s+kOXWbCuQbwCYlzLSfc6QLpTb+vFOs8Bsq3wuFo9mV9tbxmB/447/zoCIV
m5IbiMYbG9/WtTysgAzCTYhKew3ppZl5ppRx75A6njLi7MgTXeDRWaYjIAkudYDUA93QRmysB+rw
JeJ7PLTBWK6VWmSGbbIOP612c602b4oxr/X9tF1hXDAI4AOUDQRrs1dCH/EFoJl5jvFZugboD19W
bONCk6MQdfSMaJw3zCIw9tVDk/88cP76UxmVNY97YMmoumKSPN/zX6g6RKjplrDZCZpbIhW9Evl0
tLmpC08HiJRyqbyOk1mCy95wRwvz9CmWrfRqrZkKJkE4BdBNircAO36jwhIiJgiUDAV7sGLSpJoH
0DdCDiJZAEcNjPCOBKFEu6NGPkxRWLata9WOMemL7mc/90xE3LaoiZ8cOoq19HlfMPUgiEbex4AB
Eih4KqlOB9q+RH2bwH30O5PzHrZBTH9IF1buIJ4lHSm1V78YpSrU9bY9avVwlca1fIsaDwFMnvoI
RHUlT3jxs+DG8S62MPoTRULTcZxsXG4rvebXPFOsqIizQuF4tEOcT8++xP92Dz4ZiD+t0gwkxXcA
Bi6EUNB0sBlZB5l8EAzpktAM+1ni8B+dyK5SSQ9gxnG4/lBQzmrJSw1A2IuY1WSg+UMwlMVZT4rb
pQtYRU5ZExgZtPDGm+m6z4n1IqTVtlZ7b4/Nvmyp5rqvBRYTTTYIo7NqZraFDk8YG7NmrWoIsq3l
EbqFxoNh7TndqFCjnV6D2rOupTMEK3c54IsfMR+qqByplJKJdJjYy+Nptdm0qSOUBH286u5LZHHv
xEplr5JVdHHqIJHxNxCUOkixvKu1MW719s8sg1cWalg2d3Da3IQuAQUBPy8LZGs5UoV1t0S78XWM
2vson156edFzZT/LOqXx0aFUGA4hhcJicqzAf7FWsPE7/1SV1xCvY6zfkeP9ehPqNd4EPv8sIMXv
ImmeDIb0r/MCSaxGe0X8FSsyA7eKofIe6aib4d8vr4a5AFWLRsQhJFC7V1hHf/2N/J4MtAjVe+B2
ASMlgLJdaHwQGETq7ktWQCTX++nJRYNCKBVydW9kOk7uTIsqwrAWYRVs/Ppk19fPlmYp6+AaK13A
kwt6YN3oCVVwfElg7YCK8nQQoPJyrEXbpypNnkmEMge7Ag1xTJYqtncVCgw5BjNqggzRy4WNgZ+I
4SZb6sA2UWxzmPqAG4CM+TYZmp3E4OsJcEZQUATOy1v5uwqG7wcXVwJCQjUlhZhtT6R9QJmThgVp
tU61chcAQRQ++5KqzKImDBz33RqgD+1msMpTjJY3vPOcdJEs3wwyaxASNSHMAfpU4W5f4ejREMDO
w5+58qPfLNHHmGrfVpD/Kens3FR2+whFVSm2ybzmo+Izt9zRsimTWi7vM+uGvUJJEVPCnL2rfims
6xk4NvscsZSZKVOV3LlvD9Hf5Ky3M6pm3/zvUSFKRJDgI6rFsbQRGBwIC24YRsNFdlX1Lf2brAeW
hphmmEVm2vBBWKrcNEd+GOcelZI2AuyG3y/VCctMAfAiKrACDNI9Rm69kag4tpWPDBLPJA1ANeDs
RHJIIxbhc3xKu8Ndo21hO30UWk2bwjPYewsgn3xJQUMMbj5XlEI5nrqyEqXrO/2MDqf1BbsedrFG
ZWUC3erhqqgMBizXT3UsrZKMJaKTc6GXnDeyPmME6R+Dbhmxk5AvQvAalBuhJ1f3PPtcCridw8Mf
qPPgmdtY4WVyMOMrVnO6PKj/sv8FUhcZMeZKK9zO8JLTxkMvjhEVN4TP6Ay3tAOk1RdM3jtZ7C49
VGDC6E5rfkB9k4yQ45y63ldHM53lprn7NV+LrxZmZ6LKZGIBXCYK3P+PRCPSE+IDZ0pySW9vD1wg
TVQjyvSa4S0cT4/5mPth5xA2ytMP/Ho0TJOljZ2hO2yKnRWy3XlvoTkLgnLuWWOCIdMUM4V3Mw7Q
DWxiHh4JcFha5fC93orahMxAjlPoGbNA/GOvRvRMduuIHAH/8iwPfZNaJ/A2k5IVsonC/25VYNuS
E1ljPHGUPvKk7SP8M3WB67HtdeX/+YbvznRinj0dtQMO5TcYzpHmvD+3VONt/nOcXh5BjLoQA9/w
0a4MoGVjccg7RMcBpHyimsiz/8mRWqseRTgiEPW8FDg4YC5M2v1tWVOWFYE/NFB75KpwEOwsq9JM
5jlyfcwyO/Z/I3D0EimXvGO4VEZbroQ7qJJ3PWCp1kaWt/hjVM6BI5FDV30US6plfp5uZ5PEfA7P
PGPb57+k/ZI/0LZnyyG3y281EVyDaERENv4DW/eb34QtWPj9PWtmCKdhLJi+ZAOM27ef+k0+hmBU
tbuX+rpE16kuFJepbTnmlQxrZJpjxjB5iX/VTD9jlVZncgAm8s4zB8opnW6HpaJOGXw9gOlkPGvD
0g1SW+ovO8wBJqZ2WJX3HLMRgi6hiVdFkyOdjgPfv6R00gwqHWs3IjUp3RxLu9ioHgaZU2Woskz5
yMq3AuGJ4+wz42vb8Mw8PYNj+tIhhWbCTgxOCBTcEitPnBSB9pc2eQNPab6N+/bWAQMknjpnxvOE
OF4buFuIVICPieqUNMMzPswoYEff2CH2iBX/9UCEn5Vd1X7gZUqdtKn1yStJP9Be0mtl9XPOx1zU
a5//eY26FUw7/5NqZA0yeUDxNSLUTdLkZFc2K5m56DlxXyZhtvGJ1AlRsCrc6+fgqK4+M0KfenRy
PtXTPLO8MMUddgwcq4hVHUbaaQw+ZtYMmg/0QIgvTRQKnI9ze04hNebi6I/hdsHB6E4wrFnglbp8
lTW9ZB702RIXS9dzpPKD1EtJBHEC7djBdDiz+0oInTWfoPSxEq/1TexZbOySJqUve9ci4iRaWkpk
tZry9UOBhq8S6DJ6KXsRp6Q4wjhw5P5KtqSJmN1AdseaFH43z1eF/zAc4ztKg1unHSgSQOLvDsoP
STJ+ndDUiThIj2DL3/049qfXTeekHqaJLEhJGLt7/dShuzvw6F1ECqHt2Hk64yhq/QpBgW69aqNW
De7wiQkNI7IMk+EImuSQ+6WAsoUErvRfeYP7N3ZgGMkKiDYsGIhhUehLEk9B2nDjCyZecA6928eg
aZMVPlXpSCDiSfn72vU8jE/TRTXfoJMeZippxJKBnmeRkRUhzcR1JSk+LrFtkrxZpjecYLPZzPve
mTv5236Yp8e52y0158ItC9HQvywjPZVVDI9M8DuhRwxe0lg861bJcnBAuYlVcbGUr4HDUqRqE6QX
+dV7Gfvp6GjNF651xUwDrzDR1RG1wU9DfdKLJsIUM3aqUUbno1wPWJrJaK7Z68NYrOg8NV6sZusn
yiYDpwq/ZrjTc/XJxoqG7bv3BIR72albUcoUaFVGQUU+Lx3N87UlTG58/X+CRTGQYVSavvvrzfNz
gqq8Lf+ONCFiIj/EaHOeinYX84Ku6T1STQwm3Ow0WT/IvfVwhB+Y4eC+SrEwFGUtSpr2+JmTdKHj
LRn5LL4C4OF2jFNCi8HpztMtuutXuvxLh0Jt/bjP6xWLd3f/xxxyqIEVVld2rHYS9zXTcXT6rmg2
BRtEUjDCEaDzU5qnOGfJkpBL6OxofPVx7Lm8w7Iexyq5tLncXfJDr0pPRpi/JqV85/vHEGUkZc57
7CcmlYa6bP2nB3qGtyV5YTwA+vofxPLdCKHvmjMr0PBlIwy7N3NL1unNnQLeYMuYetzohma2vugn
e+MguEyR5bcv11ppwIji5oaf0eFv24mkdEYytrr7WOCb2aDDV6avW1VuqCPNS3umTfilSrBqRalG
cQeCUfOYBFt7/vUrGBm21H+4C3RXo0ZsNYkQpMN8OiRg1p/Ja+MgcpIZKxV+F938PFPwslrQViqf
rCKCRUtlZKAp53Dg+7vEgN9THKPyP/RHmN+7Xz2PZGxwUT4j7EIpQFYDoZNill2PBl9Qrskby+je
iSW3Rlu0/TwKWJbXWeHIUY8LD9Kbyme6Be/tggptsk1+lzk85NnPiQW0pJ8J9cxYN2+LxutnE/+Z
1maEeyRXbnxfm6W/aMRT14RJ4Kxr/HjwJfn2rVVsdD/EIm3XZ2nxJAR7abemyPz9X82szKJbmPPF
w4VUkqGFUexd3SHBxrOXm1FrPxsqYVECek41Sww4sBx9T+rPpNH33ldl5VxkWTPrIixJ5Z9Qo3fx
JVAPZFKfW1q2D2nUecH40uYthTMOSZL5BGKurb7/9vgdEkye7Ni9BpcBQfzdKk/SKUgFA43abgAJ
ZKi0lk1pE5cbiT9Ja1Vn1ykukhHeB3P6df/1XRBton+S0MHo8YGURWtrqjEBZi045V+ckGBdUh8q
45zwzwEkf18qgxV2e6b7YjrI82dAeI7jqJocv7KZuOFo4Fp6cpJFxFD+FQdlxApgVuWITGqUVbY+
tOAGvnCugbJsevxecBEFGfTL62cO3qnbEPn4uJvzjZenLSDrlkswJ/vahz7rgCTeg4/ZB87utaxZ
G5xu59OfFYfYoOC7+KzkH+JTcD0OtXPJ3z3GicR5KMV1tXey9E9Fa1MmuRT+x9saZ0WaA+d09xFi
mQbQIU1X+Ucfoc33NGZ7vKSoCzZTUZfInNQC/JgK2oTWQAV5wvgT8TzBxUUUDA8hTquD81KCeDaq
EHtLnZdGmxCOv1y0vUtGVnlU1v6X3XwMM7t6kGdOXs2nY3RxFatA3ABViyEkLHUTBzM5c4NIzEAJ
ins4BKjJDRkiMjSWmFKnMUCrhLEarbyTJx4qKRomL9zMKLsQhpZoLomj+D/tAdKPvdPjKK09me7h
YmpBJKpMT8ZStJml0oUhIniUHaeSI0gW33eyE/8cOAW/GX4n7uL6CpqB1/G40nqA3HNFwsJq92sz
5wvDk6hF3iASJFOYcL7bEys+7Z6P2MNp/f6nY3wSJcu0lLBfNLBH+LN7SO6ayGFHKtn2NlNGfpzX
tkXQixwpTorxExnx5BMSCToM/bbRdXmhcUYza5NAhgySGQWJVyP1z2F0rNqmuy9ry2oxsDN9MseY
lJf3LJoKht+81k8+a11seMVItB++2AP8/9+s5qO42euQk+AmIOooMLZnh3awqXRWV8pDRt8KpQIX
ZSvdaAwxPZBnsl3IWW3VH4btFYKXnjvE95apWtLiucuzVtoprtuADCdcofPXy55+kZnPfdYMPza8
XKK1hm9TuxRuDALwPajNAr95NyWtbWCLEGPCqqgPTksTdRtYD7VW/OBILGSTvEwEe/4gCQOCBpAc
GYbSCQQfMDRdZl9rTLcb5OxZOzyuyak906+xW4IGS58g03FdmOr5dwNMNhivspUQd2OKXWfR+we2
sliH8Wzwpg8vZgX/wsurPhaWByqnSVvzJwWfjGegVHJRZs501/eEByVLRjnO
`protect end_protected
