`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lli4WPcwyX02+Q1jv7oZnAubULvwsfbKSCv5DidMvyhpoDhfOp8jfvOPYU0NGpIuuURfOmuQkFhk
NGv+/UCBQw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
g5OofTPIBCB8noKS3hAUwmUrgwJ/9D15JuT6C6b9knLViEzE1tU9OEng/YwbBFySPIM+PT04jhVz
G4seOqCZlqkfAfVsBpzPXXSvginm2kIwqZ2/okA63RHYKZ//k9Qg+wjClHVlINHcaChUXI9pxKT7
j8oPAYFQ1Mrv3lgBaP4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oeGcSYSnFLfarXqLs7ewfhQv5rZIg6jAhjdk8MnfaxvbaDAU+UYovEsK2d1HXTdwNRK8UijiEOTd
8IqzBoIq3ltK45i/Ph59ikfbfVmgbRo+709fuq6b5M6oViRVDFgnd6viB+t+V3mNPdbVMThaiF7F
QhRsPVeC+m/iw5icBwCgBWHcyODTUORFzjjKLdx0Ncc97+CAKXbgQryBuvtinE4RTeuiwxXmawPP
Vd4/XSBaYIXJnqBwWR2dWl7dISC2AF/Spvz6+aFeBY3iZF1Q8ZdY3mRKEz1nViaE5ov5EQRjZOcg
Hee0zMsRnlty4x+AAqk/8jtfCn+xgd9d8i8D1A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Oa+XcrT9B5gYB6B3e6UDtBkut3ODhSN6LLpLHQpPIU+Fdwyhspto0NDXaPfx6k5xR+cbJ85of/c4
2t9E5Bc1HDHqsIvBZXBIHP9Murrt5oVCbP7W8aLU1bSrqiMlN5VwTyry1nUf6uQWIxgmatnYoN1K
AFIExMk9HNg6a9i1d1k=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
soB5JS6OY7qPSyrbICYwfBPR85NiBnycjeWdv9Sb7uc2KwVzOJpqsbhsYb1F46Wk5LoElkcsPog2
3wVYKetulbSyz6aWj/LtvoKDdJRqErLpGxBQVBo/zlmy2I7gnD7AGh39ZMwN0mhna4cjWI+Mlsq4
fweJW26Z0ZJpAVzs4N97ndahQq5Bc8HKTqGlv7RgcnYwLwm61i3+gDmJV03BUkKFV548QSkOf5er
pQka3GEIIHcwCyFJQdkUiAXP7UB/DfywrUZf8i/vNmjz4bgjKsMznMgdNii3bXKXtTJGmMxDWo4s
OHp9s5H0wRLA9l3A7fN3L36IPs8jxLl3SYMJJQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25984)
`protect data_block
jweNSrT+RhL+1BEGQVRpk2QTJpdTgnhDxvEMv8UCBtnzSJNkCqmPyzCUJKBEOvgfZ3OjcrvzthCU
yh7agcHwr6Gmyb1FEk3FITDMqDgKcv/IhpMeEiPIZDzRD6/XpWUzpwWS8L1/56rpSM6BSeDv44pg
PNT39bm+2jbZByyxiX0QHHv3Ewv2CQ04xLfdxOGFuJJV1xNKenKghoIGmpPkKeiPSua0FTgiYWZ3
LNLDlxAdZWDDvodpV5thckw0qgq+XOWt6fB3YOJKNIPQ902wDGN88dGSEfpeD6GkiYO1lMDSVJ4G
yswwMTGmvFAGUoQaU3z7QEE4MioUyVs9asTeOg5C3ZfjTmRGWoKT+dpoHEsbe6a0JPodC0paS/Dj
SDbMQPWyrjJHIARLuVE+dbTrS5Y9S/ijBQFeWODkVY1AEE3VzshIhaLiWVNmLqjExs8Z4PIT/zEd
BP1zvh+ne/9aRfSJqKhQO6ntiwVePzez9jIWtlpVjGOaQOjXMGqLFHO9xO0KS/rvbfTCpnKz81YH
XABLk4J1p6o9LAZJJsbb1gSgjtooUREyjJriSZjMj0BZeX1vCRNJMR/ROMUCmdr87KxmUlvC77HE
uk0ljinHamYJWX+grmHI3PPedNXBb6tkjf6oG6M2+2larvfvirzpWrUmBMRDEoaV98uy/2cBNng4
9d3G32OswjGpHqPc+rb9wC1sXX0eZ0FWFfxA7XE+dpRqQKNJX4xX5syDgEn7RLYYmEL5ia3M4vVK
u5eKJ4Wtkd/Tyd94RLaA2fYdHEpZT1Zc1icY5knWfoOUYwUGU6vBE1UcoDe2f25PvGH1rJXs3hyb
lsjcJbuVDE007FY2AysKSccHMI2+w1Yiuh3nimT0W67Yblb0/ZYVGCQzuhFl+3w1SRe6RqCI+trZ
2lHestY+R+2+OmtjkZAyHSzoWW8mLOFp5Ixfo/KG3xz6bq3MGd/9ga2kDQZRGPYJHdRSgOHAimVB
QnWTw8J3R1KvTA/WAhckXVtwvhVxu/FO/kLVdoVwHjtkPXAhANZZfv5QjFDE+WaicnKz/QQlCiNe
2et7V+TjhRa/NpwQHwSiqEAvjQqXivai3aW/S+1L5fJCvP8ZuPY4W7ihWfQuKy8CpMq4LV/c7lA5
8em6/9cTTAnDMjMaLrIkDi+mYEnHzdGcf1bNwGbbXtLQzn9N0pHtkVBIgfgSeNUpduR1XR8yZzEe
A/CzCfFTTngsTYIfmMo7jx4svV4bW+gyGvJc48+02aNVVh5e0MUxnRiXIVVg54k+Khqfmn/PlYBU
cpSI0GfKM+LQRfisSUnrUOTCVZvSutOR4BQkCYDghQJ3+L2NPCFOIJMRxSM3KKV/sSJOQvYi/10k
Z1RLI14XRI2CNtSICFr04liPxUe8VBjbh917LkWsZSlK1AA+jNI5qHIv2ZCMQcHxRnFJEXxplLRb
O2wwZxRLLL0umWVFx4hCNVetvaYH1irfU+4ZGpzPgW9sbVWKVZooMYSxgRvJD3K+MfnKJK6icIYB
Cp1HaYE/F83iihfVmfbkrfLiDtJ+9nZfToMN24rLKYOcIjhGJak4YZNPW9olBOdCXuXTxaZubbNe
v6UPzLSsh5UC7yiFyZRae6J1eNjrt2j8CoPXG2av9XaNwolMj98CWN2rji/EQ6IfnbiEKLvycBbP
4NDQWLGIZtDMKbxEHiMcXxyLZNRHzrTNpPTI95AsG47czzdB0O3WR3zaWzr9lYwvzGYDENJjAiKT
7dIQr/dKBkCqtwgkcBdZIDjDgYiMC6O4SdH4fgPgRV5ZVT6pcPNgnqNicY97n0raXCX2+pR0jdyw
b/4Ttr0HY9+8OL2rSN30F9YBa3VpPZrGHOo9vTDA08pB/mkG+P7VABDEGQWdBFqITiG3vUqUox00
Vre3lZQmPwOcplsBSfTSoM05xiF2BG4BL71cRDE/aBqINY/eTB/k7G6KIRZpeMlPeILC73PWn8Fk
vZTT9p7SRNlH6osLCTTi6+1lObsI6i7RsgbwPzERwoR8QAfh+wWFKwCiXPt4VZv9VAUa0fKCVtK3
3hgIXHrc+jeK2CZrsV9VD04L9HJEgj/m8v/ypIGo3ViDsCki3qWTs2rURs+5of711wPK9aGxnkbg
Su5swMnfwY3N03NvJlkQQkACVPVo0yzn8GM4seGdCtB/HRk2kFAwAYQrHJqk3v27lkrwl0Agb/dy
dgdxxGLnPWmOK9FfNYI/ny2hLVWltZobf1Fsh36YVDGm/PS35DN6Kdn2zzifYFMv+hDqwjdBwkm0
Dis4SZ97q8FqWs4WPdqSjhLGyz9CegKEWhsaDJ9T7wySbIOJQ8/onQM+Cq30c2sMB57BVIw+jBYC
6oFlG08auELfko27V5jyFu6x0i0KJqx1OdohMjirIHbklLASnmQOWBFNdbR2EkCb+qA+zi7zbloq
MPwr7SoR6+C86FEm9n0v3ykh4oCPWVcLnE9/YAzBx3mULtySaJF3wsU/dStfB/wW5K5IkAtx3i1Y
eYChHigVP3EEvRDSiAZBh0sa7dRMV1KHqOL2OZNa0H4/Arx4TOfrlVbfXhosSHQqQwvr+lAoOnxw
4MCDi/fsb2PONBMb22H9Aa2I71IHEZw3yRsS7YBxesRuBSBiaYiZM5FfGJSuQghjWGTRxGou7ODB
8Fd6wWT3PK5pIW1qgyc+7RmEGmlFbZXGX7lW0nTSdFZ+JSNOr3zcoyFuJgH/gKACTj6hlAm0NVhB
Q2vKw3UYxVueTt1g860n1kN4A8uZ7W3ZWvXShZ3cQZ9evlLynEqafUQb9id7e0bsH7eDA2EmvpZP
axER/V8XGk20relBvalRLwcZtUXFqBtdqWbQkJlGcY1wYZdgN4wwETmv703U2IGMecz3yYvhsQUb
GsyyGvRFdj1/08rWXdSgHBKiLAvbzeGqIukoVQNasRYUA9eiB8YZ8EBV+mTe/fyHdnept3mXOJNW
+fz2pVQPYMElf4djEHhL3yoAPwl/DsvGGVJSXywoNQfTqQ89KVtuM7FMJwKjz4xE7ptMlW1kp7Nj
5JmoN/fNLSQVjfrbSXT50fNuD1wVylXrk20qPme0hwXa0IvnDGiPgnZ+Si3plLveUrd4zW0skKM+
slgCffR2tusW+fdD9MQQLpk3TNEUVdiS/q+y8BOT1vjl5INpGXxkRst1xHYDEB16M7LutSEtxiui
0XnwMYeYuf9PMKMY88bOLl0QyE56RpFyglwHlvt4EzElhS4hc0SoSoZgS8MdK/iU/AOCs3SJfC4y
ZzEe6R/yYA5gEACJvHmjw9vInmnSgH5c2Ldm9es65P9xDipUgUbs3/qyk9WDIFzZnLIEv6j1mwW1
0JbY8FDs8H3OrnYf6YNhxZ+3uQJbuUCaJV+Ef1EE0BKNp9NhxNbLeNxGXZg0K/9xgIzgSi8MTXaL
fKoYlGsUlG08boo3HUxWyYlvQC17MWeiz0bHEAq67Zi42AdbdMLo3BanJEQhkaE1RzWMbkLGwq2A
oflr3r3+CO5BmMdeIZdyG6/dijvZM/yGnJ5GY8rxlLCrG4lARITR/uNyeq4rI2dlRjqUNUrpxaJ5
50QFQE/2E4NBQtF4mbuarOHXVsSTVZLuMJNXeuQoyBye6stZaAnW4KAZwDbG3KCh1lvdlDAJwFMg
3U1cL5nhGvEtCPJttqXL5r0hCGyaTmDg/mP5xQbkqJRYMPM2kR97t4j8DC/EDB3gfMK4Z6WwbQiV
7WXBKdtvfyU4gfFty9T1+fFAhEKrGTsc1+Fxrm6E6cP6Tuh2vg7G4q9el4MWUJlx/rIlanmxC0jO
nIEB7kJRKlIUL4cM0j5NTwirKdxY2nPx14L0/Bl3+X/Hbdu1UBLW9FLVGaK3rO6XoAEDB9ZBNcWc
aFUDBp/t/aFkbfcdBQeSLD9F8H2W4Y00kTLTbcXwo8SOiAK2nlvrIR2M/4r1RtvKvgaZoJDqFsgf
loQX2y1KYAlWRh2eBj6Oh8Otc62aOu/Xi5WTPR5kpKZO+6OazSPkvzoqv+melzxWNmTR4N6Bm81/
K6R8Qv/8E6ZDVz420VRhH1w4bzUbTPodcwO1gtux76Oz2i+zkzKnFjpV18JiD9khz9MfVZnIX+gz
K7U5ZtKik67unVWqd05JzpGyBVZIFejtVxSE+YwwaM1vxiBU4SBEkOiSNwfDI2OFvDnPT0/KqOq6
Nr6EeszUr4n81xds2woRool+fth4M5r6L3UNzCNu+oX5vOq3PUiBMQq+N4coORXmqRkL9fV9skki
VZLpkTYjVgGSF9yIQH0pMYGIC7aJdDdjfq5YTb0APM9mSabTTWr1ZhY3TgLgyOdPwudTlt7sTGmA
HD659lnnEdSYf371syVBEXjyjqwnl0R1lbiYRxLol4704wkJ7j+LWcAzLLb7vbv0QbGUQPWWi5V1
N0UMQmR6YZm8NnZxlwqgU8NDfcg4t0+V5wd7m0PQN9L9IOV5N/cbwBt+SOGmRORt1alQy+lbbt+A
ANv01FipoDtXv6VwPu6B7D5GxURvkd/hVnQqKrLI8gmAHRsAQ544eS38rJ6YidRVQ0td8szQNK+j
jiUkPngUOIWTPLqxQJ84aH9PqQ06MTqpWKZnL13I33SiFeA/lYjGjf28sDArvHkc9MRuamzWgCpx
QuabfWA6/+dv5XtamteNidgjrAw7AUHHh0tIolDHHVPrfsOKNxq5H+d+cwxv0h7i7IDWgbFqhSwJ
VuYDCCl0U2APgWytX7u6YAaAbAzh7ZTehouNvbmLDHXMNkQT9ahkugPcaAKYj1kK003o3AwhmvHx
wAkmqgPqGmDIg3uSHkTgBLCS0bk+1DBqrRiUJT/7IdcA5Tg+HIbNaIzJZeNeMJ6QAXe+Fq5qg0jl
d2jWMlXT0e7iF8j8lw3qajbFrhjA4z9n+/KzCr87NSAq49g2efEVAzW51B73vwubUDOlYtGV1VM3
8eKSDj8huNA55KwxO9+m6Kd9B37PUOjYqc/M6d//qVyonbHZ0FZxeCeCUPyrCfp9ZM9zYBOrU+OT
on4AtR1mge3r7W+7ptbJQdcY8YM3NM16EDYhRrJ+0v4iiI8SS8IRjC9KYj9Y2CKxK6jpnPsTehnD
WYFyubxc7DS9RVDJw/Zr5Xs6hlNp+6DxiGyPZN73oe3+aceZxXMtIXvSVVMX2mmr4ti0zFQlXZ4h
uf3KmcVceq5PFKNfPnE9U30jxBhhxZOVuiWvu8OAsqtw/xNmBpePgEPCRhKXSFx5POy622mDYwFm
qLuj0KwIJqxhNxbZvMLQfZbwP6bUB29W8U9o5fkldV1o2A4RMUROo96eAKPhBf1OZhZkvgs6Y90F
/BF/kIAiUJ1u0HngHzmgFN/e47vBw9FOiAXLpUweVFChw8Gxmuk4JJOHmjiDbEgmWiFrA10YHc+2
Hjah6uLKEkfTWYhoHmfVKnVlnkFGidnBSaJmYMA6DeTzPX2ZqySu3YEUfLyGtL9fx8s8zzXyJDly
IU8Zc3HsSLmg3U8igSKiAbQDcIrV7+5r6MwaGhU+Txo1JJkMZUPi+zXKPNBjivwRELfrNLbxP9Ra
yCYeCm+GYwX+J9tTTGuqhl+C1OlUyzX/vm3GkWT9vK4WszYzPX+6I6dWuL8bcnY5LLn3pHnWrP7K
6KBEoreplL7FAMxQnR3XMlocGdeFiZzf50kPrrjNBEd5Y/0OujvvRj1yOUyQ7b7obeiT6y7Xu3Lh
zrtNQgSh3lvSFqhVGK8C5yO70+O+Mh/pcq039bktFbM+d8hGWZschztzEvVBloqsfTgHqLXUpFtz
xs2gZyV/FaLNdbFzZo9IrgXEBAGCRhLwkkysATYulCNIPppS6GtroENWQvyOQvDy/xHH4A9VQGBt
vFzoa2ciK+lLFLLXt2ijk2W1AU7S4YX5sXXq/RUAEGTRYlIscVBxir+gFxI+1pMscKwi4dGGFMMO
BDGN+qnY0iBnkNLyU7P5h1B1CPugjzpNi2yheFwB3PiDJutoDIdU7AA12D2qgKDbPJ3Di8hmfPrH
sMK2pjDdqlXjGQsRbaWTj6pxhyVHJaRcT2qFFdvQBdwGF8eGp8CmCCAUhsa2Kz+chw+sXj34rlpd
11Tjj92M/h4TLzDM/5osj9tljqlrT4H0jKsrbtzK9ph/y3osuwc1EhiXReBI1FCCIYdDWM1+kLng
qGwhHmO8PR60BdbTTGIfNr6nfaikwmD4K+zdq0R+/xt7GHAuX72GXFcCb9oalKjBHUXUFCFCHALT
tWRQxySUdlbrDT3tnZCyjpT5tnaV0CAt0uUpMFKZ2o1+yxbCjwkFqWZI7lSYlLDXBuaJjB3697iL
6swcQ2G1KqgeWLyEMyuUguiV+nI10O3lfjg1ojIcXqGfo2d2dIBUYxyefR4UxOkzWIiif7qtq3XF
OpkcCZkwo9+mAYd6JtmNJzctwpYsRqNJmR9zj6+fu8k5JTdhh5FoxBCxmSzVPsuFlHuYaEkL6QC4
9w2GXRyWXqdqd4dsFTGPT2T/t40Eh1aJWbSgQqR1bXAchwfZeSoMb6iGa1Q6Xt8RH1vBrNK7t0g8
IoUee8vJqkJV8chzqPL3A+2hIHCi+PjOjADoQXR3s/K928UEXhLsgGWuRQyCg/Q/tse4ob5dqHks
MvbagwLXj0hZLX7Jl1rUC2C75O6pLuWGuIbYd8XIrZTcpA6ZJMLc4LjmBVIlBscw+J1zcYOGEOs/
xPiCiDAA6ogL/uI77unPme/C94uWVp05t6YqikNehl0jc74B9qFQmwYGwp57F9S1mDfrq8jWXj5a
+oFVxLip9gl4bialRf6oysZCh6hfG3sspMZf0tR3J2BS1TGxFiGw5DQTnmJ4jSQyX73vyENxu3Q/
387MyLMdBAytSGn8y/tVPaaQ/Lm5tPoCNK8jW6tHT5VvFED/2q/7ok0CqPiv4bmhwrYqdjYCKIUt
GpRJjw6llVqcdpPGZqHdoQFT3y4WAdzrP2zg1IqJ5btf7Sn3K2CJNTOiBekxPTjh3lNQ0wvdFB6F
pK7gj+y/91Q66Ilpm7rvrLuLRZlS3ZPK6sGP8IA+/ADkI0OY2YnFuwE6ZH3+6YqpCLp+yrLe/cgd
8mLL+53v0AZRh5SSui5LwqLgCMEGey188ZQH/kyOuO5igNZON8cQljqS32jpz3DTSCnKI/R8bUi/
tu9meNu+y9jNDAzoZD6RtzAI1PAhSF3Uwn3pGcxA1YyJSMHpJ3sOGolcI+LfcsPOuDf0RqKvyYxT
RKCaYjNG+E1UcLJqY1ibZ1Bf1a4OqmqzLcPcFzujlMdnV5jRSrYfBO8UYVxZhSlAGdgwrI3fuqMH
cwnhGsCZRI92MHgsDtCXmC7twiLyq7exoqp2DJ4W3m+dllhMl5hAicTKWkdCYMQjD4a+42wTtpLb
qHsGVgtD2XNTzwZRe8cg1tUZkhbupzl19wHm+u8Jp3hHFFXTKfAh7w1ZlRpC9gD2cvnjpfawe1jd
E3vCuA+lKB/TMj6/bBL7qp+TH57feDvLdyX17TvC8iQ+yKrji7wUFBAcm+OLwspfW32bzO3AiHU/
M4c7l2kfivmX2mvGRbKpkfTLmX+/9JUywqMpp6yHdAuHw96L6lw9CEW6Kko+2DuxAShZopHB+N+A
nG/ob9ut2pjCRxuh45ql3+bltVjC1lN2TF65F2/yIVys6LXrWefqjpTk9RGjv1xlr/uX1+3jRI4O
NFjqArGHHMg6bLkQFlW56Kca4clc2HqmH6dV9XMa8wpiCQpDwovv3zDeRD8WwTGWzi5ptkeu4Pwq
GLwOURvEv37q0fvVVX436Os3vlWz2xl7h7m9uvzlvZZorhawsdnkAaA6ufzl9g/GY7nCcQL2vDIL
Mu4gy9K/ex46q+No0UOI95CXBFfN2S3qHmSztpKEPMDsW2Ma5DgvL1epdUBY/In72rAMkDIRERH1
yAwQ9+vHHfYFEohgVn/xWTYhuTN5M4S2QroJsHwzvoznClqsuGZ0uWhVzuh0DjR0A3C1WPZzhdaZ
SRTmhNARMqj2ul9Cu9d0tsDEhWQrF64fDfKM/VI+lBe6k9aZdnmIM3xs13fLbXCLorSXZKZbah7L
BAxc7y/aOzjZEwAONQA6117zSovy+16vwy/rCjZtEG881ARNCzOAspBINWIRVIS8bmR4P8OWodIR
FgJbaBD0ysTN9c+cKNKmc3AfHME7lDo7Y1CDJwD5Z2qadLffSYdT0+p3VyM0c+3YuZAeYTqI1ck7
xs37AcaTKnDhnon5pJnlkKLDtX9DEIAMQuTVqQRZ1keERIXHr+N4IbluzrkhsasesD6DzF1XQTog
hUnBQR0vjkssAeIjFVjWSaeM+c5rdZjLvtOlD8t1/OdN8TTCc7Z8OQAtiDIrWcT3G34XjyP4fBtg
dwL2gfJvIDZ2JaVVmXQG/DQzkPjVJba2e8SpA7Xj0cubwREJ3/5471Ls0a5hrHUBp6LLdW0ciV/4
EtJu8lNDGeuC3ZZH2YwvuWUClK/ymw85VBRAiwFBQVMbaKoQ6CCLIEd16QMZT2IFA8uMBCk8gZv+
7dnnBy3SCA6tnm6qx4mXYME7DH9LcF0DjGRZpGwTw6ev6K0U8vGQgdXfXozxRuwMopzRITErMrXb
rClF8mAPoJssZKdxXzBAmG0p8ugNPE3n7Cx2+nt/8rhGwVLn39sFlPo5cBwuwCs/9IlUl3jbrLPh
TRPrMfKgbPuqfNA6m/TII4dLhKa1GiTY4mbKDEhYmgABMxagZi9snJsURL8PhW8PRsxtuEEbD86X
p1WMBuXt8Vf6Hhs7FRinasEQiyWBkUvZjoVhFN5OXp1a07FLIJ5GZSdE09Odf0fYORPexooyD9Yy
TbIMYp0Wod2hAuWvP6dsiZSDF3mbcLGvroDz9KnS9Bt8VEgcqwIdOVfqnn0oLC3G+YeKqUVFC/Zr
Oauy6oRDgzhMrAEXjhVuYOkW7jFwTWwRJ5MZHjCWwIRa5HVVQ//PP6uoXl2PSd9Fdb9iSjiTgkP0
GkYQSDEJi1lPl83VQvNMj1qqE6t+9EZkDrWNiNc1FJKv4GBREb2qliEz/IMkOJVC9tLE/GUXHu8I
+fLOoPTS1Obk5mUFb9aGdHf5v3QB2E+mUocv21YDUeu67ipx26HjCPDxK55hSbC2NArZDagsZ3Lx
oZDSjSKhbePldPXUK2tsB0jrAUS5P8x3f0Fs+WAWwhgFHJKAEMCHXoAZGGyhfK4KH7qEe0Ek+ySe
O0ymzfwukJt6290FFvZXcbnFhJoKlj5I23CLuhs201/p8ifCVzw2JXB8DTui1Z9Sjc8QkBgfqPwa
+4LNX8megEwXG4kiwuOwheHg5XP6sawX70rDZEJ/2gDV2GYLNXhbUQCERxNNkzS4HtpmLP4/kn4l
2Ej17yMZkQWsX1czJDeoDW2D1AwUY8TMQ4q0JDprrP2LLb35BQaaB9A4+A2j78m4oZIfhV5veDHl
NX2FXgdlLD81Z1lQD3Fisin7ZAgpUl3TBgO9vX3u/kBOZPxCl6aeyHxLn33p6CKy49XzHCZwvcw8
D9p/SkynbxsY2rXyTxMX1mhlJml4CN8zNMhERzqml4tPuMtY9dNQsC4rWdUFlSV+ql3WBu5RGP9f
FA3ElL4+aA0kpW79nGQN214IKuiFiUOZUZLXKY2CMRo+PiKY/dc0Cxd5+kVi027EPAl7GyYVxOiC
P4b7Vgo9gU5XUld8u2M9n6TbQNukNv3UkKMZqsr/qHw2U1ZidDRiHyL5OoO/FHMUjBYrdkVfZlan
Hcj+yl1zxgCZfdd1kE5EKlIUki/ZZ8Aw1o4old45D8xvkYoDGz9SM1hQO9p1fEf5zm+8DcdK0RpA
O9+AkFJT6CZ4j4Ahrgq2RB8aOJfP/kHzzhzIpFMzXGvI4Sx+/fiRdrd2ArCNlJxUkjN5b+h953Zi
i8UlSEG9ufUkUappxjOliBp0WDSGHDjJjDtfY0/oxZylfoaa4tsGAZpFDcgNURquK6nCTQouVkfP
W0KLxh0/RBTpP/saqUSC9ZVnr/u/I0clHg4w5e9NpyKIleNXCVHyiRqLqNUXkadQPUCzE7D1o6OH
8DfUNn0vXN58256DN/BOr18yMGLY7bcwZznqKrKpH0zYZXiHPfqkJWA/+j8pu0r+xUdLouxEYlK4
JYoQLR9Rxr6gue65zVDukdHfbC+LLTPcyTVL3VZeJvv3lU+6ji0sElnedGDHKKivk6F+ntU5qKfX
g2YW8gZC1IOGaXNWsyOdbVzboCE8rYHidhb3q9znox/UhPFNiSTqwUa1q+NEJtcS+x6b3otJ9kQX
+BG9MuycIFGzN+w5ryMQ2wI1MU3CBQ7Kip+baO6caAGap4l/o8FxlSbtaKJ/xFFCxGoV+yNpo2Pv
xqsrFagP3Qw0M3PzvY2JBnJitXPPQZC8o6JCK0UU4UtebYVHIe/2VBZTT21EKAU303+Zd04nA8pn
zU/EJFsVvAyukU0w0UZQcjpCv3kX6rLgzQDux/e+IDpjAD9MA+CJTe7cpfYmptvQEbl5lXtYgMSr
BWzauOpSKYMgn4bMYiu8XwlbWHXxb1g9wUD+P/YcjPs+elWRT5rvWpCUJZhZ8qzAm2pKiXW9Yh1l
rwMCLhaj5PFF6Zo/mcV3BgN/g+Kh0BeCapAJsXMQf+ASdWEMwUAmGgijBEDrLCsaskC1RuFooxHt
wYSYI27Jb9TJvoT9vGbAWxEhrRGxeZPbSTpWtTl28K8kGxjxr/4W6ZESOKtF2LYgxT7KQFOlJXKF
tOpKEMPwJUnVMq+wLVPNbHq6E5y7tPO7PAdPVLsglrXtyPfKHnHDAYrFLlY5G9qwBPzYFgiW3EBI
ey9X5Spxzsk5U/6x0+8sAFaVpCa9RnS61Z/2Jwd0XTWKF3rsIgyD0/K/5U7vGgPv3xSYm0qQ3+Ve
l1xoMQv/AzhGnUta0fwMVmpAU755bpym4Wzbomb3vvs/UDzqupa1L+kI9KyoFEFSEwweZVLWfJDQ
RwLuBNbElVS6dCr3USm8FbCmbor1u9VDsgDAGJSiSenPDSlpm3rH4afQzsGya65NyW1qvMmGnuJk
71adDkqSHDxCOGWe7upcDVPFvHfrSDMn4JVwr3jR0J6612DMH8F3rdL/5Fqm+j8vfLWVCeJYxtlw
X3wWTIaXs/xDZVuqgcmAMfUe2KWdSc1H3n1XsEBGOoiAHQhqWC0Dv+TV6gF76i2l2gnXhuOQ51Vt
+j/NJS9lbmxOjBYCpMMUmLW0q1ry2Km4/XNvMR/bQp9/KslOumj7JL+ac+SrmlgzkMSh/SaYcWTO
yXMUKVTJH2RSjlbwv9QWoR9JPQ0TAQ9h7egi0Cs8qQZTWkCVaHOrTmEzN3jLivZN0wqve9rbByYM
gHJZ+Wj4c2/2B9uIohBqTh+ej4UbEC4x01wMDLWJKmUk6IvYd0HPTtk+kQaIuMHt2SfFcvglmM+Z
cMAEb45fwXd+Hjq1+k8JsGApq9dobS0q4+IqY1TkJQPrVxU5wLB6f2LKmoUhfvLbWEn0KT8mxtPp
kMMordpRwAHPzRXYks99pSVMoUMgT0dn2xctsRZE7H3nl1hLsdG9e3hcfhlrFeE2mEK0Ipk8MjoN
nHHYvIXKb0B9bDam6p9PEIiEcLQMdBz5JHLPeo3cq8nLs+BIy1C4wNz/s5vvLoqiZIJoZQLgZ/1P
7V71G9lBfPXXVvCCz/WYRq6wESQ7PiW4pkM8z5yFKmIzzO+4ap8yFrZxrVbAUT4NSXFI359v5TW5
EQIZ09K42nTAr/09k+eOro/Ef35K12TL/+J5O4rtYuRDsF6uHVWcgATVIZjE35G6rlMqe5uakTjk
ewL2qHGIpvVq7r6bxdrgwZs+0WGzMugipb+VqwR9TMTu+iZiZMfKZ7vL7jaOZrgACQzqm+RNz/b+
fqLsNxzjKpULlcGcleUPRAq7Qgr/87fcAxDDh5zzqQLuPPj4mCkQ2TH2ouShxsnd1IdUuIavMfHN
JYuIDLiqCAETS7jyzMBS+mpHGJJwLN+RGkuYu4J+dLB2Q2lM2EbV3QG35S3dkGVkaHmvizwd68BD
W9ltrZd4NNgnanxqH0pmbXyIaJXZDMrbu+8Kn5NdkHaiMG1WaSH/SR3qoQCSOpeaOkkmQ1msJ352
G0PnxhKyNhBm2sTG8ZKppL0IFsAzmafdQoILTdw2YpaFc8UMh5XoMsrGrMEoWyu7/Gk8gZfKrt72
C6waq72yYuvhpNO/0IzpSDcRvjbW4RunRvIjCdm50aZX7bqwqffXeoBHJdS6tLql1jF2Xzz0vBFX
XKtykB8FgjeTyiS0Mnro5onzJDHk7ZO0budQLhBfgkI3lQS3ytprbG+Wg6pLu0FZWKhQiz2wNbF+
OAhpC1EVvmTkCKcBfwvGyxWNWfiC83ne4z3xehc8RENdRudjuWtsbf2ItaiG7fC78xvtiBBv3POX
WPi8WVJoBRhbjyxI2j+HGhFi5WBtovQqPl+PXjHcA/+YCBF8hRW19XonEfHfLUgGU0O68emEGLny
/VmNy83ZKHzzMFIRvwtLq4laTbO05xZoAmaAzb2GGUYCUwA82KuhPVlpGZnIri1akTVmi+PFyQw1
NiaOiUcQwGhPg/Hl8l3JT21avIdUaiqPK+mduaA0Tt37yTWIFSBVmmSsRuSr6wf9zVQYjxnOmrPm
5xFTMlssI/nI+88zJUfXg59llLqXRYRqQWwKoZu74Mt9xKc7/dwuUya8P/CsE5H82mra4T7Jbe5d
uF3bnUvMb5d/+7zaA9BQv4b+6jxdR6jQs99i9QLWgZdnEL9oUeTvu6jOs8MS5TKdmA9r1aHjEhkE
w2GS/fot6Cxl6n4jJj9yKtYRJgv7qxpBxIq8nUB6dMozmGojAzrW+0iqceAuqeFuMsqnNltHkh/1
FXfVySpVAskerIrkElJXltO1TBErxRC/WGisXxyIAPYg/nQMTlAkS9t9JDy+lbCRBeLgqFWH+QlX
5lyey56Y8+i8gCwLYmD6s/fc7+j15zPS7zEkiCPPohuBTypXTfqzdda24QKb+EBJrSHnDBWpLKGJ
PriHq+R8jqqCJMjFB+zfgPnTBCOhm2ntCZ+2flC90EL6vp7yShkX4lULoSmap0PRaqxYiNNiXOYJ
DPsNJUBHrdtuUAxfvBkU+C4nq7YN1kRIosO0a0+PuUa8EUZ0Dc1lKijpc18cVy4ycgpXiXsFOgWK
xN6Tq88d5TfPq5RFAN+3FGIdaWtZjXKBlTHc22Mr9vFhgg1cdcYs0Rr93fbjLvd71bO2hymbNqZX
igx9gs6/6kw0WVoD8orZbYp4NdhhFQupxcfyUSO7785o2r2JQyCRm6UST+23A5eXY9XC6l5uJWh2
tAJrw5mLFRJifqKAvWyneUbfNKWAiV8VdY206Qj2G0wx4Bnjv5d+wZUe56AsctdexdrlsVqFACjr
Ue+f4j1O87qXIuLdnJCOGzZUN6RhG1EWfqJVDYY7cS4JExFXY6UbnYAMItSPwkcBHyMLMymvHJFA
5JCecMeUKNYYOKcZ7F9mWTFDfyDv2OoB/RV7JD4r+OBbexEb5c8g0gdsX3YusI80D+hfXtAjWulB
0gtuQ8ZOsR2LK4JjXrIeUILyMobTdv7V2ABg6gF6BaMqOl8jYhDPGRB6/BQCcCB9YnMdRb9/800N
M6PLLh71zAXbebt9PxyGpiMSlKoi2HIjLqKNGe90TBMuUiB3BsSywCNswucoXS1nKGtwVqestrTg
DdSM3KW7HEQYdDfOUBZxP9rykazRhipeZkwQfvGn2VwG3KWmV3EJryjhxP3Iguxxe9oSKX1W+bKz
oyIPXXrRRW5CYkVyJm+keFHCGjUbD2GurFIiYEY9hk7SJajU7VwmGPoRcAL5+mwp6jnxm0ygnZYv
6s9/NFSnZz03OAdfdR8O+wT6b5tea83kEs0PBEstoP6mi85Ph1laRXM3SK+/7I8TM+WAPQZVjMDO
EG2bSt4slFtcSGCp3+CiOkUpBjv53g89ZKAgZN6zPFFdACs2pi4sNhazpi2xt0LtsCwlUoyRR5nO
G5B4gFlU4l+jlLhvuVrXMHPxEXY3g0Ruw9qjhXk7oNhEQV5rxEMiEoER9lIjHmUCXvJWdI/Gc2oE
CX7LsKyscj+mKlQPiiusFdIUykbQutPdHFtA30t89E/c3KDfCKLKRtMa0Qjt4fsk+iHcthnIPs7X
S434xHN9I8N2U1od5PJx2GusglfpKKDRngmiPt0Aa3vHiUtq5ytvxxPpRYiGer6AymxzxDIuaU60
2+7e9QW0sqcvTC6JPX1dp8GsHefF6tSCbhLcUSlM8hQqkhPFS2kkd14uS5pdzB77oqcTShsCS7p4
a361E3M1Yf3kerP8IS46dSkIuoMccP7a4JDzjft85fd44LJRLAWTWWzHKx1MmN49N80UcY95/qDQ
GGT/Ry4sCKPdCAhqK1X/KhiLaPPkkjtHhT1hzYhVBcoxeGk1EyruVvP6k9tyONk5k+7qwli6FjoE
EEbyiK1tfhk+IQTL8TovKmfsS13pdGtXhDOhmg50+hDVelC2/BKelnqv7aUGkc6jhXz+qZ82bPmd
gjUbNlpQqEytRxF9ETkgpp87V6AMbC5HME5YjsSsW8DOH90vSghUj+RMBWe+o2uTwIyEUnctLx5/
uH0x9b/Zs49PNnb5GeQiGWR64imeYJlrueXDAeobWINdC8sBDfL+UvtqlLKezTQofRR1rd9ijnOO
q6Jhu5fzl2XQdmATxoNhNrMKxKopd8ByypfA/mNlC0ZSNuRgRd7/VHza68lXalYoe1uLGILtDPAg
OgAvX7g/YTirsX87sF8Fd8SuqH8znl0LdC7/kjtS7bJqZdwx/E1IR0sQchEzjcL49Kd+iqAVRNNW
YpVXHMYx9ZDuh7+ckLmzoGmyOtSxXNEntTUmW/ppQUV8KDJhie8BL0bZJ18EiUXF5xOQkPZRXmtg
OM3xlgYZEZjG9XUSMRdKIqkYTZiGV03NtXG/diK/fbBXLgCouSvhIJ2yJY4QiO+za/5RP0XGmsIY
f96qxoGBuR56Gx/az+1XN3mFGdVA6pnX7Lm9YAcVI9Snl1GWuLN8lCN5wZbaI+RJdGpmZqVMSMV6
4uwCHCCVCvw8rBAJiaAt0g0EwEu4wtaoeknnSjU/aQ7mF/kpRWTgFfoP5qPnR67zFOznVEPy91kT
eDZFBELT6NzdyH41itAd0NfRifNIcUH/PG1lmPxX0V2Z0oSEN2toTz501j7SrFc8Qq1DXx7sdrzE
3P3mRR1yEUgsruhQXCu4q+4Q9ngHxwJZYVdg0fz3ey8B/J9m/CIQbKnUTD7Hkri7W4wAkdhRvvJP
31EAI/Jft0DFNgi1mK9C1J1LX0fbBjdmDzPaY6CyYPqL3rttea4DDMgBTtD8vnf8TyaaJOuDxS2r
PFgsfrDBMk2DDzXYGH2TAgP2k5Axj3C/r06I1A3VeZiOPGY236mDd5VPsCRQIkGWCm/JEMwkdXre
OplpfIR0yinYRorJnZNwgvURtDHro3ZEIcJaJ2p7p1yeKq+xjx0gDQidIuJnDw5dywsihA3I1ubU
U6ZtYMYTEwlzU68luQO1YIOaAvLCAN5et4cSH/H6wpiju9CDyyQJ2qhHWiAm3BnyLSDoq3xcFY81
SvkaXpgC0cCFcfKdKhEi9Ds0s/8NMLYpzmEwZvyAjmWv9HyPghd4XJuBficoEl8VK+mvKr4SlMvM
sqIyxqN9Dz/1Y1USn4kHRS/eJ+Tsz3o5WOm0ORGSNMjHJSoOGtRJR09e9utrTsX6W14gOj5TuyZ7
onceK/HjePPbwCuwPcrRijrkqiqsTjQ0MqAHwAGw7URF0DlV70XUhBy6jg+D6xD3z+9u9lC0Twpx
8kPBZxEU347aqfNgMbGr9ofceov0hUF5vmBQS5uvaJrvenwLGRaN6sH6HMdnd1Nlc7FsjkZRgG9q
3SnJ/jczN8AqVsBhDNJMWeGoU8dSKUUMfFvkkYvuZMBqjyHMlmsPg9AM3Fo/GmEimigxis7ULM/T
Bois+g/UTNU1Sp4d40JBzcr5k3+HGUP8O/KSEiiHToHQ1JfugqwywASkC94P4J9Du/hOSPi90Qcd
wGB28bGdRqzqi53SHCx8xNnze/i6UwHUeVRjShAlw+c2UmB+vyFMI/ikhGmGDRYDek/GIgSLTwhZ
P0vGSwSL8GmUnod8KbfnmJO1Rdlsap2gqeLSvW7wZ4M60SDof0oSB8X6YK6pWMLjrDpqmxfr4ux9
YPBAPGYjTBS5yaeM+jp5OXWY0jaDz7PXMCme04NYB1opniRQRZfHqBX+TlZTMiSVb1hm3RpDFke6
sDeNE7bnzW7HJogDEnD1G5qV4PxREW0Bf32PrCyjuxjKWC6QCm9wL6bmMQsfK6Qg/bJh52rbPaI3
kyjh0mpOAgpKs/yu+TH44yE+WhJ3oCihnFDIFYTxAzoXHlwTPVnmSRis1+zWxvJYHyRwPce+j3wB
KHv625kXLNd34dSMOBDdEiq8zXbERgpozQ6MpVXKZzixitUKPWcbMDWHrW35rdZ8z/m/1UUWjw7D
Pt3QN4llqSv4Ipagw3v/SxHv0epaY9qbkCdIzBbDOtRu2HpITFHADeu8HN2gyRhNpIto5X2zJyZU
IOZweduUG25xEEnqxJqQ0YhweRJ0DJNk2+S7Xvw9M/PgZLkLocXlgzQkZ5CUe3JxGvffcEJuKBja
2s9+Lqv136w8Q9GQuN0P6++GvC1uJFDIJEm1KFI/wK/ywOc50Ofrc6Q04DdEvDk2XDsL1rsTI0mu
7FTzV/h8jGThlfND7ufOjr3WUKXXu72NmY8tjEUyEZmC5WygFb4tcokV8oZAixQLsTvaSaYDakLn
p4QD1XoliIWlBe/kovWFfvk9xHnhZZ4+0YX+W1m1I0OVWJGlr/U83+6c6e942dHO4mH3yS/6e1Cl
WzYMMaH8a+J7TedwEyYuXgq/IOZvzC7bPdkk/t/CX4Jg+EWn2Q8i7b7JqUivMj5funwo4Hs1uP2r
E6Wtcx8hR+ewDe3DsS6dfttBB+ljeYaJTnZrqoQRS2t85iZNUPEqzaxCqatr9MU1hGRc/ruGnuyK
dZ5C8BX+WNL6cNNMwJWgs2YlsSbJngqCcoTELniyCT5akq8cP312K0Okomb1KF1dWhJr2zFWreZJ
lObYrCB7kF1nka/79igATfqkN8Z3vXXMQu7qfcdf9DuBmjrvT0gWEWfGKCTBp/ZcgHDyfDUKfdeh
SNAgbocHUb+pdUngWM4wLthPkC8l99803vu8Yt+wD7UqniWdQqdqc1Qt37w+xcPsyj+T4VEzpjC7
GA2GoO0Lqkxdjrmzwx9OWfttrJ+hksXdDxFSOwhiUlkT/2tTlH1WwW1FnPxR8xFwf54mVKjdjzwL
OiKLJ1+6a7sJ2t8cCTeZQ1p5Z4s7LXt65sh1/TqUxx7h/MEzpuQvGvA/p+B+6hC003zDJAy2QBNK
PPotuxaiHIcgVZEAjr4Ukd+BUCO1b5+IMXbwK/6R2e2Rb+WtaheO1ccqhmb9rWUJcV7z8UyNARz+
yzVQoIfNxS342twk7rhY2/1G40PJqrejgUPi0APcTuSh7IuWezyyNZ0jFSHgfDRyToBK0AJo0nee
dKkNKvlT6f87jQt5CLgDr3xTmzi8gAzp606epgKvNuEeS60yJXO9VVqKWP9RCVNpiqrj+ECBz+M3
wfCCASo8lLL8LsI1h9JiJpvKUPh3B1zBId5iimG3+MeexGsnYtpfKfysUEbIhibqPB9cUYeqbiWB
13c5tA9yUyQH1dcDFJPPDu/mMV1Py1LPijpPp/lJ6NlgqsDg5tnu0/4nW5PuXOYwKXq0417eGi4o
0xCITIvvm1LDxBM8E4U9Jkht5MQYREg78QJ5WBxv2+9jT84HP/hcfg5fG+LzuZ0Yan9ujKriQGdb
o4chq6AZLXc8HHliVlqwwaQw45qx47Kafi0TFQHKHGEWG2m1+ASKh0wOsVKjImAQcskP7X8vvyOa
tdH662PL6Cbybzm++/KPUiPeTof97Qg8pQXwylMxzcp7KQuSI37B8REHXItJsttyT2EgyUl1maNm
k8f9HHkE641tBu2tYetrWwL6jTqTgDV+x3U3w+IXTiEXWQ+9AXB1olXU6NiA45f0ILXkXIPPH9VX
04xKXkRAcP6RuUrk6rriVm/rVXZbbON0MAS0U+m+cqHMuALfbJ3tsCiSfB2jrfUfxnfFMRnPUAOm
a56LPtiNuuIM1hHUyX8vGjX8ZkPkr7XuBDZKhJZYMoSTUfc2Rm4m6HUh1FG+Vd/PaFy+Qr8eKYiE
wS3YZRCLSTzOq5Nd5uHGT2Zmdxcn/lT/NNHUDWuHVNSYcVQphzFl1CdqdYU7dKaiIjAXXV2uj/6y
q2I+U+oR91E2gXHvc9y/Dh8eC0cz1IYXxXJPYErk3ZYiejReRFeF6a6zH5XkY2ZCd8MyQ9d32etQ
vxVhFw5IzZx+/BtDT0XcH0zov3R1KI1Pj2IiY6oJoXOzpmbldK+ExJwG8/TG+CSyGyPrqrRrvs2r
0vG5R74Ts2M37g+vLvzPIg7QmnFKDl5nR7fn8azapPth+mm5vt2IJWJROvYnNOesFrv4lTU28hBM
CltpG4SU5uCETCL7+ba6hZa1bXTeeYUesUgDOFwSPLq8lfC7a7tnf5JsyU+ivTaJdwZn+GUOcXEh
e17MwvRCu+v1lUFz8GcmQBvDkSbAOlDg3f1bFYktNVcvIS7Kg9aqppi7vaMWhrT6FueNErdN3J14
7CaucwkP3uY0/eibsrNJgubUn70W9rGJRuBmw413ldSaMGF7DK8EPalplYjoHNVABRDP7vOD2Xc2
ob/O3j+5yFHq6b4Cvm857tU7Zn/t6X4oCdU1Qy6bG9Mc+ekvA/k3SI/90QY/35DBDgv4igtXJ827
hScH9De2cTtA0vepZKt/W/pBK3OFj1+zkeu5f2tYp/y2hB3VtG09X2hn8hk7Y3+dJh+rfKxGzttK
SfibczaJreon/vfwTMPlh7UAM50vVhNpzBUn6qjNDacpqvy5henahBHcb/AQSoKhpUEdlbsUdvYY
iz9Q06GlEyN6lzBc1XC70SyIX4sfHX83o3PdRoP60/62PfhKiNc35Xn07GCQyaZKqPWp2bWvlAg1
jAmcRKZlKBdAv1pnMpbGim+gz+FDo8Y1wazosjERO2wk4i/uERTslluSggBlugGC7Aq+qFAWtyjr
HUZWdN6ZNFt5RTdzM+3jcGK9MSoZxmNinAJZh/vwVOV/hBkCBv4oFuIGDeW78S8EopZ1Oyn6HOsa
RcfJIDYi1008K7SNLUbbN3rrqXId1rPSLYmznmMavbNhWNZQKG4xmx/rFLRb8vWYr/+ahMnsTaPd
P4PHZVsnXaPrOX+rsk1ZbYw25042jt2dS2j2Csg0Aap4cxYnqG83GTJCDigfAr37PgYkAGw99sBs
WAKZhi4j3oafQvb3HH2yH4Ob5DFEJQxRV/57tcF85vJa1mPZ1+ByNpvtNR88lQEmz7Rm6Z4OrXbD
gKQ3a4GD7hjUJdExZKDyzBJ+6PWx2UCVbR5b6F4sL4NL3woswpVQ49NqS9o+ywtIfuYbeKSEIJK8
e9gcx0V2VgNrxVZuN3HE8cbCYke9fuJ+9S1wxQHg6AF4oeFtdUCQ76O2M0LDpwgAosykFvlavbie
KhPcPxiRrWkexXX0141A+KfC/DpGwFk8GwckLvnSwGL58WSAUNwMCj+xpJ3zP23Q+Z0at2NNcAC3
bXwSjWhGqkMRkUJ5/f+uXFleZ0hDRvc8r7nF3T5llKfhdzhnLhqkg92qvCplPqikjO6ohqZrtqGR
Vyas4uGbNvXQ0FDeQKYJ5zH4YsTMIvb6Xhsn/gR87ooDSecUx7kdrI0stvmRedHB1+tDoRSmzfC1
vlft8tt2b9L8MzfEIbwaQxk5KnTZeEpS/mMdzk6DHz8jNie7Idox354l8gzS5/CQvtdKaqPkFr20
ldKnU1VydhDtDsPofcwJQYoPt0qfK0xFZ9tVWlAnl8u8zD+u1wHFjDtmhEW1T73pviB5+Vq0Zm/E
zgJJ4W7NGUeKn7dQzrEKgS/Suynyn1s/yd8PqL1YJcJtJ1V0PJnR6wBUIz02JHYIVcbWmGNeUQxs
fxfipFeEd8/Sg+SpDbp2GqW9xUSamo/l1mr/TAq6gwGnkz7p+gYB4lyrE0TiPV/hpYyRbAnYs5Pt
DATLnKOfoH4R0ZfELCE3aD9i5vBn7X3vG/SM+FjnrpX/ToPHQo4zBPwnPz6HyEKr+kfH0cvrib/a
bjmw8kTAwAX/sl4LqjGvMQ3oci8Jx9Pn16f87K3GfBZSoo1xj/VipVg9rNqzMY0rErNBO9oQdSyD
n38BfksO7C3QNufbbm1TBsY0MyDgcMK1yPMX21IsJxBiZOpC2zvmUdZJtcnGdKGKCYC8/k4nrjuh
S9TlnrYk4vyKiywVWS+oFSPUZ500TYOFowxtoFzpEBt9Z7drWooDITO/2P6eOp78KQtaPG8bTzyW
sDjjDlUMxZ2FVAFGErot2n6OpvLBb5jT4K6U50DHEfNaVshYYGes7PJTkNl3vq2DBPn+/qH6bE+c
x8T8MUJLBl1XMrCec8lXiMnN63oBnpu9ftmi9ME4/LgTJuhG2RPfrePsAKNSe7EEBESTO0lVKVBj
BY1/QZg4o2xTR69+2iKU4kwoqNSS0G56w1Y00KSAsgpkKsjcfGxiuuTW6W4yz/ULcZErCNGWBu3D
mwD6xJzcSjszU+Ze3AagcHtEj8xwgS31uTD7F1gaeuMyyys8NoXqhrGNKHgy+0cR3x2b+iwnMyRr
LYdWQkH+IgHM+U4FGkxpuyXyY9KuRJ0UeVdnsLQtxcJMjw9urcY4vEaLMZooB1q/7M9m0D2jE9Ur
zg63JHH3TPx3NqhgNZu4hkzwbZOuqcxGsrflrXzb1fCZwsl5YJveTapWswjI8pkSsICPcRnAJvt6
vV4RGu2pdeCHmYgUqyls8sH7rZD31BlE4c7VazEUVzqQdxZY5BoBxteu+4jaWyA9mTTMlwLG5Rhj
9sAByAsqu8wur5n++AqlTU/e8QXXNtvzXHdJtpoHhrKN6QYFznJJwXfCL2tzn0PyjWxvcWt7Ky/I
lk3nQ5PvEMLlJVOV8x/60am1bHYEA4AfjznGllHEWrCk0FSO6Ehtw/e3XBZmbpKI1x18FC+4zJSD
9Htt6Unb5X4bRxDB9bi4p/FBgIqyg2qsW0afXb7BrJcsC3KtYAYYVcMAGyBJlf3OQ92p2Sd3fwXL
4aJjL5ZMpj6qXJkiKkXEHzsxlSVgYeXbyezln13Dmb38kT6haPOhkuPgclPByfRqu1/VvQ8bl26I
S6wYkaSJL+ziFLUczWr67ZO1ffEtIfp3ebYLmyoGFKl/uWAk0X4EP976RxBU1B5USqlFiweQYOF9
QqZv9V7gAtEW4grnbc0G65Yso81S5WH17PK43H5Q2RTMNvVlKhXOXS6IYZd6i/lNwfbno0W2cVuE
0aHvwnrwD+iMZT20iFpMN4+AP/of38bEyPtRCmktJ5xyUYXW3qDu85RGsEVTQVriXPsRo3Ww1eH6
B0l007o0/v7W/kY/E7VJ0B2l6J9vSs2JEmvcU/8ArOwStQveitlYkAZa6nzRdAW0whyyknOclVBq
7BCm0FwnSCX7QliootS/MDlCtvIkRFy6UmfVYxjckUYd08NexYXZpI0ZC09i0XRqCHbE56NHISdG
cWL2+zIPVBuQ51VK1eFlzWWNQF0NFSjXksTBkOvP5YXNVwi/bFtBriaoSa8Aq2X8UuhsUO1E5FEO
ONVL2yzPjsUpFISlYqUgkTiBhlC6u4D1EaGkKfGEuZAxgqbXV/YB2BJnjP16EdKeCkVrS4rBp4bu
auBf5O4JR+mQ0UBiJK5w+vzm69b/LFmcBFiSSNGlRT95VXWEXt/ChD1iF59NCys6qTkZoSZ65LFp
gWTTz9kyJ2ME4e6HT4h4xm1+Bg+oHXDm9OZCXPYhSlbik4R4bNuk3auGDr5ME0ThGaXYJjmysYf9
edHrSzY0S6ENgBDgXaHWJH8xrX1MrDbotidW4dm4MLY0EDnXPBKVUAKjw6ojUmCB1d3YoLFXstD8
22MFiNL8hblFd2jTD/BNKiR7OHLj4qy19nuLBod6Skp4DZhWgy5jy3mu5fDm125ts+CgbsV/YzEe
Y2OrRLGzXXECpuJ2CcFSGvnicowwe07cDUR23t9cAecRoRG92bFN8+Mwv2pBGHRIGHvRDtb0CsFk
hDzm66qdELhvP0rdE04ofie/JkCsv3zT0WS3LNKiIPny4C5YQvurbQXDWY03ehO0YGI6EMvFZ2vY
cHRY9da59or4E6Y8LlSKKKZCAXvRZg+G/KoRhA28SSL4c80rt1EOMvx2pv7apwlXIXybf2myZUzP
1svntkY3Dmrma4C2PcxqymXX9sLMQCcTdzoJJWSOVxJ2WKgj6SLlajz0LJ9+o+jsU/a+3hl35BOk
lcsQ454DLry003Te/nEroFc1SurfzMeZXc7+SMrhJ1e/Y+dQthpeB1ezhuF1LaWpMS6iQS1ca7+e
xTWivDMR2akj9sYnLbCElogr7GeD1zHFTgEYVN+PubrbOtbyj9eLPstU2Zat3MyWxAkGVT8xIX+U
jb3NXw8pMucorh76Obwh6/yETCrLylUMx2XdxXHfnyQz5bSuHNopHf7UJKxTz8Saqhs6BS3YGrix
MPlBy49NZ4ZLRjtP+OfMwbjxDd9nZbKHvQ+BHRxVs2LpPuJ/TNKkTAonLCzj6SGiihnE/+OHTjvs
tP3ya24tt0qynLEdEuc4yOserJ4jZarYPSFojoh8v4aDf3ucTpie553pCS+2SCceZhQrjWRPl/eM
4eCHCW88mrdXr+5CkdQ+CaahE7pZkct0m4LFtpj8m3anHLSQ0IpkAONyAOrAoTbLgy8fSLd+kjZj
aP/TL5eyVBKBIQdWioTybExsTSyrRes9FWdz9enngc4LvJWxfqdg3T5yKLVBkuOZgv2W5xws2a9r
IFwc9zUYGNxtF0p+AFMpnwuGAyH+mEqfxRGmrAinU+btFRPPos4xGFX2JDJ3qXo2aVuJ9AMszpq5
wF/z0N5PdCpky8ExrkvfWGdha+oioCgD8ke7mQwlgYSmIOAvAEXESKBgTsfxRdhujJQGX1prutw3
9UeKbjOl04Sl1XEB7Lygu7fK/12lBNpuePGNNzhrJfZITAxQ0rgxd6uUHKk+xvDzEDkl6/zxRz1R
F00+zhno4rH42bu+fDd9piTJby6t3H1odkODslWv7fqzXiMvjrI5XiweoLGQ28HhdFZqvP+Od661
Q1uYt27vPdOfUBlLRdw7/FGZyQbvEZRnlYJKLi17nBny03amSsANPJxtkPPmWRKHjfsJ/ObwnYYK
oTjrK3/beP6qTAvdDcIOdvuxghZXPyvMa2wudf7JLmlinTHRweZaXVJFRGcFQQvs+sw6DUY4G40n
Upg90OOwdVBwDctxlJ/BD9mCjmvYo0yuPpg5a2CktbxqF9TvVjmYWE1xk9rRtNONDOKYeIqp+zXd
F8lMHsAEpfRTruBl3rVAPEXighmIJQxJIKHVPJY8rr0FYEU2h0vz277BbBKovfklYSlpB14GI2tl
gJQaTv6uier+iAGioBjHzgOT68Va9gr1yOCo6HdMEw5Bvh1+uHwRUJADIRD7V/FzT2a5fBOo99iU
5NIqnMxzBu+sjhhmwsAAgObVGBULryUHV9B/tv2EvbojTCxNSHLJTWErmSOoHjlkZsV04sS0mxPN
paPHMkbeTUqRtI/vH+JMJtc6WHsWFkXKIEk66CY3a+XsXqotwh8jXS/J2JevXV4KeMDMncID6Qcs
bfPrfnDYkOtPQKdby+cgeQSwj1uIGBn1C9MpI6YQQkrhvvsmyhJsKDcW5vy3DkwtyDzPlw4z7RPX
Bc3SuXKDrrFxNvrF/ZlJr0J55GKrrE5R2Km4xlJegY8V4sabJPgBCzMDM34eIZgNTRPIp2trjyz4
1ivcQSBshT+FvlGnjcCQkLqIiAQBj148zNIYPPDRd5A9DZiG1U0SBizzAd9eBq7oV1nIX14eUlGr
j774LZwB8ETpJZZ/b/YMaV6CyyQW+Rak3Y4ovQQqkDXYv2jiyxUKxSdn92rKUbX11XZffgr8vEcI
5Rgrci2WsKuOf9a6NvQUkEQ8yp6DC6Z71Gxt4DUeqopc6Gb82hrYY7pQT7pP2mTih5+J1sb+HObq
xR9pjvpCTG8IeZ81NqRMrVNegDqDRdtKextGlzRcS/i3q01e205wImdc9HkExDwDp1MW3+419vYW
q6AJ/2LK2NwDpF7bDEQ9pNyTpRb+d+1w2CEO2PijDxdgQ3B12HLpnzHMik+DrxG/TCNR2mTsG5HM
SBfEIkmWkiYytFVXV9nRjOFbQFfPclQiReFPS1cEWGRjH4rUkF/xPyMUH6spOb22N4xKBe9tg4MK
9ydsnRFb8/kDTl3t1TJ3INW0vWS5bfNynORQAjTQ6Faze9WOgcub3alTd4wfrg7YhISr0plha4QN
2MEanpK8JOdwqeHH1I9AmiIQ+KIHIhvxHcMP5qidQbBQjyTaIjs2EAjb8uV2fjcXKVbYrDAbJszB
yL6sfmqc/qT2LAqsCkzyfasATtcbc9JG+NgUGCVcPL8F1wxcE9M8EhjsS+p9yC8xYZBXTisjoUk0
IphDFlDaAtyA6vHlMsHG3YwXTFIPYMyLm6mLmOKa8lVNzNxNnMMY7p6gn0gODoKTI4K7ue35DL68
nS51UjJVrvSilgg80HkSzI3OKBKw9BrEsdb3WCDq4uktrTM1ka17lDjQOZ8iSbfMPs9BlDCRQrAu
O8lR3qXrmr3atEYypp+l1NkThpF0+83T5HG82jFdy2gXNekRmkN5mvynnKhgDVeFzi9yyiOlgBkb
QZke5LCSSYFiVuFIQ1/WOvJwJELK1WXqGVA2pSzE05/l7zm7e3e0plztWTMtsTYeHZhB4mto0OGj
dtYw2sDqReTqTuVDYuJLkz0LK1PQoE+Y0YamMzfY8AhsGkbp4Z8GIx4kN92fSTbcvA+4DB+6vSUv
1NyAHu35w7zg7F3QI2eeypho6v4nfIcNhTF8Bjy17Pldebyv4sGE2xLlHzIfFhVnz578Qg/Ijeo1
sInipeckp75jmeOwBxQZNhdkAcPUOyud6CO2prwyen4QHDxCVcLyaX7Gy6lVH5Kvds3k+yhXT3gB
KYzwKQXblIOPvuKHUlrY+MgPNVQow4mLaEiRw89VMC9vZC78o47oj2Iq/88gg4AYmrQaKKq4yCgG
Js8x4uG8m9I8UpC94gksTzczSBlh3Oj/cf0eB0VVT3CoHkkNc3ANPEw1ra/8j58F1ZF3W5lyEuvu
tQjNaqQKckmcCE/1aVsIH59aWpOW46KCn3wQM25u/fNjtquqq9kB8FnGlRUjyxOFpjTmgTE1K8of
GR4KHWqN+vd0ZNhH2nfNvpRLhgus6FDHE9sWPec47+mZkiyHCbRwUmURyC1fRPMcZJLZ8VJQAm5a
wW4SFL7TuA3wVTR8em2A+keKeQT8KIgwvfmZSgf0LgbZ1E8J2Gs9utqiEmgGU1cbOezpssr4ui0d
GOZWrCKAr8YUgKBEZ2SbHmrTbWa0NrW/wRCsCPEuwrCoLIypFuszijz6vux6UmorM7ylXVJsPgVL
vyy2m9H9I2X1yhSJ6D0tgNi6nw9r4A+Wh8NTC5mbDnHRi+vM2D/xlbh8hTsH/amfgPYYBUKp1/AH
IIi0dlTQDn5hVQ1lSWMA/nHhEAWBbaTh5mz96UcHp2zlJj04t5RreP+joE/IAq+d61OOdL9NPpUk
daLaQS/BXwhrE9aQEduFerzD8lIafbjOexIegUyOV5PrnZilLUqgrn64AbrNqoaedmbwHY3ALpMv
a5+lvg3fZpqp487hjnPNjJBebfKDDg8ZyJER53ib04KqSGi64NAVTa58o+RGkKNWlF4UC684rcTN
zFCSwcgKoCFLuA7RR2mt2dCu5hySKk5y/4SVvUDs6mnIR11atdSC2WgnZPhvyYAmLmHZcDp9YqRn
eBS3FmHLTbgBPTXGj9LwQ3yYvL+sJM3QCmLquzGel8ijLj6KPvh/YeS75p1YkupdPG2bJD/f0j48
xXm+Fuojc01iVWRsUeVM7P7PKUTAZcUHWNMLF43FcUFoLQSjHUyUtFeAXvvBM/f5QOYMsva1S1+y
duD72atMTzgzasAbFSquEG2rADEmi/t0v188SSqtb+5GqpGmjGYmvU8lw5SKpm2LYWEuDtf/twnT
jMjeRJPTlt2gxkEljCJ8Aj1zmDvAK6h1+taiMrX0RHpc+qpXuntrqpfv3VqsI3xRd8w3zaUWpU2S
YRtvCo2tMQfTEvX4uV0Q7qDdqQReIxhNYurZbxBMaztG/nYmoGeGRmODIgvwdeFLpJGeIvuQOYKs
jxAOZTelAK0b2XhB7DBEUJz5tzB1Xd2j6tfse2fsrw2rODc+w+JmlIz53PkvJQVp3yCGK5eYREWo
uKkqZ6k2GXAw4DJxueAnnT8dsTiY+agy3mHM7Uqq2yBzCGDI02mGqYxrrbPaF1p3R9Z7kenU+ZUV
u9GMC8U7aEX9ihl5Is9x0Nl8OSWzmsUnB3xmXWVi5SagHqEMsJIuQJ7Ub6i4DnkHdEMmshYIDb32
w4Jkap4KpN5KspMUpKc8SklfmlAflnHR0wXtyZalNcLviVH83bLY1dWTe5vVw85RJP0xx5gfVBpu
tT/pFrruokhF80dOsoXVPc9pPWAu8enWr0SsvP1442wMuTyOxRaxvGZWinZagiGRKLcVvNJ1shCw
k6nT0PckhrfOscl4/syQZqB5F5vupPuhc1fmf54KkMeteIDmuYJWYmAGn0oLUwb3cxUgBEwfy++Q
koWIEc4hMI7ANSVj/SnV9pue63Kp4IgkOJKRKUv0XXSCcnuZp+1mh7qCB0W0LlMH7HMip4Z7sYn3
t3L9R286AKv2H7VVgqOn+vDPKFjglUmfw7CqYFHe6pR5AGxTIh6edbca9kRatCd1DTJ0d9wXiI3M
x3NdB43KbENChRUnJtIegdHo47Cb3fiA45mLEqQyVrPSfhnQhoVEdlEeKNivQQZBSGYXesijZHn1
Au7A/LnT5uzem24ymKKt+Pq1ncaL1mCRy/U6JwSAoIA3A1wIbp8wqWAqlqqoyJ+FnwzF4GL68nti
oP5T9qg6SpLcNF1x7xuFYGjkPpjGCY7nmZIAgPzkvZkL2JBpqeQ3Owj5KgauLebJ7hLcYCyaVoHu
5yvvDbquA8Tx0UatPNadBVMwfAAtlAT+r9htjX6ttEdE/X7Buh2c2rAfCcxBQbJxwNUSOb0VJAUL
2GQ/yRGkwrwvp/wDPqxNerq4cwbS8N5v0V8HYf8vn7/JhcsQQIDwqiaa4IzaZ0NOaffzryN7Xm+Q
sl4Zu5JXwwTifNU0z8entp4N5IY0Emp+rpF3d5BKCbTGeIw1hNKmJxHNGUbNl7gFAax7dO3PYeiS
QqMVhyfCm3E/okHRBqDFa8xPdyq7U1mHxqOTGD4QG4nm7nC4nHHM0hiv7tvGd+2aNs/0o4/cXGRB
IOLgSonkHWm2XRgvO3WhzC/aMSOUKr/gpHmfjdVPAdJPste+qMJDw1VmwrxGfLGU+7w7NQdNuYpO
jHD8T69Xek8y5y6mDuhz8AXcmjSDiGZd65oF2wciEhD4nO57QMvWZZmutrf97KxoNsVje8X/8Opy
ACKTZmMgfMtc6H3APhCnCwmWSlQY7GJRLeQocbCjeC6qUDj1vGt+70+O9csz9R8R8r7dHaDXjvHd
8DEZRGti/TpcJCppuK1hnazx1/PDQxZudkGJIvMkPlAfvlwPS/OfCR3VO0UQ+7CwDQR9v4SR0XJK
ujm4TKFYDtjJqlLQa3nKCUZbe9PhJHYPBz5l6edOSvxNneU2IOQVnZDWgxcUeERiZ2C9+KTRNK9O
Eyl813x41x9OTkXf/CSw7UbE8h61NgCBiDj9Mbz9s2setMSPwABqXQv7fIdHoqN1U20kfPEUOQH/
H7NprSP3F2uUpy8RH7gFRwflQEduNs/uVu9y/cGWwboMJ35Zfmieha0yoUi3G1keSQ+d/M9JllGG
4lt7+rAVkvlSW2h9nXEi4pBZaPbeB9u7DZF3lkGvXuKi5/z3O/M2AQYgDmRomNVDSL7+3N1ZMvND
HweIYGHIzf97YuxdZBIs3bzvZTf9UCWqWNuSabxM+Qn0Jk4TEm4ogblzQ99COIm7Qj23PzbA5Ult
P5zoMFi/ZmilbrWbRRKmEDBNIPhlznCKQRCNmq4LpCD2439+S3cZUUd6KbY1fPNHgUKRRLKxgYnO
hIwp5YGMgh+lxAKauDQhjZGCfUzBnLQGC4QGP6/StGiB4P0sihUyUbbyXx8FZD6F4Aa6Rp0tuxzZ
fuaHhimuU22BAmNhgAMnGAC5ZpgDY4wxqGQln01kTqmqFtH22U9J2YDrEWkVSd48lHYdfgfL83Yk
DjYq+1EpWK/4OUL6DUss/R4KW6qYzgDELWJRcHLKdD0SR/cbOcX4yOSLeGqty0vDbhh4Gvtb2L8S
QaKnG+O0cQdsJWFkJzCxMSotMl0zdCxaAp353LJ00U9O+pQUt9V463QMbkls9DVAhyQwvdr7HiTF
wmsgpbl1pggqd1lwE4rKZ12b86DKyFWregxsPUAQhexBy4VmN9wm+3OR5uXzd32RWnsqCepkVsrp
AGiYL5xcvie+cvlpcbCgInUBzcSG71Mpq0Dx5Hx++t8PQyShTvLS72AFnxseuNbmhoryq+WzPnbZ
itfp8KYyHCImuCpbDXu+klLOXAwZksBuVis2NUFw9nHPC6RChqjcoObqvMV9kTOYOMHFELm3fwXe
hHJWFuSfsdnrZcqOrOwvGuq38CshKsuDD42csVkmboXIEPUV+dqELyeXamfMwXZR4atqKT+kBmdX
n9sBuluSQpRUivjuqhFddhfiKvcndaBubXOzNYbB6MKoLdCEN/qF14wUdYAX6877xQRSU/l+pAep
TF4Cz6JUcU6wJ2q8sIgID1kZHfFXu52znqGAUpnR6XpV6jMLUhRwhqUffhQ+tFfsBStvwczUbl/1
rzcXXPVtAc97OgQSGlUQ9nE/1L3c6QSVZvr2bFQQ4GEETdWBy7wCD+VCd9UY0ZMxSZxCMYh4VJgJ
1uJ4N5QUF3tp/0nZQNpoVvez3kqQKronzAFn3mlD8XozbwtKvRjAvc4jCWXQSw53M8TnV1IYGsQB
UHXV1GexYx/O9jvSdcMvYfd78w6LzwHIGiVaCwOgsJ/fPEO5Ps4fZsc+GaUxogfatTzgty5HBwRU
/3+6c2YiXXt+Zhtiw9r4wqW3PB79nDP7+uynnn9S5b+ZYdE+623djeabhoQzXw5SuGmGk+52X/hh
fRX2pa2VpJWjXW+/xuag7k4MbrKqy0JuFm18sY3LA9YAOcvwiuC+fXYnqq6vvJAg3JVszK/26wwR
TG5sMVOvy+kUoPNWyQjuFXa9I0UbR9MvnKfh+s8bEYbsn81qao4hp1+jC3VIKA6tCV84DJA3nZxq
fovVGxNauHEZf9XXOmpR5yBHlwFLA7+4KJ2DIGm4hrXYYXNjIPcQUEEnFs7fIpTcexv+Lkkl9Vj5
NK8R0TGN7KI5/VWykZFH3B4aONlFEcXm5DGfTkS3p6wqm59L7hPxCsNUk/qt2XdGYGUY29US3EF/
HtgFUre6IqM7ofowqQ2nN8JJkMyBZoy+FZG6bQLTjqprqGvHZR0yKApyjMrAMuJ4L5birb0SzDO9
2GMiJCXhgrG1z9gpAvelGefh0hty69XE8E1lrZ3DVIivkeYbfLev2RLcEFUHjd+FvvZi8koMS7sA
jPCQd5EW8MIUEjnqJRbrt0h0mOpgH1BeKl4W2xj+O0575LwqM1KJgaCVrQv2oCipLnQsNmK0791P
eZNsQCUupKRKlGS1XcfGSOAP20X53e/VcjZ/C8FaguRrAuSs1acnRoWYepar8uB7CP1pp1K5L6tk
2MKomJ5YcxX6UepFV5fDs+QOptGJgyOEYOneeCnPzeOvxC3hjGrFcuAv/xcqdknqEjKXfQBJ6RvU
vmTr6OPgOtGMb29KFOlhwQTzd4+Hjhamt6tov3ksO6N7SboYu2b0JSaeo8krOhwXIknhdjT1dN4Z
hrhuNqMP/ouwua9FwKeGxqxR7Ucpb6cC+Bo9qa7uYk6+4MQa/sr9kYbkeihKytNCMuhzslawXl19
6YXbOk6IlGDlfELlsZ7fDSp4TzUUjXogT4VrqIraqxAKIfsvCz3xrkYIResznz6EDy6l2Ox3RdNU
5qElN0L0fU/5i1YiFiN87IwMymAVxVYssBaIkHa31icwVd7RGVxjHd1jVgiLMGe3RBxb/AlkgUTR
hmhJDt81bA4//UTWTb/wHtni5Alqhy4CJfoG+JAxkWsuGtRjh12GPlp5hboqGhImFQpMY3A+Jfkv
Jv0vuzdg4fYqwSCp8uYUce1N0BDJpfxaPOQp/SgVLDfaDTA/BtVDStxwHrCh6l9K9DkUyNwmlW9r
Klao8WiclJ9gUQAKR9qJc6L0CA/Y+RbSSKhU5cnJuiW95MrSKr7XgrxQ9Lmh3rI2Igw29HvHVZij
ryBFKk3kPJW9t/IN5toIrO5VzxNJ232BmThAlWkPzxige0i6BFX+ZydsjkzW5KvFFb8tMu6E+bYm
v7/b7EylRMrbUAIDL2KMzS7SvRj9ndlhhOfMKQUEoSlLlSfwJtLGYudKcKzMVWsM/PBuFeRqHkJl
IsoMJ+Kc2UXu7ThTk+oPZmxaEkTbygSavCxiiStd2Xsksa0fPEb6p2BU/tjpOdQ+E/V2HSn7oKgY
O+zUmEt3jRsxq+sZpc2mlIEs+1i1Z9OqZyZUgHmk05akOyizu7/yv4/QDVvgNNTEulLTJdRHShee
z6Vn8nBgiol8v2cBV1yzKzIRdh2yWAHjtLCyuZNrbH3BaqeNuVPL0W4PPRzkp1da9f1a2HPQEZ8N
/SlS40U6To3skJUXJ0I9fbcWVMPw/+dKXpG5CEJ+p78ySkpcHM1ygU+Vg0+5vg6UK9pLUi3WDcMi
xHbZggu1XHlvcAv4I/8oOmH8UYC8Fy68HTnFdGbBUKcmV30Z1tsNJbQgcNHCjyCOgBlCup/E1da6
A+j0kNNhexx6ew6YUQASI1uRzrZerf7DHkZCccULtuowA48swaJ3RKwB/CXGNp1d8R8GEMi/gfZM
ucS40GHT89L80OcWrHyaH1wx4s/bUTxiCAVI2Yb11Fwnj/00A9e1Pp38n41YXBO2/cQE1gpy1Pfw
X3dn3z+2iGxjwnOd01wcZ2HhBtx7Z1frJvABBTRZQYvZs6SEzmNiwqElEd94VPFjwPuU/JmEzKDN
MY1VuJuqytHLWYoZnAqn/rsAshNwuDnZNOv2pvLrLPGmDUN+PPIt05o9+hTEgbmtLCYrGVEzDnYd
+sjJDAIfn9s1zCU6cYrAKoCkd18E09A7ncjP5jdNGdWiEFlvUIcyb7ccEbAWQsiwy2MyfUn0LyBZ
ABsHcLw+6NsQ6+d2wXe9W6h4xfCI+teUgDjCPGeMAXlJ/m9/rh4dGvoDAbSFExCkiUc9Ygebpsno
Rw+MPcvxAVrJaRUiwSA1L/InsoZuSVHhUoIci2qsjrP5ECqevQRpIdQ0DQfkJKBtPSLivUaEqz8M
Q9NyOImnJ2dNRDdQ2zpM5GPIaXOt79wAk401k66G9ScQLNqqEcfufFEWy9/ePYugv6nM4I0m+mvs
Zf/633Z5BiPNwFoEkqaw3oTR0eWDASfsmwn8pehO1ez4npro14cgIrZh36KZC0N10WjV58ukKQVU
N/M/AftA7GjYd330+xYXWjxnPnJQ5ZNdj3lehuHkyyQNmNPpci2RdNq33kLmj8jH4G+SlihgXYMT
/bpgx8mMJqUXbCNoNo19q38qgykymDwyShN86Zy4sGU96KMbkLHRAgX5QaQPvXkA2CKxOVlR8/vt
2B7g9qYjNhVOeVc7L/Wnns+3j4Pb5pkG4ov5pqeJzNQQsmub6ClxRHAbx3fUDt08nOvh1SWaTR+/
IziKSGM1a5Hgle27dAKRtet2kH5c70f8i5U17ktzY6iywl44z+vdJ1yXHFnBJTmfGpOhbhIr60Np
6d+SLFOYXnMvHOVbjirX9GdAE5g/0/oUiC7jmaFlFh1lYpa88GG1fVidIUSCzpFWWmAqrtgzOa5/
D84vh1CHAzx8Pgzfk9egJFjymWywlA4a80MFj1eyw5Jx8J6wnuh6g/X8tv9yLBxjKBSJvmRQqJ8y
duVYS+rEQEPG0QX5swhzXtLuaSsSEnMprVxp4AA63qnAcRV6oaMCD5Nec5KZ008psjr44vyK6QYX
AebOkKp/g2FrFflg3QBTuwkkvOKVZaunm785WY9wuX3wRgSQ+SsDYiDMULlEzjXq4gK8PCuuQSWE
46nt3ZfWLr5Wm3vUGTiOPZltM6KwBsh4wiM2ZpAiMvkz5vX2xsb/9T4txqnIw9ef0KjKt7F06Jee
RcpNAu53jdAqf4yhxGpGFcKzOfyiR/7JnPnAQdB/PK/9LSQJZTT7B6QFKh45aWGYM2JwP1HTCqqt
RzyBhoLbywoCJR23I5morM/FFaalL6QnIFllqsm/iUiQOSwTYqum1d8Xb655V2uG+yTAeJPQWcBx
2lioW+zQF9eTqVkbCP/vIWNx911jtNWjID1jEaUQf82V1SRU4RtJL7a81NUcAQdzo/5dQuWgYRjh
AKfdjnbEJumWeOGYkOsTFdXhs3ATERXQ0jFvAosh1U10fkbvO9gHg19BI3R0mIBEnkhUS/7ja/4o
3dKG02HG9NczLm/ClrO5H1qgreXopW4nUtIw+y9z0JCNhh6ccbZ1wIBFVjnvTcC0dwxIMhsRAicY
vXfTT0noRfq5JtI0nEt6UwJZJuF5aHulhBhZnpkbzKxMb5QKGhHrbDYxVVd4r27oLcytjDWpoyR9
48TfDO0mpE1agpozWjLHrVyEG3e9n9nTRS7BR4csGTNBj6QoOlKYBrgujO75P1Yha9UOwq8fQEDO
2N9McZGewkix49Am0uyfV6S2xy7H4AGQMKkg4D0Y9RQCmDXz3x0YdvM7nWd7T0ZJ9tlmRzGSZqYv
ioDcBNE/6T9zZ/cEhzbfADaCAnS/Gr5CGvl6uIcD6qSHnaD3u9j9xVjsYdVzTYhFS5Z8A2d9lekl
D6yT1w4w27RZ7ZE1R4LqdOHMw/igz0y2eLHlif1d+ZNsufZcp3dzHJt/AUuVcUcK0WqksVqb3qav
XWxcZnwUZN8rGxMqN4M3XnhNlcceZQgeOqss/CevowRLBLBexMrPApLl9ztPIj5W8rbYIxkUqlop
gNeBGqJvp3ZMxGncX0C1XUYMSjNHeeQCxY/+hys2e17G0J1u1Yb9VJuAQWhG4wcd/XzqnW+wzOyr
s1ZidYOnRSGcIa2raYnW5erjYxZYHr/uEJVQmmdz+PtHog4k2D05JsTtqpLJFhH2FvS8y6e0elRc
SCieNIUj2K4DUXTY2dx/5N1KlEwGj5Bj/GiA1ZpegrZGf1gk5F4x6GAQPsXmtIMkBaSexB5p9xJZ
ulU5I5+Pofp/4+RO3awokhfTU5aF/d18In6itP303i6PMCKDsyefz4JbL27T0iNsCAR0EqtCXQx0
dEvpcuwVGELSJDq9IKreu/lTWYE7OEftwedCBRx9Lx9vF5gMcKLKqlk6G/6hPgTVofPSIBV+SQ9m
mxNR+rsE0N+xFBBLTByF1oSRAib3jvb1cVTArcHlJ3iHd6we5Nej+EfHmZRKy5MVBt81KV7h56Lo
OiTmizjLbiLEY3HTE9g/DjjMlFwUuA86Keeo69Feu+PEz+C3SntBN7MhcAezqrcwsZ2JZEV/F4Fq
vd6QKcx9lr2W7aD45tH1ChzWfZ+T3dGNfiG/hl1lGlLpr+Mo2mjscDhl0heV5BcaZ7ncxmzTpiuc
qze0eSR8pEY01jO+1uBLb9qUJwcktJc67hI1kgnDNOX4dgasvWL67Zn74DhckJSAiosUYiYL2vJn
ZK1WnvxXa4LhxmbnNzJmZ/sWoUvi9zSBtkIoVOZaur+N0MjxYeOuwm8T/6/o24Aa+PWcZiO4WW/i
XrmavDL5Oqw133/DqkbG4yQ+SZSShj70nvME4e085qA3uPE/gd8+E1sih5vyImGOOKorFuxyqWBe
dAJCLd5aNxUi238N8RaqUJfq3INx42tp0LCSkgYsbZvwIYItGf271SSbGHo+whnfO/94olDwPL7F
wVZC956zqjJW1QhnJEhvdUAehijXtNver63doV5p/8+4wAzocIIgpo5ubzRV5nIN7jF8OIoHHJmU
K9VUjbVledxj5vKdNXg+BG/AnNC/qFrYL0L2Qj2Cl0gbsUFWE6+egtiF5WWC85RVMB03E7lQ2pkQ
QORZvDdtvGfi2jFTHwvu74HJh0n7rcbLXJ9+qHnM95DEQe33f35z8lnkoI6zheeFeMZDGUfX0pFS
77umMrDkAnAC9gBaro8h5CHY0zXbsrPzGud1xAYGHSLkR4f8Bwr1lW2jrDxqCJBZVGe+/zrmW6dM
eutnkD/8jh+07Na04RYYMbZg9xaMdXjeBHnxG9UL0rxZ6ILF8uqVTf8tArn3psiZCdsxikcDcX3+
sdt82LSMh/djuJ6bdObsZEJuF2KS6St/kuhPMA7QVVkeS0Tv2DIIdDoct3FD7Q0BCA==
`protect end_protected
