`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ovZC2QWJKasEP0rHP/XmhuRFVOmBa7999Io0U+MMoVKf5ltkIcI0SrzQpkOGaEb9KNSoWmWZb6HM
g1NZfNeTOg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OVltOIaz8HWc64LPvNvkJWmZtTAan1LhqF2SIxsSIFkpHXuA5q0bUvYnd8Ql69Mbj/Z2e85wT4pw
ekcAlhCPgH5wp5iYje9PF9Q+AUJyunOtXRKgeMZGZVzKMV6oKPYS8/thrOJgXpGyTvNfgeoCTd+6
Bm9Mx6M+vjcSZROcZSA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SzbbZ+M8EEvvE41qnGbuDapHEF6NddRavn83xVqSDfjS8x1IjE2T6ypnjyaW13aF8xxOA6Ildo4x
/0Uy4CfGmGgno4IVCPbwaVngq1QwHqoHIvFovmJxMphtT5y1H3E09qyZuSLhl/XIVKwODZqU9OBp
zneG/tlcaqgFpSE11lS97hsWznIyG7oRzPN/woAQNbh3KHB0OIE0XuZXX87GR7NU7MQ7M9HuEIWM
ifECnnhGjhqQL6TIjIIlBZs7Von8chXZdvcIuyDtoPInoB4nS9DDQ3HOYzJWwEWx7/zMva7Wyuxo
WSYpdkFuC84dFRSoInlzk5LozakpZCUMWf0COQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Of+htpAL7TxZgOfvS0pgoQzX0ymCovnOmoI1rnPvcenq7Y19zYsNlG9KKPcuI+JEx3OnOrmJOijz
uCtrSL2Gl1m5deQOv00IGzsJq1O8h8sDzfNoSBB60BgQWZFjqyZRdNYI52ud0wCo/7KpuyZkpee8
AKeK0WwWJq//SenFhLI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eoC3vGHEuICK4U4bYm4blG0o5RnhfwoMq5D5oRD61vWMky2mOvLilS6/NlB+XaF+FsK4OSIQHeMm
k3VzI8BaRu9xLPzGzM4c+2xFQ3R0X4t+gMl4u6oYV3WkRtFzn3rPyA4qXDLRiCIkM/aSjIliGcSq
mDBaP4MeLDg9Lg7WKY9voHFu08GknDwNDPepYSqrWojrX1eJ9hWDddQW3HgWinBxHQsNghMpSJUK
hqxOcswDyV8g2ZUfkU3c3NPeY6g7jhVbZQH/K8rILqX5CXbZbSACktgMqDMD+VIE4LLQ/9xWXcxs
KYLqBnbhSjXJcMk0IoP2NL8UVE+8dgKkYsWaEA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54896)
`protect data_block
9tUAPRZtaSkHHJWZidt58QIZ1dKs2XH1YyTCVWITPrGEXyeLPia1uUoUaeCVK0Q9In43uzmc/xWR
1qwdVqBxv3E1LicS0/DFeczVQGatXpWmMyd59PyvUnYuMK/EONJd8POk9JDDSKgVrUVfLIV2t3C/
iF/Qzb3/AADdh6EpHiR25G3LtVNUPc0o9M2/ZtxFB+/RxezeNYV0TehZQTiROjzcBypbf9a3C3n1
uClSw+fC3H/7UWzNCpPtQR9R5VJj7tYnJQ+yKWVX0TmtCG+nat0X6jeFFcxye0H+U5peEIL/2sGS
LuW6yrA/QpeXMw3wZMrIBfHp0E5OZycYndjOO8ojhZkCsmSB0yRCwoU08Us4ErZj/R80LbVFiXLy
oolDstw9gdYIKj22r4RVI1Jom1QFkI3Mvd0BNBHsChlc6VMveSUBW4Zmh8hOjFmpzwU1QqSOwVvH
ATcvVGPPRaMdom3ckyiPcbxr+dF38bmJtz8JGZ0IvYZwx7mADFUjaaDhSO61SoZsd96XfOOwTWjb
w0pKNTdMcfOx5+bfNUlGtYUzxhccbnyM2RL3ufg3aXHHXXiXi2UlvA2Fs+UYxkspeyquFw+JsCNS
h/T6kGcPr760rrv9bjjFpUY82YGBJT7OzaK+Vo9v7vDKIqe6b8zd7PAN/MrZa+0i/zHGmLfGeSFN
E1LuvOIeIQQBXc1f7o/wI/i52fWTWca6gYe670565QulrSu3qx6nBvj8e3CyW/ie2HHmTbvWfHDM
eDRK5n8lmGIZcdJgM6VI6SfckxRU1d12bCcmcMSl8Y9ksnELGrGXFVTcNDhNkMyJZ1sYZGhALwxH
EMFwEQtos41vdZNxc/8VZ4Aff5PMXy6RpUyp3DpghgufpoAfor23S1tfewlFWzyfpMIeEItRUYik
oVsBVEsa3vj5o4ivPhnNMjj+QsFBAKi+/AF5Q5dcfwBS+oDghXV4Zqn5dtDkRJfdrAqpS2gPYq0z
HGYdB7MNH3adNEkCXMvDoWPQ6shMM+vKBRBVFz3yhBbFoFNwesKUHrIJ5EGxeD7cLE72W1mQW8o1
cCP3/+J4pj/pGSceGTLREpaIYckkUGO0vahMXVr7Esks0nQe7FG0MMQH+QzuNfzyqKZlScOuhAWJ
Rvx4K2jtaE0mBLJ00/J51/wBKVkCjZyMjqYw6aS5xEYKthihsdcZAuhugw89C7rmmZTEvOwIUano
5cW+QZiCe18G4tTDdq25Qx5+iaUfH2VWWneBXLFDngwMQsYJgemV7XIsR1+9NKujEZsrLWi0cSPR
msTG6rmqbTWIk180oXghpngwEaf3DV33kIo9eODNKOqL/Y0ujj7uUATxXYOXoxfu+QaPtYufLFyL
MPVtgGYTH5Yqqynufj4gTmo+OUyigsnw6YbF3+oYE0Irx8Sox2lc6GrS3kg8e/QyRF6n5mX8/Kt9
3QICkgqOKRy0xfVRNJCDwbsd4rvJyNBJQwWBrQWps01URvfwN1dx1L+YsUQQDNMR4idPd/RQL9yL
FpnWZnL+rV8xPZ5YlGmddRi7dqHk+M6PEHRyehn/ZyBtn1FyaCXfB/yc4YQkao22q9KnB0/tpzJR
gk8iJHjN6D6ySFaED2kGIVT2Dm7Ax54QNuXtyzD0YhPOWcNTtvGXVtF/DdY5gnMdrW8FxVO//j5w
uoAo9atu18vKux7gxbwzMsv74CePjreGToJzRglzXV+SlM86YYyA3hDGN1WS5GCigzNKQ6OnZbY4
y2nKQlctIGAEmR40fJc4X6PEvuyucLpXchNouc+wnhfAl1n17gdcOU/1PyL+Sfz8tGKgBf2JN79E
bymLC45zRYAdT5PL4q2eaoZZjPtPBz5Ds+wocAG6i4GK7ysBixauZgW0Y6hYiAqa9/TdUqwpPsyq
ZkeHPPQ4Sz1E/50NwJuN56FTZg7yVvcvK4rlQM9VvOq9Thuj3kT0TVAYkUKbLTAiblZxamDmu9vp
1no9xQNqDsoB2/PjJQWlHJWgkfCBgeTtL7Dxibtgb/eZDRMX4x0R1Adh3szCucF8OjAvPQ7vQkvu
/xsTjojmG50KNhv/emqt4uQPiieX7EfzvvIn8aQ8TBke3Lau0n4CbuEMoGl/5nxEPHqHc/t2U7As
dwBby03C0PLm/kH6vDoIMn5CfOCQRsEhHAop8C/DKbuezsgADXeilIXXUorjpzxLRsSn0CjgHLZ1
QVDQJ1rDuNeLmmWXb4lN+2799Xq+KTet4RFW9EuAK4RRRM0mIjyYahfgSueFKiu2UKozrX3NWFG1
gZLqR0DNEFkCfoSXnaascEuShgGDiIZhoGCfmU1BW9cxhsfTOJp0K+qzIcVyXdDi5XQTwP3aFilN
BZexH9Ea8mJQtQ+jerb7efGyyJzYXPszIH6e6KXktTb5Gb50ySGr+ZB8HJ4IJuvLIqzOz7tw/0Rz
fQ4Je48Gj15QWeY1ZzCSyUonlqLsuBSduqFXkE02clo8M5rJ4aPkprDvSm4wk89QkHQUAAeE/q7r
zW7g99uc0HOmkvEnmUxy5C7+wdNlTQsyTEC/9ixTWkAIPl84K7ZPxpyY75d/xwPTjXbl2bgaYvTw
XCH/covlhM23+qPs/7PWrJs5b02ua3FhUoWvc5JY31R0fhGovMcWa2LWFC9NTwsD6GKMZt28p9+W
ce7eJ6ghVzz+IBBZv4Eu/rm8fk0U5UOgSDCPbtl6NM5fJScFRr2xQJkrUs4U+gNgwj9xanRcCq4z
ho6IyO6CivsSZEUxlt5Ot22pYsI6y8GdMoLNAuhjQ1Oycp+Bfur0vIG2U6DqWcZpdqmOxrztrQg0
QQhsOHXYU2CGkE0eM4JTBNWP+sdH7541NeSYyuUTyDwnQ/8w7uW3rPaJ86QxFNpNwIdAHivTGvNa
ax4L8NoRedbfg8hdU37q76AARLIUcXYHrfWVrTX9pSOMObLv/mAm/EcM2maavyXjDh1Ouf+XTIiC
xyz5k74mm/jtZZiEYOmaapZjiAdHOFTEXJy/HNZ6dad6ZqpeII/IS9qCaeAQjP/UfFWpjhBmENKg
7kU6mDyDVd2CMhOnhVGg/b5tEN/X2G7k+l4kTEBMVPhpQWNP5sBBTBTHwKIxtqoYxkgNxDH/0gzi
QLBB42jMwei5/5rB83cXGw1i/TUUlRM/3Cb23vEGiN/zYKPVHPnkEucPcevZDkFJ2UgRPYC7+0CC
CfyqVLNPCmNvKRIKHQOoGKuIQibWJQDODkFG/2G0eWObiIcxk6gVWBATC7LQArcVdWvcMmbLseSx
b2Py0yZJEy1ZC77yagMnWciMLEukTbUnQdOlHUee8lwIezU+Dslk0T46cAXc/zuLRN1G1cpcwrv5
64RjdWvye1Uv8awS+LZF/LabWMbD1Q14lAmvISLZdFgUzAcehhVDGVx/1lst1hKie+DOdyXnW7ui
8AiMIpCEKYfQbh7hcuEjZAdx3D9euKZj8y2T9p3ugAf9rgOv3H0nn6jOLpE/WBlMb7UJX3RfYRD7
LoYavJsnKxVs3nVTB+A7SSUsNXkdsUTIChF4PMbzyNHr/TQWNrF/SLSuN/8KBe+NZFTIQiH39U4n
RQGwuiwU6ql7waZBGwm1MZ0G4RH6FEIHCLziBP+E11IT8vsedRZXQpNB+MiqTkNUpvJW1Fg53w4K
yX5BC7IC5lQuDSLd//Uk2SXl8c0BvhzfedT7Imnqn0EMO/25Yb9lnxMfkH5xGg0XShAwsl3f2/Ns
6Ni05M52QcHAeSEG5nQRi9Aa7n44yPGfalmEdXbanaOfCFFOULgCsYTd4DCKDd65CHPfzGGnbrOI
6fG2hGnCaZAZMugw8enwf3pP4g8P0iIgxzBP9dNpYVXcoRQFFw5o6hZoSH1k+9f0ruv78uO6kUW9
rmImIvbszFuKD60Q+SBn9Jup4wHUcoyTSVLkeA6b4Mt68lAxcT7hHWFnlqvUWdACKR8hT+U29YqS
yiPDZh9TS5XVvuCY+Xj/XOrqjyQHTyFeewu01SBSSx8aEY1rB3UcOTpHAgsDiS9//RuP19jOVsFz
wtxTv8jZrr3VjpnetmSfg+PoK9yB0D5iS9urZ/RZ5fVgA2kpHNgOP0Z26ZyeV6duC9uiEtzx1P+U
xhoGWIuZhV1tct48d1w+UApxwVjgH/5pii3bF4dzXPq4hcHjkhSRYTubJ7z79pylsGQg/eKVi/R6
ezyLB467jWpC4s931JAimj3jRbUKlci2pHsHN+1WbX53SQVEnbv11eNPKF5Cm1Khl1l3ZcKTdFnW
1//dBu7NsG3+mhXiK+Vu7CvrrERMXKpgeTrY2Eyf3CtJHi3Sx7dP4SuUKqGpAI/maHOvHcgZphTN
l15xp5Zgd5YVqLxp7h6b/+cefg4rzV1cXLeuFwB/3tMAYR8IeBRD1/m0q4gIiIbbu4l0v46eyHwu
WTR3/tAHzAaSOTriYYiRGg+9+7osMMTA0gXkkAtAS9ZJhm7eg81/TqBWvHc3tDNtOzp+B44lQyAX
TJqqO27zUB8o/gdm0SVHt9dCli1rr7tIib8dTzX5WHY35WuQk7YBWjgKQ1w2IRPtU+RVeyeTEzE2
tbFO5qk1PftVa48xa05f764PK0oVTuuwmU7xy3Wv6nAF5cdyxnEWBJHnWt66XdPTiTB0t5GdNlyV
u/CzYXUEjQq/ZSKtk6uLrXeV4jS+4+5n9LZm9+a4eqqRW2oV+lSG5MQAAyTQk1hryH8wCQhQERga
YPrSkCHv9FZLo+ZWvBTnoUf3zDsOnq4/Fa280kEozfAySvaLfFbHIh80NLwE5ZxTnztyy0Vy4r3o
5ON7lS43TB12QJkoksb4yGlqhcniQcPFPfGVTb9G25YnCpnCxkOGtLre6loGeEgy7lrul+6LbPPO
LkUdAJU4qhrty6qzOoZ2GnoJ3Umz0JmH67WrGlwwuF11sT1HUev8JrQF4Q6kyEFi5jq43tgJRW/7
kMDS4GpU9PfgY5hJ4LpvWJzLY2rH/QskuK3LN6wBTQoNyvDz22or+lionMBva82PnsjYct/Oeqxv
bPwyC5xzooY3/eZ1TiPzA9gIBha73yvs79fpX+Ps0urlhgbS0yvJnOB3cEW8zf5NgpSw69vvACcI
2/SH7DRxNJ3IVv01yl/1UtHMllcXD/1FwQGofp68GJlIf7zfhLit31IiUO3XhY2vKtwhKbc9r5D7
abZmjOqCBynCDvhh6JDAJ54lPJSAQd85WCHa0phfcVJpJ2E+zY2zVaHiHVUeHt2ygWov/vOZFrf1
M6uQNDYlK8sLsD1yDjgzu14RN0s1LmGxfM4ay+lpiVAUsrOmccdo1No6RbohnohkKG3NthQlsiA5
zj72hNGVF/HOm9hRVAkycQ3IvhbK+2QcYkF/RwZkj1TyDPWBAZ0ELu4qaN6zDeW+gxru0IJ81h20
IASOLAcpWqO4sR0Sv7MlpKj2gXVWznmE+OPk/fU9hEccmDx8CrrJMLtJRARH0pgy8n1AlNDcbFwL
oqjzl5mYkuVV2KijiI+YJuN/SiiiIFp6l4MAIgX/tz7GHwdejV5DoK88d9VhRnLH+8Gg5w9qClPc
LK/lzegbwjvd1kr775GXNAxAd/T1+4qA8YcfnNDecBK0fljFO38eMzTbyQC4PkHCCp12F+bdxjnF
3q4LSvIuNNfMXjpoYLQyJUkuMiQMBd2G0SHJguFPjsfNVHGAMiDDFpqWD1hSXkWXEeCjAUelK1Dr
Ys/D9O8QBnjjl3pmdVeO4aQpoxYKfyeRAJKZxH409VZh1uzOa+45q/OIT/mF9BWBF0uxmCImU7w3
wS5BDq8z6KsQE8SVWtP6WdNUSk6P/1KGfRHub/3036CMraw0eJekQSLWyHZuQCY4rjr/MJ4EFLOO
2DwvXH/sb8mVpXZWLrt2K3icv47cP+F/RS0UMchW2SF/XPr7d1Fz9bzwj3IrkVl4v8zGlai9Pb4V
ToyTuygCxmddm8HXKzlHDh5uOM+2Q8JFEt5vcR3k+zyp+9Lphh9uCmIFAzKAH/JAOk0XrI0Etdih
HbU6dKgJ5p9Cq1VjP6n0cq5QaEvqPW/zoH5NTTNFl8ZAhNFDrTanibw0877y3QkQkyXu8XfDVgOn
rmTKDDHdhh+FCYoYv6zK9Wgx7Z5a9EKZZNOvgucbUz2MmwViPBWarXACQ7nk7zBZvrQWc3mqXk7J
ZUkWjShDPv47isFlLlTQoiAbt6+b2JQCM6Q7DGA/nfjB2ocVVSbDgX5G25tfx8ULHuAmhg2tx58G
qK7ZkCUgSw8x7yWdFq6aQ63KynqMqXKi7/8LcG/I/Ju7zPD/a32Lq8M/EEcs/i634Zg70O+CApwX
DM6S4hTbH9Ps966OJ/fUHDabJKhtEzzOomNY8BmYJqP28qN+PvlHlLRC86zFHWzdvvt3tHaAditM
5iAuZiUEyfaLN70gG+I7/E4OehFc0ySyN6riMWHSO1HVDBZtPvQm/cL9sSZSFuEGXAtI5k+0fxuS
Bl625KWrb1EAxnDKD1Y5mRnrdYmBUs8zIH1Dk1WZQ15oVSsypT+GMWBkvWV7yqL7z171Cwl9otkM
x1+M7xIeJoflkSpfEPikG9dHAKttczN4DuLOmQrRVHil8MboRtZ4KUu62hQCHb67h8yIs3MHO67u
My3maK+UJevE2cUqckpHkxSPAat0kQQ8X9MF1MASlrrB0TespwwpZct59pCsZK2hYC9/ACEaEl3z
jiTjPPDfkWIDzT17D2g0rT3B9Vz2qlVFNyRcW5Mpg4HEmeRPHxChPnc7m8LVvXc4xeVzAN8fk89j
xZhTZqpYQKSIDYJ64fsTibHXSc1Cnk++8md9rdoY3u5+2QH5jchNfc0H+dO4aP1InswwJ/moRO/E
fCXfETZJxiK6QD4DleusNqfD4VXHMh1OFFrFI6yOOmM+r0FhQjNG6ZI54gNvBcRJxaK1H9j/ffa1
n4coaLk3y8YI49qcwWVLbCWy20d4drnMv1NWQtMsBR4Es/G4MxMRLu60/UlAI/DIqc4sWSBq8k86
I3yNzD/SCvIpG95FCY2ynM12kwVEtrMbqAT4rw07L6DZxwaCv/V5z3B/h3gvo7SJI5W9JlUbJ8FY
7o5Lox/TKWqJQiQJ4Nae2EbFw1apz2YJzAMibHTt07VKRWCXjhqsyngJGiWubn4kxQq7hFL9i+Ys
Q5G63/3n2Q8RHf96W1IWCa5MhFHiQ8IaRrR4QIDq3FsHwQYE9bbY/JLfIbxk44R72hhtZsxILHU4
0nda7MPMAvQvEs3tdhfRH/KA1k8S24Erfk6zFj9jLfrPyO6cAorknbQcP2kVJR0MNREQVuYuJpQ4
9+hoDLgRZ1WWxa73O5m4Iz3GX0Q2mgG3QYiELkKzVRW1+K2LIg8R+p01FWkIFjeonuT7umgBan3D
rEFhkzAZwFi5udh6RUMbEV1ezuEdopdeMEDvHs9Dgr0jQf8gdV/X/KKb5mZ6Wqi+HMGfaZzXMNLO
OOhMI/cs50rWx5KN2DDRURB3jP4Zi/BDeNFBrr8oNCz7qW60yYRZ8DYVQQfTVMkhWGKVV0zaNqOJ
CHrLtwKlbRd67UpNgS34DKCuarvX8NxmlHSEp3IxtozAe5Q8Lmo+Niy0vRkIacZEBPDIkBUBu3w8
9mVNxQBW11aBO1JaLB6w8tHOgA1flkkYu7p8TiEthKD+mwGC/EmdZMZOSOsGVCfWJgFS6ZEGKcBo
LJ8lV7c4dgT+neZi5mqGKYCCobdajiCKq8xYtyCXwiSu5kG94WwwelztJ0PyaMPD962RbQOAHLce
TCcHEmm1fLmQwfEzxlJfGv4OsLMFy7FaoMKD6WdPcUcyFMOq23Z/mmAqdGjHMvwR1hD70dOUGm9M
BBilEMCwGVPz4Nq0OrhbTgVQiS8wQqfWSY/trJN5jxhCXqJ5j7wT5zrfMH7TKxa5VEAnZpV69Qse
ZCCviwYKihHsvoUYdHTMeIYWIfRhaDEaufaBo7nFl15MGuEPM1Ak2i1XM8pp824bxuvJgt5ybRJ2
d9gdQfQz+a7MKlubpreuB0XYHOsQ6lAeoIetwk5ucM9ubV2TIWLhwC0+RP0O4RonADJoa8D8g0wM
ay/XoZDiWlWR2x/8I1hXexM4Rlkx61Di6bUWI0oM9L0unOvHHdFxbeMJtRXoHnN7gM0TLy9+WQ09
StPVelw2WHQlE/e2GAaJNFnWyIwMQKoxTSZ8WxPfuIq0KklZ8L6foFwDcPXqn3I1XV89b+ur/Yoo
B0lvVYsGaBq35jiLdOTk0fAgYTia2VByQiwRpIGI2QwB7f5Bx6tbUubMIhWypzAqZZQGgpsPp4b/
Xzs7crtiGU5RHXiWfiPcvwkeaJxP03NQJBBTUS/KQ6+fy1w8F5P4M+2JMjVTnizS6bHKhZsunkHV
7PCEHz8U+EHIYuAMLsiazWpBiu8vxkwomI+cUO7G1KM7EwGCcSuvmt8S5GZnSTeWjcEHDk5Jg3SY
vIPgHC0Vhvmrbo5X5F7xgngtRaNuhMjuZWTr8v3uejE5UaoRU7b1M7d4wysmtucGOMpoMtEi4pRh
OWMKu1RLKC7cbUrtSVQ2Y/wgWQ1n/hCFrHN1JKpEPbUTbq0kQBpy3ar/aSK7zwJL4mQ23aHm8+j9
9jAv+XrAk8NsmsXOqTQlS30exSRlsSUJIqy7TFNrG3HsmKrcpmqSDMtf4axjENZ0lDXfK48Ob8DJ
d5AUC+7EInCVkYEY1mpJ4U7zNUFHPp5O2G79HeB11YWJpwK+qg+Uhc1PpBX41/Q3odyv4vUI7ckC
YfsAUosXbwjk0grmjayx3Mrh6/XMXT65Y/MN1/7E756kLpIMxTzGgfrpZT1H1ttjHrUiXZ589Psl
gN1gZGTS8gZonTuMcS5y8nHIbXa6fL1aOADVy9hjoefEUgQnWnIXL4oW3Kj0Ir5qfKftqOoazbbK
BCjUfDA5U1gwmYaO2UOot2B6hm7BX18R8J8kgWXAMZJbkfoWb7GETUAGLz7tZFHSbNzMJTTj3qXa
wY0hJ98RL2kYeWY3Cfb4z9RUyfzXQk+8ANltwTRVqupSH2rCrLjwFpN0Yru4eXtprNJIGSFdEt0t
1w2zbgatwbbQdGTJygbiEFCdrbGa3oW6+IpmO92Nsr/ApeK9x0U37mMIAe3xGBQL70j7EIj1Ak40
pEkc/A5rStvnLabIVRK9xQW/dLf4FLOK2FinfDmwY1LuLKzkSHR/oFqVsuV3Iu5GVxsGx1U24cux
veqAcsTllEEAgntPftZnXFcvByBzlNOEG8luUVsSHS0L48YrPyZ1dMQ0V40lQ8LoZD40mSeVjuXB
CyBoiCB4KnpRJKD0M8W8ByygyuzZu5XxkPh7cZG6mSd5SRyYV2/YGUhxixORageR1zfHsMguyPR5
JqFMrzNG/HddlK9WI7rI+rQaWuoFDoSiRRhDnxJkZVIf8ePyGEf1xFe8MrNmB7CE3ogjsI+zUSBb
E8WyCPD3RVuSQthLZhe/igt2fwAEKXiRBsomrsXMiZWnkug2WSSsfdfY7nFlli/r3bPAZmjLwsl3
KswegPewE1TTQTF9caJSMfAJKhnlhEDQyEVb/FDH0j90F6OCYCWemNvCd8R1p4u/sTFI4D0Gpw0C
iKl98tHAyFNfX9xp2mKr5YZgnfFtM02GpIpJ3KE7F/MYmOcu/SqeqSQ/lWhVKdqepRhVHHbFRcQY
Xdq3APVo3AADJNSK5LMF/ztnu6zBcfRyPugFJd7kOT373DM1ML7sBqOTYbHvQC07F4/kvnZ5UA+K
zHssViExbTBIc748xMHfIDUd3PpOMKik/nZFQNn9NYWpDpNzWF1u5jmYv1HA8Tl+BrORdtVlgo74
oNGGD40Hd5mMI8VgROxEd35zIZs81EYrXiRmWILKiU1hb+h6EY7czyPBFdEkoVWVnQ4mjuA9VCaX
lHazSBbsNA3AKGY56d2OJZpNZIYKg5OclbzSVjxNIXrSyQ+xpdPm+86d2alNShj5evrnXaTewAM8
jzyQ4CQFHgJDndcqpQYq7Kaywr0UPvHOMZ3ylbXbqQiiovzhYWL6TEiqTMP0Cm9qarNM+ykE9Itl
GLkIuLk1FeiiJ2/N1ATrX7FwqIKabyiLhA5LzLhccH49STwD2l9N7d1Stn5BkfHaURrEGjxUCm0f
JZPaNs+LWrCPT6HV4Qq0UcUkXc0+KZffwSGFMzgv+C08PXglWVZn51YWeLNM5A9J0nJnEH0Kz1vQ
4eb4/G+d6wgYR4mHRPJRQm9Zv5HBGwOTtfNSnexiHI5y1xViNJJqaNhPp5tPjodsR7ukGvVNnmrk
1T+ZsKMEk9unolzey0DpNAdwhfpiy3h5a3bzA1ifWTgGoz0OiMvHEBMOqviDhao5I6mR6unxKbhB
YNCo/BMJcaTJUHYt1DthdqAXjWkg4sRg1NxgXwFfIUxc49JLhoPMVtIoKc5by25ZwkwVIercRjE2
LmgJljrZE0AnZnObKU03ykdiDN8KwmW6LB+hHbv4VjfBB+28wzEHiMXGvkF8lWKhp7xlxPT66Y5p
xfTsZvI5PELku8N0kCiVPgSpSh8wIIZvkvF4rJWB/ImyENwTpX47+Z5X3W0jQ+ioHPUYUJY9Kdwr
uOqm+tDLKYGwXH9q2olxTwemlW3U3BzvlmhXlBuOn4Pr6WQ1mU5DU36evKuYTe+a6qWA7qCQpR1W
J2iYNqtHz35sdOSmiA32ZPNOH2MsikLaFrjtdeZ7VO/u0CVadUXK/XHusCgBpGfSAKAJYYtxSfxV
irj6I+/Gf0b7I2q5SLjond1eW9G48rBBzo70+te0kUD+Zn8eZM1js+5jqBPvhUb7ghAQWsxhq/aB
dwoddKsydiwM74c5PyeSvLKb8Y7xOVdmqAAyQDNgJzK2BLwrgL0pvSjSF0ZpbWmvwqbo+zRMNWzR
D4/xIOZuopOqYUXi3fYLV8J0Q4Ak86Fl1xLgUTepE4gpLFF5YMJKnTI3WJJ7PjlCpHoy5D/GKojx
RRMokqV+e/znH0KptqFhf8bNYca7q0Fh8/C08OpLyg2y0OT9QaPIakUxwoPLXWgvZ1Xb9BdMmss2
RJvh/honUn077piwGGlUj8RbQJovFMg5j2PnNhcT7RqWiIQr12C7y2nh2xAI6jwutekvGUnpxT3N
M+anWC6o54xfOwIdCM2SnSI+toraI1tZaFP7AYBc8QkMw3r9BJzZmiYLVArBxmLOBTHXX/bDZDKR
azx5t4md6hntbAJtLwB57WJOfXekOlFsXIAkyAyQxDHc1qLW9AfeX0aTojNRaQds6++SdX0XlnOe
RsByYSt/LCMrSYEWXoJvP6OCT2EDpdHOHk04k8jAVqqxJVvge7TU4TM/LNL/JKNFlXrcwpW64kQ8
7DOev6PMcd59cm6r2e/GQ7V8qm89jda/qdcKCCfdCX9Pcpv8Bcqg7ALv0i0K6Xb2fMp7G8Wu1qE0
yjOrMy/cF6SUNqmPcw709SotflnfECAAaYhHdzBgtLLwyol8EphUmy3fkbbGM3g3wOIrI2H88tqq
u//41pXVdJifbWt9V+gVIhiHQ7/chlyKUOX1r8BPaIs6waYwG0UwLv4vrhbcqRuY7gCS+KVvkDmd
eMyG9/JM4B3Tjjq6n5YYUYaKckRoAxkT5JABzeBgT//J4CIjpLck/QUY+KyRVKehPCI4jZWkEykX
lIYGUnNZj55Bp6NISAQGsc6abbveRbMV+ysH99op2+RbDZqdbK+SASdynPBd1O8c2movTtYYXR/D
qeAVGNcPb3FrXJLn/1f4jzNucKGLOdQmFpNipskrhaEUsAlr11rmo4bM2lhHp9dnrW6Modi1cTaw
QSSrMYVBbx+XVNCmX2dqf/PBHeCt8mW6cytlwJ9rW7aI9U586th7IzbGLvpp6K5l8ZG/PRutHyqK
CWf2zxWYiBe9VRe9Xe0DIl1K91SUrr7LdkmpRe+YmkX6hqk4oUVW7Miqtbtm7F12F780EptcJ5O/
K5LEJFktJw6tgzcilYd/5Dy+CC5KxjRT07+MXnmrunX8zeJ0VvN0s1rB2tx1FFA/AVPvyb0xyeXe
jDXW45/AQ4uqpWZKMqCiBoLK4GDIT4Gi6QaXOK2BfooSXwHRDUty6jRjh1pW5TzQ5rBaQBL9xBQO
QyqYECQC6TP60WpHxhnt5gHovJ9ccuP78pY+erJsQWTeaL5JtXb7U0yjIiqemNO1sh8M535OcaSI
0ps5uJVbn5Kfk9du4YpDOw10TH+bC7AzsllqNo0KHILGPoOlhYe/kIhTfSZzV92hbibQuRMNH24r
K1458crW+Wug/i19q9bFx6Nsi2lI4PsRuRzvjvwWOXvSq4M9i+ZnDJCQNQCE0HF3Tve2NyVp+4o/
yBtB83KoeXSdIc9dgjHASiFt6wQbFwLdic3f9TzbpOBrVNFXqNIV/zaXBzDd7A+QRY4DbKDvpMR4
T0KK079rFia4efrzhdyHsFVsHSQ4Cl0LRq9YAmZjJChB+e2sLnTh3j9bK8O67UxKe6YTwekPI7GP
ZqoQKmMX6mQOAZ+DI8bXEI1gdSSJa5luMQIbtiArh7jfkyGGBYedNnv0SbuqkwdI0AjNZX/zJhrR
e8duTY84UFI0QXUdzqqdq/hFZgNogSIrkbIGjP19cGU64bBklRywrRSQt+68A8Dh7QtPPbT8/71S
qwvZ4FlsfgZ5Yj852YYdkwQ66FrX6PeKa4JmDhub4jcMTbgXLBidg5rjs0ObhfaUbSBaGkeYudLV
0RFGvwR78j/8PhEeX+4J9+XVDl9TCMqnwVYGfBdo1Di/Te0Pu2NDTzujvk00qmQWpArba5pbB8BU
7naXO5bPnfMgCJTXv70rI4PEbgZ6/I8VdYMUdu94WWqCKRzYXZ3cXmElrlGBlKgfZPF8we/3Kto/
DBW56lcUn4y/FOE2e8JQMKQyWq69OC2SX39EgV2CcE/XDxjSn//gfD4/XrRgevn2KHzETEqimbux
UhFyXBhmJRN1Jy9sWqG8F4iLz5/4kSapDFX8q7FCGZPn3DGKbUunfSYtg8KslrGuc0WxaJUFb9Yg
LOLJ3WqLo1MaahdW1HIKEBAFT29d8woU46pS2LXip8g9qJTYDu0D3ijgy+jIvxtrian6qXax2BIN
Z8ihztn3mO5WVjweIhdErttUDV202Wrx5RcAOiRo4GTQFbpmxnE7RJ/+CmnKRZZblmcbAPJFdC2r
SE5cZgdKxmTWJSr+760Pk8zS7cXaqjcSnA8ORjZxvvL2D5YGzdGcVmPO3E+E24ZV9v/If2u+virv
K1JCaEWd2uCiSoYxFy4WHffWa8ahsOT4k4ztumjiJz3TqCE9i4apOIw9gd9A6G/+7CwUYkOocpyr
C2uE2iBw7UtxzGFJpk8G4mRHbMp/wXGl0Ph4yd79uOth9+kpjC2n8M1hOMAHHuuKszKuoooKpfW3
nvORPAAlfjNvE2O6yfKfWmsWfgaLyyvo8AoE6eLXbdhvD3wvBuY1quur4VNcsIyppDH4d/btwxMF
FBmWCBr9SmZC1/LwVcP2ADFcXoEqcTd6vtx4APYDK84pssWGFgMt2gdvl4lNWsjJc7ywOrqr8aNB
YW9YM5m98PvFrjjmRTrfL/VQueTetD1cPrBV7G2YDtyROs8GCukOg6n97qJqk3vhwhOclnn8Bnu9
uS/DipM40f7onIOtTuQCwI2X+TdybnKyDrE7rOlymQEAWxUW1/HkiR8y9ugUOxEIhXrFZ8gS5JXM
GbGHftK4VJLhpn9O/1fLWHZYPR8OtKHM7mL/W1ntCyTT1yw69OlejjWpOvQvvvWump+c8uz3O7nP
bbY9IpvBhhaD1+cFiSRckihiJdqumhyUE2ZZ1SAmpmXn/Jm7/Wr0RWYOHM+4AMZVx5KHqbey7PI7
C1S0Hukaah4x/QEeUNOr8Hu1HbFQXdO+nH2LKhYE0cZJOTZ6mLC/COlYtt8KjJRrVWpV1MuvHpn8
30EEX8XpWPnu/oToj7flHkXibhszBfGRa4rCIYVh+uPUbBhCRJ14wqqjJiS6wjvoG2jdJ2KpOeHR
CFP/OVoIW3Aip3A+GHAPX8kZFW5dILilmaar5Vz8jp0f3+1fqcGBdmaGgxyvuKWyxkcxJRkEa+1n
9AdODMKlFkrkGJ5WkWHtAPTvplcybb1e5930LrD6sFoQb7qFL8AAKQjvLFIqXn5uiUQPL4elDpmt
PcuMhv6bDxlLJeYI4Y01FyWgMBjYdZP7T/xxHvM0Y20p+1yvOnkf8NZ4IsZAm5CI5qIMswGNqpem
vabcbEs777rHopL+v47Ic1gmdm8iE02nzzBuns+gjF63EYUGHZw8rEdYbdIOo5bt0UBzreKZSGag
/AWGSiiJPQvHf4TXGR/7FSOZ4uzYXQqFIUzaBIB7BrlU878tgqYxXbRBthYoV5vec7uGTSYKoSOd
iNYsK35SuFFDzZxargVbNp7sZmaTvV1lX0WpJRBsXkdjaA/qO48XHAK41rw1ceU3YwvN6zoTNnOV
ruyAkPFAEUMcmRBS6+va8lJ+4DCeV2pQecIcidFmWiOJAM9iedEpEShS+1Pjcu3IzFDnbXL3hopZ
PVNgO5SShFX17CWCX3TtYKM+GSK5s3K0Qvr7AV50d5k2u0YL8P+3/EAeZzuOHJoaAhqk2amQqQfC
a2cqcLgKGS2fV2OUelxw2/3PNtN3WPMHS0MWR3QNK0utpfUw42AvFdcaogm6BCz1owA0sPe9tDF9
v3ZCunZGYgMoY/Ip80Ku5qXHt+is06jJ1AZ7/crYkL+iIcNRozLjxc0G9BowIGaUSMMwxTIx7cwO
mFqzCzkSWxlAVWrg1lsrsqNiJNIDXjkc4oJSx0Sua1mpv3NQjziZ/P9pIm6Te0PyRc8um9dzjw2p
2vnD9rqaEL1H0d0FYP/52tabKu84SL2VoVBeYsOaw9bxAbRWh1iIwSHGikbItbuG80yCKm7uPjNN
C4c1fXEbDM4wrkZpoiRm1vUuTC5V6zKimSk0kOj1g4bis8sldZsSlzqJXJWl80APNmlfFxCcR3/N
QLhrcc/ShpW+p4OxYnCpZzmp9UpBDu+RgErGjrqUu/W0sP6GPsZ1MsbXABJC23jI5oRkgRPNNKBd
hoJbxD8TxmRPb9tOQGtOg6kQDNKE6rkafmMGtPppo6rKYy3+KwH6KLo9IjTWlCZ4dO02lbh6uLJM
uLPnt/6Lg5XLIp/0hLYIf38Q7NWsyWNQfuah6KZKG5nxBThoG3DXIz72APm0LNcJAEVsYMjvdatP
xWUTBpXEKBoV9Gp5bHOJgXpFQvU291osSc9GIRImBuJgqRSDE975WJkWE5ShKZf0h9FPlOg4Qitw
QM1Jy61VwqoayDK5jPBXXPuQxI3HGKH7jC62tFHTmv9ckmCVNQUO+kpM/6zh2wLvj1+psfLwbE//
dEYBrZf0VXs0eywy+PUD/i5Y8uikWiyHk3aQXnQtyCPBUsF8roLs+PZFLY/+FDSJVOGY6F/Oba+Q
nLIWtOth6kc229wrM+LWwqkh2hXDAosJS+xSd2AjgKRMMTHeDBO+kaSMIK5/aC4vIfZtHIYK5DQE
JIfGfFyRJWrGljyJvjMdFJCA5kX3ZLgywBJL5kSkdxgTmscalpREmB1eMxj5e+VuXf8StJhZ7DyG
fIDfXXp4SBw/3QwNviaE4zLWV2u9+vLR8DWyKMu7gSmCo9iG1jLx8oBxsxRWVFzSLAPgJ2UkYGkY
vw6W4eBjp8jfnZn4++GTAFYBsZc10ZOy/zANPAzRwk8QTixeFp1lz3/joUm8QsOj1YRkouOpp2k5
mlB8d9BRQ0IQ0eaYyWSN08qTtjRfaMIiYggE1Y0CsWfgmxg//xQlRCgvkQwgTtlto+I8V/g3fP8A
s4Ahhy5HJWP5yDh03VQbovGG7UMwRAr3k7mI95NkU+g8PeYRO6amVUCLo8vsKogvpZmCl6wnQpN+
yI2vfJ1L19qM0zJkivHpA/u1Y1DXuRKRpf/3dkal99Pw6BammKCOP2iVKtIZKhN+iXo0iZLyDalY
YJPaVKbbTLC2eLw5AIGej9Rx0sF6L0IUngL2KP7Ax00I23Np4Mfh5ZLCVWaFjmOav8vlnWk/4XIW
AUntKhF8TKyM9iOLTuz7UC3ajTeaJWBzKvQWO3XZcsygXaG6n2VnpZ4qd8IZCHSA/62jpFFrD7lA
EZ7TTxXqYaR3VuXXTsRCcYS/b1BOyZGpb0EhfpcCnKLT8s3m8iFVLlBq7CpqW5zFwPxN+qVU9xbd
izGQmVJSsFRpXbtDxsqDLDb1CoEqRP56ogyU/GaqoGuC+6wsRHDgOBVp+Fp9Pku8b8+IAp6iJBZ/
YE3uB3nyaywXkMdxmVhDOszSB7mqpshMiXhbJHbrwapfdOh1LLaRSd1jBZM4xFDehvlbFuoLTsGK
n+x0hRHzeW8LFCGTuLtBbtXhAUF66gcyTmGET1qZq5YypxCL+8FjRRJB5JgDv9IEOUjc0yf1IJIz
zSHW0qBgdjds5oe07OP+rSFymCfXYZSnOQv/gS8EiKk93PeUZQvm/rLMZ6GdtJD/fRD5386FoVNU
UiGfTCYBhTIWX/unyl5Ybg+BRgyOqaWgzg2HJF8OmxFqua2c9FK+vgjvUPxmB5JY0xSc+MgYyUIi
jo0L+6PXC9nAL5q3mIzoMg4w9pVi+wdr4hReKHIjqbQ+F06nIqqF+ozc/FzPJx6lk20HL/zt/wAv
+K2zs4bNKWsrovOAhWsXXPTCE2F24rzjPLM0hXKNtbq8naTyscs9Zbhvm+rf3h5mgYDmKzM4mxEx
FkokPJ7xXyh4OGKCbpr+4z9miTQJzg3EU6hvHd4npviIeSU+clGwPMUNjBgPokZL2GzBEgea+9/J
UtolWlxLPB1QRQNwc1ZG+wmm6CsQnDLxYqjYlE/EGbJWvNR9XMKy2C7OKdy70GEXCgt2cD3UX2vD
rFi5B6gCpl17X14cRaOngqwSUziIYtZZuK46+gLPk5uDazoDyzqE4SaiUG9bBy8nur4NY7HtX3FY
VwDubZ8IKK6OBAEZGe4M3/fC4I9NLDjHh0kYlGnVSAeXkG0wL7CP1itgtuGVvNPCZIxq7eYAbqDk
upDg8sE0I/3DDcbd+64csHHwAziOfhNTRQPnGDzVN2Xz/hKMjsaRdqObfamth3vsgp7PkIbKltLv
zGuQiEUD2r2+rZhAmqR21uLUr/lVmgmYdGdVuj+O7/h6mpOtIA2QboJISRhpu/+t0f+fIbT6qj2K
wCp6SEHtDMsuc1G0gIVNiLkMDPikzVv1l8ftxfGspSbdWW4ojO9MDdV7GTZ5e3CFRKYEiHBjCnU5
Jwa1qUt8MROUUodzUL+lPfTufYEJBP3Vnsr+y9Tj1PBhd6Sq6BRgcaHHsmt8cOSiLgXkUCLr1Clk
pO4CXlqZArovD7sMGejoJpAVCPeukOO2dcSxNbjyTiEW3nOo5AKFzPUs+FSPGC8tcoCs0NytHa7U
N4BvvRLqPC1J7fLqI1/9YlFWo385onW0uMtyrljCj/+7+0g/DlVpTtksVUmXthlxJDAPVvn9Oaq/
DVA4/Xsnht1UZtvnLNR9Owhwenz2O5ar7BBfSZfyLOCuEpmR86FJCu9eApLjvkfNd6kHmbeit1ew
IAIOzrZ6HZmNx/RaLuPBpJcQRW10iXfd4DX/suudqLUaGYfTr4AQp5QGGYzgggC6orol9jBPwYcb
4N9FlSJ2NRJ8Qz1QjTRaTUetAUy97h2DzmcE2cob1Q2o2NXwfR8iNmjXQ56uSA1Drw26Coz0CTMy
fqj1v75pPk0CGp7+Jx25wnpnpuAqIVhP9jP3HAe/yllZDeRVlAj8FGw4SpVKnTB4KECCyWYWBEw3
Ao1ouL+BM8cApdn9/7qESyLC+AQ2ENL70aKdYlLWAbztzuiJzr5g8w7Uu4+P3K1RLgdMd+90M+OH
LNl8+DQB0wkPKf5nfeFebLtJlZ1O7tCR7R1UVF6KGgJJuBc+EVrhIYQTUIPuN1PApvKyapjo15vd
Ac0uOQ4oj3opxepB+HN2m+4Q0eMZ53C4U5UCSECZIKYfVw+Jj2/iEJZqK3t/tvLOD2uO4iYRptdX
966RIaP3T4zS1whgmxsqSYPOSYGSqLEJRhdCErExYnSyeFiX+n6BevzENL7WzmrtJkHgxeQjisNX
HqFwJ2UhXI0Mwy/k3Dv8/RqTu8onnfjjeS5ygPU3/t8rcnN1LyemBfhMQWuV7uy4aeUyLm57D3XH
59gB8XarQaFNCJ0ESq0fKPDxg4J/Z05JArKu2s4dHXi/KuIcRWSOy+LQoR32D8b9iTNkTBTX9GzH
94k930qCcnsw2iigbCM0NVeJw92E9JiGowaUy1xPB52cgoehj82DgwBPIKM2vFVYPVdqLrnb3TlT
z4I+Xd9hg5yB/Yr4tc7GN+oRWM9tDqt7mYTknoZPOYp8s+ZlkxUBv2w9nBLUhRBJ1k/igh+/SMvQ
ZJAEvI3A7/D/+cwQJaXcqQXzaRmnWyc6er85h2I45vqlA8Nr4nIDOu55uQQ/etFn8qOpNmCQ9T+E
hTv25kL8qU9Ai2n7LaN6YMU6+e7Kr+DcyaOz0R2qfdQDT17Rln6iuoit596dl4sqYj6rbqyObKa7
yrSGz4/MvGShCk9Q2aDFIr6F+DKERC82q+J/GIOz7BrIX24Exn55bSfpFeFYpjtVBcGmpWwvLSHB
+CsF4/SAGdKgzGSO/3ss+o4ji1BTfRi980t+uTaksmiI1Wf6AtRcdzBOR0wu/WJKkCmlXr8GNkT5
bYZlTNYitNIQzSojndget9D5s7PVkrQHQcOZsXSMvCOq8X09wpK79H2hoefxumV8t8EiHO1r5MOs
cOdPz1f13DEopek1dovC2ngpOW03Ew3MY8UUqqBzHyszwey/MbQwkvnuxCmFVTC/0314iNY8ytk7
CUtXhqticVo0Fm9Chgf2M5lNvjSXpia8honGBf/QTJo+cHDGoa02m5B7LhqOXrmBIhCgYvY1E+YY
Co7Rt6YQijNZfIUe9XH56Hdl/W1/pBjoDzML2Wp1OsuTTSuJhpGOsJQXcOgBhMjSbjCNg7YD1RXN
KNlV7jyk6SJv6j5Ov4fYNjUonkVb0tPn2JuVfhho2yXCpKinDogzdYCoiOOiyKIznmgPnwjHZpCK
f69/koyfAe8uI/sL5U5paqhMub+8iR48a0X5lJWq3DVfF2jNZ+qgugjoalR5aTE9lnGJLYOwqKuu
u8ElrJd6IL67V7R1YwzztOjLvdrTvD9b4hfGgfBTKpOWpd5BY+E1MNO317AjQ68Pw2fs3TekM6sk
Dj2w9ZabKIaghFdiFF4fYy5X2qQejNszc4cBszMpSVWmHk6Ix1pztKZKzeJWoVFq2SeycLNdu9Sw
lwIOG9pjlUa+20GpFVX2pfE8R1VPuBCmX0ZGxBg+BOfZt11j5znCbKnNe+oOlNW7fuEoHNa4uV6j
FLrv1Z1Uk5e6jKM2sCtj+9HZak18bInUXpFHmTGlPLRUV2ijweSsNfZN/4NetdvUYntsfQUJSWbQ
/Si305v1KRPhqfb0NKqZlwrhffq+chuXiB/T6Ctimq5yThXyQQpcoAJarM8VJWwgTaPCu2ZBjXQo
FYneiusGUzT4lBkvbthLielbq/4QIcuNAQ7ktUgraKwkhTOmw/lEkifilYUv3JsIe2adb19rLyqw
wgYf41Tb9iB+hmwUHWR59dtIL2LcrVn7sYudELwC9qD/KbA7hzxIrLwqs6eVFcWcklX+LNogrUqr
XSOqv+hfP/KXsXDYX6zeCcm+9oA528vXlyrw/23/P5RN6P0ZXSBBc+czMReiJ+LKbdXlbqUs8aGe
3n8EYW5hxpYnWdVXkEJ9SvvXH+vLDeKB/QVL7mdZ1Y4qdY+y9neuWDljzqdCaIdXH/1NtCoFlSy0
fZ7ARRNE1DlXbPf3ynayxYhnEi2iTUSszODuWvXpDaB1V+5a1ARGOffbSyVrdnqNtrnk7EoKyrA5
2hmrnMthtgl8URW36iesv46A/n50uRk7E1vJRfIyJwASxd8ajeybXgYrYIJBADvFLTSBy7zYDviI
6uYCdjanbXcz1DrVocmbSnvDids1wEYrxKBQzCapUtMziYAcEIdPz+5ND9kyIR3B10QzuQQJCQmh
pgYb+698N+HjUnqy/je4yL0oK6NHhc+j1LLbBLpwQCyYkgPhoFI0OkHNSK66hAs0WNa/61aJGiuU
9aEQGi/xUM5DQJtXSpm5N0clqKW4h69dIeo3lD6m0O54Emv4ZXz7cYP7w6hVli940hfqJpXXnmds
pkdCZ2adPUrwlE28cVvKqfYIY6aE/UM1wCRbu3L7N2nooHxhiPnRKqDQZsiLDw2zUQP9Wc8dtCG5
gFMR7ep1+LDmm/WZbG4YBribuDWP2D4GX9Cnx35g3TZQpv/KuEgcjit3zln9zXEG5vOwur5gis2j
KTgGAubmjvEuiZaEuurSGw2/sss3mCqeZCv3T1r3P4U+o68rScrnYBzM4S1nFLEQ9siBcF2aIxNn
h3jtTqAGpq5aOX2HKLUse3y1x505C79atTlni71cv6h35khCfw3grxk0bHBayWs5mnOF8UtncI2w
fTWptH0E0XZwOYxEDd1KmQSh6MtVRjdOVs5rga0E5ypnqYlvOMfuVaryP1NwIKKd+G1TJQMvnjUh
RhAIbGubKqYBVeR7mT4PDVNGOvrAPEQuntuxMQMdNQMNAQTspHh2m04QNUEOGtPeCZ/Sk80TQGga
KP7N1/R7X515Kmm2WNDqKYRTgECbYpX+fUYA9iHvyS43fJNqW+U6LSXxRXErvXz4h0aCw+dCMeDD
OEuTw67K5Os3fFkhuZ1Pz+t6wtIialtY0bUMb/M7BAZJl/+JNoYnnT7dLLebVbEkZ1Oj4uz5+X6y
m8YnHzcqMuDuEd+vqPbdyDS7jJTo5pdx4R265RyqzVrVmAwoyvTjjR/x5C430jN6VDWub96dUKDE
ybblW+zpjXbDsUwyhlFPvqzlmst0dAYhKgKmx4aJB4kzP6Eci4i0f1QJQY7/u7FrEwuoUM+QxnmX
rpmaaFDM6riPcWBuF4OIwqCrm5UYpnY9sAFFLe+kGx4dGRVkR0H/QeU0RGH/aJmsZMAMmHHtfaGO
yuuQMQonUg3ofT8HQF5QgX6O8nciyl5bmzaXUnbfALUnXbvtm1VfYYOVLLxkywk04amV365fFhIn
eICgqjVfejEJD8yPW7h3s5ykdT2WVLiLBSv9VPuKyVlhiT2vaUWZX8S5jA1phQ/CINba/ZZlUVod
shp17wb+Ir41nmW2edAHoOQY+58I7WLCzBOSRlmVqJAOLsTHJJkVAGkuPi4lOgMocTb/WSWmu6nw
2c6QIjKSDwe/uFzODgzEKL01nZeDlEP+2u6cuSdliPrekDCT+yQVatwJfjFlvXhZZ7Zs7KmXX2FJ
8xeUNa1JVDTn69Ow92SPs8jNO/za1QWGpefmi3/HOw/j5JcTzsHlOItquz/z+jcHKnKW8SWMmBXK
xFAlNbU3R0YrFdh9pqn/5SGEHABej+KCFLKXkatZSUM96vOIby+0U2qUzdnkeSkCjkNtHiTBbY+9
7LUtRA/I9o3LgGcERF72pudzNFrClcKlHd8JQi7+ySXcM69DOOOXGpVTlGJkLGYLKSbcZFAFPyuw
WPgoFuuDU+qe1loiwGPqxzeV/IzBW+s4fm5dvlXwSpDuQjWrcK55wmEiYsKSx6SoQ6zBPvQ1GGj2
BuWdGBZl2eiddi2Eo4Qeko7Mco8NmkR2GV1D4WP6a3CMNIFfAYGgTfVinq2R4y13lj75NV5saWmI
GizPk+5TA/OM9vUldC9ssQORbJ3IfpNVW9vHtYBnqDC9TDLKUJqE69CRaJRYnGSCpG5MxIjt6WjM
vaFz1M1qYjB2ktoqZB50R2sOSI1EVtlgR7lxgtImKVBtLU8gC12fb2WD+Oiidl9Iks01hLQ+KSpt
oP9FQBNlDMIWNHqMVIdaRUG+bEZSJigH2hhBBIDLkmxPFgmFvq/hFMPN5NH1dcA5htRVox6wJyhA
HndNLwcaOL4VsrWSulM86qx3DLOCTifrIMzXJT4UpdFtjoRJA9k/pSw4qhz6D6dWMMIEBkKllibf
jEq8WH7ZRUJM5ftNmH0AAYQhMDeKmVxB1iUoM3JA4FlTbskNpucsTmZaEmVWJwuJEnHcoT7LsVSe
oJmojEIHj3mdOAwah/ir+/zEcMOgmsBzykTilLmiKgxL0vlzSSI2n84+OAoDAKmGgEdCKKLcJta1
PkppFZyndzIChGCA3OgYLl4odPVzCwkx8yQ7bNLaLRWUROnIQuhO7foSTLGMLA5PQuFl2C6cR6LS
9YtGO09iduW55bou0LaCbZa305mtDZlrA3mf4IdOkyPnXF4Y9LNEGNmWZ1C6p78grGIWjSk9gATf
zP0JRFbP2XP4jaqhdt6e1mCcQeGUHPCX+EsRQwU7KqAErFIl5S3lLNCpskfanNJFxcjGctN9OECi
P7OrWWd9tPfKel+dN1ghpCjNZemuWsiaUtsHja1KDP5SUrOOB2aOHoID+Q1BjYF8rUQW5I5+z5pk
dRx4O4CzrDVzg8huGKoraTT7nukh8tzpo8C9At+zVA0QXoZSFdMHg6+Y4TWqtVVB5wsiIjjDhHKx
0oCtnOoN7MuA83EOVT/jyrtq73ce+WKcKj5M6M2GMy7XEQknzBBwAkRUsAZdMHcAEQfjEv93rlLI
eqrwseL7CdPg6QwST1SbWyQqlTgtfzQGb0gn3i9Cs9elGdTV6NH5I4oZBuNdjpUxtlb9SeaU4tPp
jW1Bjd3E28/vTJxgRZHGPM/IUuU7JAPdyFSYhvu0KxjtNcvN/A7rtPCqheVggNfLu3jJVj64F+8i
d4+ziz7KSZUAqjJL7e0XpAH9iub79f/dhT77FJ9i/i5ufazZie+PkTOvA+yL3PrjIobQkLp91J/A
clE49y0ZmrIpDzKs6ODNRbSXCzs+foOvbNKie2bi4XfKOuqXJbxpSuiyG1HZ8utcFogmLatR5pfD
Qg062HnjFkSXayIRzeNUFNkhMZdqrYY6GQjAoVndU3XtnnRa8D5JAh92l9UeNz8t7/MfNNg9g1vw
MWTaw9Oxq/aRV3lqAy78G+nDadx9sAZQoDPEIoO2k5nH1ArI6QqPQL8XtL1kl1ZJNPd4p09X9F0C
UP/3ik4RYT1EvwWz6WkAqTx07FEGYGHQDcR0N4Eg0gkAJDbspPqThJNshVa3alMHHEr7lDrzlW1i
r9259IWDxhet13sSNon6H/B6k1GijvCphWvmkQ+BEQ5hV6Nu52bNVFwLDBw8qs7Lt5p7YI3/snu2
ngsAswOD+uxLqB82j5zwp8jSElLv6GKmWB2pZZ60PlazUVEf6pTO+yba3vmBpR2I1Tp9BVevCmG3
F7/Q8kvk1eJ2IvQBapGO8j1ME898bmpcIdWkBtYOJZwzZgmkxwY5L62uQDVFqBjRU3gpwI3XSgrG
ndtMidIuTssuSxpPF/qLeD2Vs1sFjuPs0y93dRfEvOjZr6MwpZIbrixFO8XUkSUiIVVaEva0cann
zu60R2ZlUH0dup3Yqq4K7OKx8AD+NkN60i9HwavJCh/dsLN8QN3q786JZGPTTazb1SJSjg4VuR39
hZwZfqUxulYmcGlnzYYJ/G9vGwQP1tI8+fWyYRZ4BqIGB4GuZBY0eixOxOceGRMzP1/1/WgZEhdE
+qNHoMb77DmFcSnjMLkBk/4luEddxmRSp1y2DQX83cPO/3Ewq+63w088iLzTy32l5H0J2vWf3qcq
QoEyx/bRU/+710uOLDi6UZaHCM5dDxS+PPUbHGECEd0iw+FBP6BUQIngUor2rhcIzrLPHbO3LM/d
06oBP0fZU0fV1PzombBRgc7BhSKOaVgh+462M8iIDQdV+ggHAz7KrANfBiaTCDD3EqENqZRIWl3K
tGYaDIGdKjQz37j26a9tkpux+OjQ6790/JrGdi82TOQejhMJxarbCQHpkkHAc4bacySRFMnhOHew
3BwPv/MB2YrJIYtIaJLBbVn0a2rdVZ96fVgsqrwWov0H7luLkostg1GrUGozv+PJEdJv1/mUwq0r
xChOhdNAgy2kHvDR1cZ4/jGUd/AKyV9xfDZJmVJyiQ0s51U9PeE/qJl2abaHKyUSf61iyNLf80Fp
Fp1smq0b8Ip/nt8DrIXPbAfo1N5D5OU/lGn6vRMMbdJmooDPmlK6gCBvJdlHT6oVuBd/S4oAXmH5
vRuADHpg1Zb4tCr4Je8QXdCeTn1iB5r3STawR4Qz5G0uWF+7ELekOH+FzJRqfcpQFsPZT2h1nHnN
r9zdp7gpZQAauEVaDWFrNRzA08Zo/BmzCtF7YcNaVz1PMuy0238v2pLTLLKJGa5zRneHsoSHFAe3
sVGyQ4RtR60QTK7ohq1MryL/upkosRJ5Avlv100bOR9yH3jVDFlbdkGZEN9h8scPsxLkp/zg+fC1
IlMjNUAyuQ/GCRufhHEQQAdSwf2Gh7q1gCAOrDtmqSO1RaH6rPAHTJSYZJB2HCk/cdQCGRQAggP0
f8XIlXQGvSiGCvm53OTJLm5SedOBsYWOb6xEWB7QqEg5xTbzAXngavNigbrnJQXF0ib7JdNCzYNT
xn4GLppd0aJAXUWMV5XuIN+IvWYAenJflOxqG57FEsZ+P7phffmfxSb1uEIgzG2IlfmhmuF/2lmL
Kp54sHIl0zzr1XEu14gHXXVGooP9wEH5D0ESI0/QnvYrf9qVWjRRDsOS5oWvc8rPK4dF70ifgped
8X6J6+KMV1xFcnQuS4PYUxC9GikAqdx+1tHout4Mu3YNeeMrP66D9cOVJpAljb133aH7RrlZViBe
odcmdZ6gD6DRC3une3omdoOCGLDO06G3feAmLewTbUMl65BmC+/8svdXSZucBALp625eDIPoN0Qn
v0Tn8T7rLjqoImmLJqA8KM6l9HLN9yBYALR66RMTtFSMRxJwOfqm/+ZD+GRAdbPa/43LuaG/c/+w
+XBl1jsUj8lpPQXZ19L/BqfOrwZke54H248c7bc7fKsbLSsNMTUItVtgZHtd4ddhQ5ZF6MNetwQu
HZyJ2DYZQzzn/vU+6whSmNVQPsWk3ei2zuqMhdm++riocvc9Of/D/nRsFPBJ+qqAmmyZPwKn+c7g
iNK1LwxKLVihFGPOHMY+tpyDMvf6j9HySwnNQ51La/wIxzVN1CdkjkwC/DxvaSO5yCEmxt3Bu/vI
tVq+I0weFA4bJk1B1I5Uxn4MFOm/HWAU2r+YsvyUV6fUhk8T9k211c3/TKbuO44zz+95xkPIQmO6
jeFRxwn3+GvBFr5jV6Q/R2TaxWcA/f5R8Yqicz/K7qOL3bonTnbLL2bEMVvMP9QnjNlIo1Qk9WoR
WRsFJlHX1PTnq55pR/gZfyCLaXYcfcO2X1oMWf56Yl+zKqfjE+rijbvXa/mRBN81zY+HClTGTCLt
fLZ1X+125QXOZSWhDJdwWMpPzEzUE/SaPUZYrsSoPJVTIetsxfM37p446tSJcLzs2V5XKsnbj+JH
F85jziVCzNejEDOeJ/b8tfNm/HR7mu0QbRMDaTHphmfymUS+pLVKEXdPGaYoUUHLZODoFZdLFkN7
tqz3Aj06wBBcTgFhsioLOLFQsV6FASyHQblHf2NTPr+kkTRhpHTAecFaopRXsPn6mzceGLlzkYYd
mBcsX7P0acjqvatF8fVsNRH+zWutsB8eb++hDottrejGkzpmsyn//Xo4i52kSygHsvNdmPwJ8Vls
eBIETnMtxuY+6ZEdBdyX9WMOeVsS8xHDwxZ9+IksQVDv0OS/dJKAZE25mDbP2C1iaU4jDkeZjZcv
zDeREMyW+D2goE7TlvFTwCd6g8th1hqyjwHIZykDDSwfsrFqKSDUX5FGPkkAhPf6wpwiN8uJoQvM
YC8nGxccEBIu/TWTdpDykh3FUogbVEyQuQjiNYJj6MWom7VihvKvLx+d485fI+iC3M32WeMr1JMK
Jd3HOOC7aS8We+Z4odNf3gMAc5o/UHdX3aIkoFXzJ8v2ILcm0FOBmLF0VVrVKck6t9bxF6IQDoAy
g4nqTRUtsiA9vMMMJWBxCQ4MS4sHUS2SXgNeQUGzsh1C4rWY93Cn2rXG82wUUJUJYkike1SbmmvA
UNvL7v62NFZ4yA+8zMSuNb8hZfYwuCcc+o8ojphUKiCakI3zHY0Satkit1NddyMwWhboRzyBH5u+
yaOfJeudx697EbrQN0bYww84bp/dTQug5jFibbALGHSxnhatR7B1oAVXxYEdULLfKt/1oQ1EIIOL
ZTj3XYL7I3pYKbCo/Cgw8kYJv1d4gKA3i6fmQu79mE4ZIcUTSWpp4qKqEwzG8FqAnOImorqRfhE7
X4TJMOUINh0YaFP/P9H5yPyXX1+9lRv+QzX1BNVo1BVt88Xrh9DMLCij33dZiT0o/TrH5wbj4snq
DLyLCz8MmChiYA6e/dYv+mA+Dpte1nGvlqWTrhQ1ZZaT3LtjoK6J9Ek0RXxhLSJJubot2uAbFeWl
+uoGrsfytF2zH0l0D8B5sw3FC4OXEQfxDFpsg3K2pBB+ijbfwgxoG2LDi3YGKjUhEyA/M1vEBWaG
yH+23Wm0/LoAVvl7Nq/rvnhl4tggWzKnD1AuzRnqe7Z+uuCTW6ZmiS9Q++sUqw/k78S+9awH27k3
yaZTDNtCNPBKeN0SPPIgFzGYo+4HxIE2+DMNb4FUw0ku6ScARCVUYidL5LYKvp1mdrLdZus+kNIy
gfjrq70swVZ+leONzEVxbqZzbZ/qfVMuPKlRq5dv+b2hvx0cMBk1wc6QvziTS/D024YaVkIwhNnp
oly6bahRWiLa4NwLmS4sCy9GHGI6KzVgBEMRvpnBKboqUTHOBSdwEFbDuPhz+L8tao6KmihDKHGu
t2y1VoA3E6t7hALOxWZNz9L4bWhi+qJx0j7OShT2fiRooHemS6R8afIh9QB9OPOGkcz3kfD/A4Qb
vCqzSuoc0wtX6evyR3yU5djf5DLFZB19HGtgHizrn/HVI9skCZ/wKCp5psRuQj3z4NjMT1GqXjFq
lGqfiQN3SzqifwXBoTqQWFYBBys3P1lYwuyttkKRE1Z/EbyKpd3d3QjPMng/n0xzmM9Xn3TZeoCR
fZHAtvtStNgzf7MCvPysU09nPk002dG+n2NfOFaKoPkuWQxHi4o23VolcIrTvjiKwthK6r9qgivJ
kOQcU20KlLTuBeOja0sHUk/BNbWW/np0q8xXp7CR5hnwuDgCoGpA3rspW4eJ5cSYKrMmP30946+c
BbrribcZakokAxxdd5Isz96vN4PnoNlIISZTKXI5BXbj3eF7bksz0bnyOQ1tYthEAqhrsX00V7MO
nWVWM6ZWiIBnYxIBbpwR1TKzRmgAX3GnMH7fgHawacnEwsDqBhs9mXQlxpedv0p4yShKwYVTegsb
3PKDcjXH+H794w80nbRo+GYw57o2qhyS72L0ISLfV8DkOZbV7Jt9DG5qc06paPGde4Rwx6ilrzbM
a8/0pkeGR7E43bhoSv3HEVohPocH6vUvL4Ja+LYJgqq/p8NgsDGLW6T3o0Gwb+s5NVWt74fakLMw
bz+YyMVPqWqOI+c1bg1yiAEhcQd7Uxxy2m2K8lUgyD0NAb7bmmMenl1Hqf0dNcMs85fw2B3rn66Y
3kyBziiNYuDHjSHnb3zeJzatyn5IsF+CNwOzJaSw4sIRUdUxrMo+w3vzZGevKEUEm2g8SUqlz8I6
GGpjx343YxcM9gCslJyih41g5m1UG3uVUH6S10Qkh+N1GvpLpmEtL9hBJJEY4BnD6ms0VnUOSwQL
ZewPAT6kyvZ4WZ8FLmt0bSBWpOzepiYP+qcK8FQ01V3JMiXsjU/OFRfbDciP31NF+WaOobOMgkF/
jlw+yqY5KHIjB3hBzFMvvz/tXaCu28e5flvE2bTI5IwbPQ/9gksH6i6lCImVFhHmDIOct7mtmvh7
P0hZ2wsUoudO1xpmi4jRMjt3aIgjBwHxCTjYo9MyFptsXx8TV8DwECVGUMtjyweW6z8XR+AI99tK
i2m4VY95w6aL/9hSVhm2ZYxLgLf5LGMF3M5BeCqzOd5ecZiS2hE8akm5PiELUlfh6IimYy4ZPVBW
3+9rz9XyxYI5LJQvoahfelRMfl3D8wQlqLzV1IjVevSssoY2uoGM8dStY0FKFt9TKQavtQ+E9YPa
1mFSfP8hnl3rtiCPQEsKsAc9z51h5egYhtnUiij3soInxCCOmGmmEv7JQ7Mf9mUPGJbqPXO1N/Sf
xvgbqACLbL4qXRaf1EDFH9UqX4xiLP0YTwFFm1gtN9R1voc7/7Ba6lGiFEF/XA7keoPVWtP8KJFS
M2GKbn0DT7fWFxGYMlaXqNxUzjJtVCjjDm5e8/H4txQiT+3wEZ6GEDGD8etXzF5aN/RH2sOBp604
zCdJieX/ol28crQNGryrRCrP7reYAPSFqF6LJ704qhohJ4oELQO9XgJKuLmgGZYCowVFj4OU1Pac
XA+mEmsdMJNqfGNNVsz3lZECjHy243cMpHUsNgOqwOLxC3I3XCuTBebWSAt9cVfu3ciO7zRAe5mu
e5+bT0FQn1IjpvNP4M15yFIUgiR8JP9XYwsZVPwbl4abH1BeqjIhgzWCztkSkeWoe4ynJo+hQqxs
0HScHCXagiWPWg3ZguhQOkNPHjtkV7DbImPYGdlDuovv3kZ++8L5UERkOsUm0OutR/+NkUjLQpCb
24LektacAUwnnrvH9O4RpkNsJfdhlnseWA8H9Noy8+yevYJxgFcqmT88uEs4SM8Cw+WKYnFMxpiJ
9E1a0oYRM83GrdnLmW0MAjDclIk4LDLJ1Z2DBv5/ABjhePQ/ESae0prJ6c3m6eYHxfcLyuGuQ9jM
tM4OyVdN75YFqhybVj8/p3obaL251OyHgLfOjKJb2fCCrURQXq4JZq4YkZWu3acw73ba21EhzbQJ
96R8Ne5XWuZPeuh8kAMptmHLRfkYXb7UUaSfSpu8954Y28V8kghJy+/hZe2NAg2Op74nbeSCUK8U
0zv6sdFlkofxUfh5PX1PzZ01PCvQsT9QZz3RPioOy66u9UmfAh4pIi7kI5gbFDX4F/nURdIeInTY
g4buyOmHGkOfvOfd7exUSvcSN8eDLz2yXPhOG64TQKRWgQVvRwR/0eQN2KAsZseMIGGRiSMEDErY
YL0LWEC3rfX+xGXv1nmt0Gk/rtJBM0SmNSMvVqOe5mnZIsYh08BFSgfRbJgi8aKAZxvZGmnnHnaC
bHvQb4iJycgVVpKfn/chuLL4whyHhOH0Enn23sihF3Pz2HVBbpgKcvCfw7JUncQalrmy95JeugbL
OG461NHmAlpAqrphOV5lGsy4VAGhQoNthCS1RZzqLMx/Eo4eAZZKa6nCADfkiCsuKiATtsR9g95T
s2Hlk25/7Lh3m3meeo04EGkytFL+GrN0vhN1eVixIwz404MD8BjRvXS1X4MchF7qcgG57aBpxjdh
DtQALCRlGETDat9s4tSSx6A0zO6kxe0OQIOj1QqGqFrzN1rITH4ehNHwSTveaQP20Od+Z6Z0fS9P
+0C1+RmQfuYwMYLBZx+k1x6oc3+EafEm/5e7LBxKvZs8ksZdVOfpws62g3D/1v+jQgv3WRIWBBuF
/YWauRZeeczudDrAiXqPcw255PMgfqDxVM0QqdtD/x+sQQeYf6MCsVuAmDLYQ6Di/jitjdGif9sR
44gwO07dzNNQfdHbNCthraDh2fuI65O2kAYNLhRJnJ035yNQZvC591uyf9T1CsL4pqkbIboGU5T/
cz+xdoqLnQC4fB2nEwF94GzAw+fexwDGlpy0rlsoh56+GOVpVQ1Sm/buwmi4tZ+MDL+huD96kZE7
nERFdR+6LlotQx6vG/GQelQZSzucHjHi51MD0b6o7vqvOzGRKpTrCoBH5GgH8IqYQfaIDoF6Hh4y
EAvrINkCjKjo8g+4SH4mZhiBZcRSX0oT63e1FK9EFOkeJKxum6LY9yhmOD9zQMkFuX8PC/42NYjb
G/CiBSvBYMPVZ4KeuwbfV39RZUf9GifnrY8kL9fFYu+XZv3TYB2KIXn7twf3j306NkSw2Vw/8pbG
54xcZ57chN/sPudCXlKyKheuP2s2o0NXf9qY51y2r0FVPOFE9nXQ1pS2mFczUUoHjPDmALqWgQoT
x2EEjubbLyh0Lal+H6D4/nnkN32ftBMAg9Iq4izj6uWYxm67f6lz8a1jZ0paa+z3Aws202TWKhZ7
Rqs0nB6m7MkDJ/43QJcwmArhGUc5N2LoxHc8U5AxdUm5j7NzLfCH76jRV32x8QvCCLi+Q78LW568
Wd+wwyJIzWNOYFvHwiTzK8BwlN/VajtVb1dXIrVLw/ABKNWZQoQwzDjcvOQhin/tuUwGS7i9tWXr
Wnu0tc+IR/cxUQXI5L36J16Cyb2Xkdbf9EnkSew7mCFtjybQZU5wvon/GoUkLl4EJ2ATXCRRsYJL
XNPQXEIUCrMzv8u0hOnQIGz2pBfAamKv4FPkNyqFrvMbPm0UgO/XBmAPOFsHARVz7GZzdh5qfE2N
FRk4mVYx5ZSQeuM9AdpeTDiNkGVzrweuHhAC1zowQhb4z8BUOb/EkBKhYWtuwV3rdx2JVbWlaB6a
e1rSpl/lcksoXCmaTdJzFq0BCRJIpj0aNEGoRIQsPKNUidpAqCNyRzyH1XIjsaiOhpploDcuaIiA
cXmOEoXACi9eb8ELGAAo0DDzt4vsuTSWkChcT5FUuLSI3Zv2bFq5opAFYaeTRGELPl0BSk8XqOaB
3PAmgJm5Y5GTScTDdwld5rvzjFNysNLJpYwgXYzdazzz3v8WJc7VxyaHHN9yz+E5V1RHQzJWEZlm
VNdW6vUJEW65sC2yG78OTC9AxbVQIajM9LAPZ53meGSNzaFLpsDEe468iVt8pA2mBBva0auLk1MG
O4Y/8AF1WHpgqJaXOsmJ09CqP8PXX//0Lr+iKn+K0+sQtKiLIKuCq0eKsmqz5t0s+a7mrVjDUiRw
xFcLpN9EGcyuSeOLrnwfXlR0gNOD2ubmPa1uGAeZfWxLKnE8/3X/aEJBEAuZAfvcYBaPnB2JPZw4
lWMDJAoBfL8OHLaQ/bAX6witB3QxDUuj9PP1dG+wAmEwkCT+NajJF4amtglI6oHW5tokfU5E/luf
zYNuX9Ten5ZZT0yuFk6PldOp7K98yJZNpkRaSM+zOZtFSYnT1tHCq/Zrs8iynoUIvbhOeIg+lvAP
4L4WM0mYLkr7/cxnYf6g5mEiQuDvJuuctSPmMSv0vpKMkyU2q3SrVjC/fWk2NN7DXxPuzlVl2VHI
VB7lkDwiDEYSzwRf3IYJsNRVKSgSfEhvj68NeKZCM0+pWp3SExL3ZZ4uBa0az5k/VtSR+Le38LQD
ucFBSMb5z/G2A2DrQ4wEQimrWmy+BqE9A5f9M2NYLbcdQjOvqIUGXJP1zPfgjtUNHVlrfvC1JM8Z
MKxpSuVjuyigv4RdK2J7mzuKWqUHTK5STE9Ea0PCkg7v82tK17A5w1eJoi2A29nT2UvtD/A5eXlO
ze0KAsDWLfZj/VMmYJRidEK442EVZ9bW9MCMQpHS/IM5ANrMx5xFAs4PLdLPsOKNP7LPREtZCef1
fdxvrbUyYlPcKhuQ/6kKzeHPC7YJ/p8w1VdAh90s7J1q+nwm+EhGk+A39B1sQaaCt8GuSh9JSqDT
Q689MUfVb1dT4Iq6qqPYyKVkoKtOJF5JJV6Xl8JdYGrti1sd1dI4cYGGskKwH15RmT7HW3/PO3PI
ANzsXAHu9BeILalNCCRTkrwIJ6WwxfyzCqKX3rpHS5pJX4NeiRiPCMEudm8E37nFYoxGM24LP5AG
5R0ziUYlaDrOd+nABzM1sTkxftL9cT907fLGBsuIRnFrJGxy+naYy0tZGfzG/2Kt/iXKUTP/Bcog
h1uB0lLx+NCVrkiN+xuqrD+QeCec5Pnr6zcg+la+XpBC77Yyt6BJVrn55+gnlZsYJnjh9PpbaqiI
VBKjjblolAS8mVTKgT31tLu5Bm8hyYN2tdMS2lhjwHweni2QUemI+eUWX+dMioxJ0E3WYIa7/jeD
pCNsISTF6U9RLPnErRGgB3shnGCcJZHs3jg9X1/v7zFjEF/ZFdS8BFlEWSkNl1OyLpH50eC2gPQZ
vbu3PUJG4J+nMX6+HVNVhb1XZFWLwfh1faqu4WuRLXzHVWtJtbYxx42qtKCEp+QvJdLBnhMJ8md8
9qCM4JPtSJIxORybUzqiDwVkKHQM/Am8EFIuAmMkSShnVg3Wo8/uuHQ2RDqH+oAc5gcygsGNarDA
yAZS1nXRzBf/JGnn8TWi1DZgBu1VTKSRAkbPgb+sm7agerqJTdp8S7OPdg+U+4Uu/YLlKr0MAzVX
Y76kV3YcjrtqtVUyrMxi7Z7nqeka2EYabeVHsdrMNhU+qGln0PXTbjZtb0pjnOXXjC+qMMk7Fa2p
oBi8rYhgrHItNzIyYOLuwkOWyxEhmFxxgVqmvosaAy/hpH0swI1vl1A8znD40dPGlAGWS1TsBhH3
PzUG4B8ppLbJU6HoCZ+yhZssj5eETpy0PnPstCqc/YraIBewC4gJ+o6jjLVYxUrEOV+n7ihnBReJ
AgI45ZFpa2ml+0SYGRK+HeFxlCxTt2lKRaBJX01xWpbfYMp1HRlUItjwfAhpcfdWqvUkzPtLJTC9
iTVn7szJPZ/dCyPT8xnfe3S9mhMt9a0N1io7qouKa7YDZ8pMs88D2M6n7vIUlOGk4XXd4IhrkUNk
3hoi8uUBKxDRZAUJkSKAO9Qac2GqSFXQomfP2r5/kBmNaQ0bi7Q/O/eoG/Y7tUZsQrzgkOdJXnl6
ql9Em3XqlGz6BQfsLzEoAr8Ta0pxLvCipCPtBVAgeae7ZsPusvWZdE2F/QyJap7tt58ai/H7wANX
ih8/9TbEp/1ZBkwHc45DJY9mV/Bjv3UWIi/klKK7qCc06948NiR6avK+RFyQfFD88kR9JTYaRzUj
HTCkITP2PSX0iwOHJ2QbMxAHv5oULOcaqbFjr8+Mp5PHFhU8CHRn0SKVuJOZ9iHlGGiNpiwgQzvR
6XxaKVnIbZhKSUefeDLw+/qkUd+J74P2H5mYqK0AncVbT+J7w+jv9Y+8J7qZENMB7Caw56F2MXo+
SoBHN4Iy4ccyvR3jfxOcMb9AmC8C4y4HURisDuvTsDx1y5HLc5hUYmAJ5MiNX937k09iGSeEHcnJ
mNYfxb+QDnUuJLe2KcCWX02eIsBzsjXOyLLZ+2Zqx48IZRO9dxNpgNQ6qNc4q4th9OEKptpdPq2c
iYaG0393pJjD054yM6NMRGCawtvCQTiqJr6EQ91KEvvEcjEOVmHscuEpR8r3HLB4SFCeUV+UHCsY
cdX3fwpXPfVuSX5WIpN+7CMa3uDWAx2Gie5NTam0Jbi75h2oHFFsnSGp7h5PBERaZZuFNGHZtNJY
Y0pbmQfYJ8S74LKWH5uJ0nMyWzx2QqOxugRShiTLK5VZFXKpi+wRHi+0tvtxQqIaJTZAsK3wIigG
1DExraIYqGsbXO/kOGvEjhfzVuG9IggsTTVZHWxaodtCMD+j5cwZUN8lAd5UfVJ+CQKbn66FMUml
cGaDEj/18fQimCNBIO58EmBMfVNznpCVlJhHASGufLcgjzcxriSAy6rr983L1CZHNb/939xRo6Jf
AF0jRcg+PqV7gYok1xGuzsl3+eNnDcxB4aHiZPlLegY2mru9JapGhGQFEJHnEg4Tr07Ns0Sn7nKq
R/smNme34CFKVa/nQqPBYWM1mr6fHN0xeo78VYNV9Q5QIthvK12oZeCLPJ/DiCxbwlNCW3uLq9Wm
4SAoNIFLc8CHvZCPiN9sT1vuweJcAB9b5Mm7zH5tqeHDG4UIbaoGIr1rHnh43Klr96qvT56P00py
8CJ3BAEJDhwVkMwKCqLDHBIGfSCI1N10NgFwcFGIn96tLFdoi+TbSjjOhZLBWRmSTWd66KtQQkkS
HTsElfah1l5gP9ipjGMLfEOvypXdSPOPxVAda68T2JckyL3RPxyjCMbBxi2NxmRvoBdqAnpY+9uI
d7ZdDdQNRmwAHl9OGxdtEiMdp945HKgvhJnXklQYuBOqapyFvoJcd65e/wJw0z04IyAs2XgfF8Sm
VJTpjP1cGYxNvtSc4k3idVCYQ9IlkCXc33gB1IqPBva1cs3Pz32d5V/GkdR5MxIq5Tipw9M1eqMd
p7pO0YXTuzGCKPKKqTfU7TzwAim8bt07tWgBsnuq51kPfaJTQqHNhi+rpO8LApZ37FGC6P3+FaYD
BHi8Eelfmxr/1HoXbsa2xJGjIXKVdOa890bFtc6HzU0judI+H1Vv0UEBUYzwfCk4Ig9eXOSUOBDl
PG4euLmVX6zOc+VnKkxtFa4gvojsczU3r5sZvINuRme2xAFEUvRk/6/KsRzE009QT2Ijk2T31m8H
rbCVK4/b+P8n6BZk/CziEv6gM2cfZEIPQ9Rg+Bi5GV+8pVZxaMog1pIpZSX43/6RNZ8Umt1J3mQD
c/EF63k25RumI/vjqcXcmunoJCOgoB8FhYYRe2hDF1divlsFzsiwcQ/5bSm5STJHrnKfbLDexWGL
3eAMbhfRrRzh6VvL/tsN471BsvUyHQVBIL8WFb1pYRPXerMTtssA5zAoJnzPNZuF3bL1eUGYbrBq
+0klK9vvcQX9l4lX/zVuTwMmHIhwEWQkADzyl8gxS8Ed9THLW6Gc+Hw18xxXoAEjHBKh8Nc0T7Ac
JFODfIlW4vSoPfDvDm9IKnk1Z4bY0QxAlX9o3ES8A69gS9gmTiFnzEx3BYgJxMSRRIgDHiiuAwhP
ENfRaGMBXI6iCrNi9xUT5eohKidxgt69vp7LDCqcQa7V5TapN+wx8Bs4uCFbysEGNMO0cjUIyPRm
GAcdQYAGt7pVq0hEeggaBlhTVXeN6dps0b6ZbmbmjwfmF0AAEYPUw+6ND9KyygClVfEgQ3HCxork
UXQBdNV+IHEUQ5USEUnYKh/Yd4xu0Mz7CM52vCFWqU6fW8lShx0ZotIdUAPA/Zf0L92KyJD1v5kN
6vqlcj6losjJiLQcs4g2ioxuG3+e1caf7ZvNP3/6id7t43lpbC33MKFiLNE/q90DJxI1XxImoQty
8TAHwXbDcZj5piwlfpXoYyHkSQ8zyRjJF/D67Xr0L3Srr0zDF1BAWTbuxg9SOYgbhYPOkuPvdIPq
4RA2wXDVlsI3mLPMVBxt17tLuiHjCk3K8USZ31Sjb7UcSB1WGbDSIBdTU1BBnSwAt9TBp+WVk+tB
MYUeLFwlByswMOs0a7bI+VykaZnOgaHdJ8qSRaZy/xQ9PgadHVJBVZR+Cyb+kbhO4Wb4tdsBtAW7
wY1vNfVJHg+6LKL1e5G2tfUZrGvji7JOtSh7njv7ZuwMo8gjkGOTndbBOzp2cbhB84JQWPYoy/5l
P+zwTSKEEjHCSC0vfGdsMj6B5xk0mbdrMW2Q5W0unhEG791W2HbXJvy0Bav1k4M1ANRVCZ91Bjqu
yLuXiiKm/gCutTuoHLfA7TLp8wuFkwxc4lbphRuGNj+Forj5lwDhEYUiuy+7JqGGNIL7Kt9qpZI9
+Mb0Ynx4fpHRxg86lEwWmiThjdTMMYkAjae171eo9yGiKbJcQlIynBbQOn3eO+wMI5ox0pN4we3T
ZgkSK4a4cz054jYKxA9+pVEdrDYRSRtC86aFH9qpEEu4dAZ681MDXt8GUhn/U14ZUiQ4exEVv65B
7pr+nNkEp39UjHLiKCQ+yM/yibygLoatP1n5xZwAILsKBNOl/nsUfnQDIA1nWQI158p2QzzOfZQp
TzKwjlI3Jyeyt/Fxj33eJQnzoFSP1aV6B3BpZQyk4ulkMhd8r0SYxN7wFMCAb9f5aPOAvtIN7ms6
Q8TqRe6mJL9gmYJ5ix8bsSrerRJwC6oSkA4YLJQjBFEWECSvcCFDfhViXMCGR+GYnDHu8JhbonhC
kFsqf1chIYVeiEXY6DFoxaUrchr18mIShMtFI3rCetNonfciAyJSY3p97JqK5jSrgXC1LuKMlGPM
GjkL0DARfc/OIwZ9bhBQO8YfLAR2rZki9zo28yVd2jpR61/xxgD2pkzoPip4M1phXZ+jbS+/Ezvm
HYhnNW+im/9gE+5rllDa/psc+hX+SEm0l0F+jiSZ7pX7lp4s2hUQyxa3siuDjssTb9jk70HmPrhO
6kFio8hrcJFFOc4etpsxObMJPyXJYZ0fIjQJJZAypdnwv5izJYO/r+wiCnXg1Q8Oo4kHodIIQYmp
g3/SRCpK5zgbKpxQ9U4XKXUrt7YhE4FLIhLl/zrvnGvk5ZoqgTRutzgtPpG2nfv7tYvQ3imboTxm
ZXfKxQgguiojncMPHMAylDv2Xu8BYO+u94ZD4IXd25Bjriptm5I71ubtyD9v7v49ElwP7wT3CHFK
YucsN6jVziWgEYQqkx8hDWUx6GNtJPLjy1fhFbmLaeEXIb2Ev/Q/SGtWAVtgrs2HdRtcU4RY+3mJ
+O/Q+9M0b+OIomL29onWuBCRCvdWP0fWWt2PZY35wmXuavQLy1UFBk/CYn/sZUqRFmxN3oxQ7aaA
ZwiWCUewGuvp0/3XzeWyLnKPdHDu5AnfDrI4SD/ghA2wcK0ms5XoSAzoRTuAe2zT0ogTazz97/gv
QWkevJ3DeI9uImLMoeRqyTzbwdj5KQXub16XikpPfJNh8aGiwbw1M3pX3iBkvZAW32p6B7a5YQaK
OtmdarTY/6baDmIK1ZrSuLKk+4VR0aH4dynLgrdS1+vWUoL9Y1Ns8IoNBAsXerA5C8Re7vwcjCzt
J6w9v3zky1HltH1PmVkKXpsJo3LTrVZ6iapz/hEXqNs3bg2uCt87whwukavS1AmkGGKNYdnujaha
CJHjK60e49oHN/TmhzmQ3fD4cUtjUYjOrun727xurN9M8M/HXFD1YemMpmEVYOieX8ieWLoZRVDq
ewfQdn4MlPW+ZGr853kHbaRKQAshOUX3Gvx8P3iD++xLEjMyC/Pfd12PKLEQ+8XD1DgoZ12rNNeL
dgl1iohsGjWp6g650dsg+/4W1fvQ1LKL4Jb1pLDa8EwW5txATRnsnIS36MxNq3OzHrKkBqWOVjLh
yws527tkKwoo+dkr28ypxUu20kUp8i2VwMJDbhrCH/tkTo1WonieprXmHnG44ICDSTMsLx2hb+uY
ur8Ue+pHS500iK2lLqKFOPcI0gZFmea+DZbzhj4X8GICWBBI4mhj+t9Xffvuzu4QC8sHMKLmuYli
lWRknSLXKZDd5+95FTJdoqhtc6EhRmGJhViW7yhAaadwTjKMRmfJReUMDwojRQ8bbdBzrtKcedH3
RfbSz8NLT0HuHE7V5CD499WmcUj2WLKGKg/F4D+jNdS7aKQqJgfXgLh7lEYucK7bdlw0E2LBUjed
RnCCi1rB+vEEsq5o0UJ5IJ+GWeOYEwA2Oquc/zkXuFMgzO3Uua0N+HfjVLAYO8mO8MTLQp8iGBUi
B6kewCV0OzAgojSTI3OhwvOCOWuDbDfJhSl9Tql5zyGPMYggtNxt44XUtBVKpYNL0Jk8Ne62PVPX
Kksmr6VmGzKN4qg3sP44OfnGI6ULqR/KuM8ZrMkoFa8EZaPEetqch9KH3ki5ekiSb2VQD+8Lin3L
vBBd+XzAYPIRYeNZ4/0KJiGPjvci/wZe4AB2hTl3xg1kxR8j5shANGZVXnuKV5k6thqplnxwPcqE
aHIy5Ev81At9jUstNSGzDOVvH5Jb/uaYsBsUX+gl6xXGj3sW8uVd2MMLiu9+3z5c6DxTVhbM0w2C
UO/kK1G0U4nMQc3OihMktbAyDocSCGdpYlQV2xVCMoYxEblq57JrZdU41oRvi3AHdy+TBcaYMr14
ZggTyQJjrsowoKz5zkc37/9bvx1lBMSaZWNn7GIuHYjOL3zeLy/MUQe+R6ijWORwXe1UwhsEl0ay
XEK+cx/hezG+HOWHXMjOuC+KQDUhXwF6SAhEn+tw0UqKmPGlkOz7MnbSa8mzQmyOHDInJtzjfEiu
EBo9CCRbZUx6OpN+DETFyboP3UQyxknRpkYUWLDaTes/3b+DlKvJ0r5UHtPqdVltOZTkhrHo8+Ad
N/4ITpOHXnac/6QNpAqM22a+9LoCW6nmhmQaito94Jyq17phQyi6d2VEsI3uLxjcqAeeAePkN/T0
v3mG8eloeS0+JA9qCImGPbnNJtGSOfaZBFoq0laV8YODS0xPA1iKu2fTdL24kPoVnx7bUPCmC06e
tomPNGPiTyGt/wdgCAvBq3JWvsXv8o6h1GCdipgTdwynnVILMN6FFaODXzBpHZVLF1PmUa+xPJKG
EsLifIwCNwYMXIvSGV3n8+Of2+xY97fXlKDwVR6UxqCWqFhYynXT7Vq2VJYedV2VEPWAzei21MU5
xAxRZFZwR/Q7+1DtoHPrykEBJmndH4lVuEk9CFUU8/XHv36wlN1NCZPhmF4FQKNDhhYfEoPYOaWa
wJuiFLMFe+uaFkCOCortEiKfJdsZXlG3xbvRCqaPGKGRslU81sndJnTILLhRaKmtyxCpD03DU1y/
6tzJt7nJfT6mxWPfpnIDk3T2OFxuDa6Yg6K7C+GMrjoI3eYQWI/8VhoLfTzpZ6aCVKROPPwH3XDs
qEGZdy/TuPw3lMsYAsEHSAIf44OXMIqPjg6nYUxRA114xmm5RW3bjAm29jwp1nTyW2cOsIWA4stQ
t/Z7RjkRBEWaTLwfPvxS72AATwyWVHFqPIqtQqDBVhE2dbuSKu+olV7aJdUeWI9NfigoKD26lYsF
XBCv9mn1v+xHZmd1bvo10fQkFAfjrepAVmQr5Bec/s6wG6pWWyJQ+3PUasdCehPg7ct/WNfQrkg8
fz07ISQyxWa0sT0ktV1pvqFBlU7zM0luabjBd579idJUaEu2Cxyxe6vNZRyRwl5QtAjX+caEcYeV
JknmThCTc7zWQPkdZskVHR7hMARx5dW3OK5jPdKAbWWwueI7ZaHdjZ8z0R9FO5AkrPW8PnBsT/qA
kVvboNjeERT4Q6MsrrJ7y0Q+ZBG7Iaf8HdeyrxmBUr4KDTaOl5fSPgVgB8A21wJcWivkcA689MVh
1KCTpb+GAT/EXFImYnXOLugyvuw1eoJG4+9EAZO45Dn5pnxEB+7L7i6bv2pmtaQJ4HIfZwizI/ze
tRWSOpDfwCfMCvJ2fvO87n+CVuc3BNiBJVhGRVSFraQD7+597g8vyWyL6+tgvQ9MXIZW9Y++G5nr
czFO2T4f+W8MFdn3Gsbz0qaaFEjz0fU/kVc1suAJaocU/ulfJiyNp221OFr/3MwRgskMtIM7YT8V
Uo0TRAuJ7LaXOGATjdofDPpKwb97BJ7vB0mpFFib9sqoAr0SkFYZG370U6Ep+fCYMUNJ3xB+CXh/
9FmoeubcLUAmBWT455n4hh/Jg+SnhNtDoFiEXA3cfcA5XP8n53t3tsuYe9tIUHkvH7fW9a5zLo/K
PDs6UaNyn9qOLQ3gZjie3MIF1A0QpIwm1Mu63pCXww1BinQ4ra1QPpXIIx7nQp/PwNvB0W8vfjhO
JBdZ7oZFD2aRPXRL1BUkCijX6iIA5AHsg0siHr2EiTscxK2RdMCsJe3eucI4J1wOS+QChi2vTXY8
4tigvu+lsDhCnEKFPVVQUfNs0+vCIXFYj9xBZTdeeKmqYQyex3u9p1RoJkOjB5VPQNXNjpkIviiS
eTWGVVm9+NQpF38F+PiN1UynZ3m/bAq0S3t9hn9UP7GXdeuGMKeD5FlnlTTNGds4rCP/dyaQXIRN
pDKQ+8KkKSIkgfLGhbzpQexgStsTVfi3As7WU/mR4hwhoh5LJ2SzWKlF8p0KBjcC0f6xa4r2cb7M
fvuzxVaSqdeKPQduyc9YpjgbUVKVtmD/dUiMy/KEegkjHxu1bRsO/Yd61n/odS8E1+z6GrtUU3+y
+M/VZTBFIUhrhhG/7nAsYMniVq+YG1XLdD8N6T3Kb1ZGcYLJ04iOiPy2q0AzemkkApljm7nUBoh+
CVqbh49xxVPqYpXjvyawobOi9fiWSYb8iQBAkdkRoUoXKSf1npLoS9i+jBBIbF+z4LoDkhsRA57Y
TaBk954LjQT/LYakD/uvCVS2mSk5Qwh7RaRDBzwpyoMHDmWJcJEDiyCA4IxuFR+s+Y14y0prfd4A
yZ0IUL4N0Iy3KQIUOhcbZJXpuaFMsMJMTE9db3jLzwNpfHiea93wAzi3g04Dq9U7omg22hWpRAKv
5gi22kRzyeFaEtPEUYFtl9CpzIU2T05Ta+uB+n3Tn4AvISATSG9n4Y6JFsXrxPIg8n+szS8oj2K/
VSgBY+ytTsNbqXLJlaProC2iYUoJai9Llvs9QzYsRaSr1p7Vk0yn8H8tRCWjiwn4GkSklje+/rvS
7bg9eLJPEL+u7d+PSqnSPQ1ObXeBC7c3Txna9EHW98V1an+BF+Byr7BhXNHl/TIB30ToXcOE/pJM
rxmajG0TLWlPwqIta83BsVb2FqN6DkiQuq0AKBNC+NpWTEhYA8lN+Am259j4Wy36xl965edZl5Mu
AxZ75l+1fcVR3U0NocNPN2nTZyTq9X1NnQjiv0DWUm8jselHmVtlQwplblh3wfU3KLv8egCEb7JD
7qyMMVTBeEU8c2vOc2tVp2BTev/mzcefngacXv4VtPYJihBEcVma88RYAIV3v1GsY3HFGaNqcSsy
i4rnuuxTFCuQNdZ4vuvbvfIbUD8awjiOATQEa79tkq7CMq8zFz2dNEn/iYn4V7MnbS3sQzDFa+mc
zv1K8I6g058QVZRGJs/W3Mvd8C4/5tgm5iKwzAw+0M7h1QZsLzc007PX4im1ua5Df5AEvCPUPFaN
pWsPTgqBBU+5NPOSZCmW3Y19jmqS43QTW4xFOJc7yfmhisQGUg1BXfV8ekr6tnIyAreKuItI+G5V
INhVzC4AD7h/mpAWJ3Wyma5BWgLoHohm12eUtVMdunywee+o5i8E59tWkW3Wd1GZEizvPOIILvun
Bb7YRdu0RrhAHjkIsh4TcGcqWx/Jz7HLpYC6MajuqG5hT5zErFSQL8FVKWdoV4ir2sy2QYXl8sc3
ATQ7C3wH5RZeCYrxV0fBJ1j0MW635iVpo4/QqXjttwRUlHWfbcJIPY8MVDW8+IxC1T5X1s9RUSkH
3Lzbu4X/HSGLpvOfffNnWaIY7EaASSLKuKp6LyYFoql2ExFjZbsWIX2eXjAbrT3acYZ8y+6y3/t9
EMgv/Be1Ul6l4CiiVQwF6hiyR6NGsSAucxRMggcVvo01yDaLMiLFmAhhd2YK5UuLW0Ubm8hhfLay
dMQ0n2bzqwZl81EXFpM6NJk1Ww47DsCQE3ESWjG44nog3t/uJ8BrJnpsQYdaa2PUlsJyNSeOhXpt
MGo1aqa41JhxDimE/m23m6Ihe9mbCJRlGifWhuYoRFIaiQPoCLuYkvvvhABaDW4uPOlz0Whx5m9w
1e097Z1wMv87S7FJGMHPlJ3Dh2AZ2qSxlZLxM8YSiUbUlIm3+M/zErRhqMndak7SP2pXp9g7A2rV
5EBoDV8zKB1j+6UrmcL1lprjFzy/iOqWdM9OxWy/LmbXXHhTphsKaWFMhFlJcrKLNr88DRi/IJHA
FD2ogLxjqKXodyYky+MwUy5wQqB553zwiB1mEccFhquGZ0n7WPJawglfl1vX/6l/LYpUqm/xw1BU
oyAFuM9QE8W0/KeE5aO14RNEAvLNx5vFCVpFz02SIcWV3Yqa43aLFAbf8cQZ7fMMxkBcnqmiTVSo
NSDzrpOaefIUfa/snHe3pPjRfDfFauQvYX6kqO4mqA9E83FLQADDW8n7eBDJQ6q6ooCN40WF/Xzl
bSIs00Amu2ROF5FO4vskxtK+C+V/YGz/P21EGvYSfHL7+UIukWLJ/x1vYkKKMIHfJ5eHlgCOy596
4vAphIIlfp+qY63lw6ak0iNA0Z1CwOaHI8u51Xx6hnA88VzMMV+8dL1erzYFnvLEteokjHkgFAcO
xZzX04dI7qOM2JlC3vE5brxU+CNTTa3jz4tS8Of3w3iv6UikZaIeHJB4slTN/jrPEXGr48wnUIJJ
f8ZSviSbNzw2khTe0M+uuPQNHWD399q18hwLu5KXu5NlSsYgwmOYfR/KY3JItLnaXGEaXFhOsbB8
RZiQG8lAAw9Q9ZbdVXElHrDFxklecQbp6smZvIGQoBpsDoLpHUu73WN6b56LeIzjzjdLKLhSMiZu
3BjG7PC9U+LA95IJTM2Jlhw5f2t1+uQIawmGZHGkqTw4Vy7QUqYqXfGwFmsYtTXefRQD5GGYyIHW
yJL1FjElZosOCt8+mzCdRRkcWwtQ3Vz0CRG5U1guT5ZZ4XjG7ZgpM2VZQBkf68SSvLttJPUIdydv
pCQSap6cFR8LMI3PZKbwKAMQ9kEEGuU1AxWbDyoK+zv3+C8RL4aU8EoY3HANPOFit2IgrXX28tox
lOFQNc2EonkqlqMT3r2wWDZWq6wA596xcV7us5om/pvorNyZrSQLf67aYnnurfAJwKl0GeICO5oL
t/Vc8IZMMFKhUn81eyH+FkOa3+nW6YuR8uwJQ/mxYp50jqSr/RAE8NQ1xBN7/Xhzq8IuYm463YZJ
B23AYn6Ol5StBu5jnDFYp8YNhaT9LmIDZnrGqXSEvGrIMiYnuSERIopXODpgpcwfYmvglIu1AFrV
Z+avsCF2qPBtkkpx0eMwf+EOpJcLITXlfl8sh2YYvgHsnCeumi0VylpkfN4pvAo0opq0odfbPLsE
8SdskLdkUrB91/7hzEZfMcKuAOHtmi6sYVcRJ+SPZtgQV3b1aGQkb0eAGfliZS6QOpCVJbb21jYZ
v4ZxfmoQMW/jm/iMPLFDo//4pPu88G5KpW+3hchjGrIuBpfT/XkXYtz5+qrkQCL7QPmUuWYzNOJ5
F/ZWrz8fDVlcQ7PcmBnAg+fPoEKQlt8Z75FcBEfZJwQqq1VChyu+4lQjhL0CqVMAji3PGOM2DCzz
RtXkT5Z6meqP+3bBH08iUap7G6c7dkE7MDufadwU5AQtAQfV6BLMZRTByQbYGgo/bE2MCyovUgNI
rNuMQo9AFuYc2zu2Q6ute9PdRhH//66nPjW4EwCUi8lxijiOPcg1EF9l2Ka8H2ZTqbwdKsuxlIiZ
H4bBHdGP9ilEIi0j93Jb5Pc2BBNPrFvZPgXn+TDDo59fQ44pINAdaqeNs/LikEw/bk386lip6R4o
avjBajOzwqhw1/tnajsdze56PcjP7KDlLSUYv6Alh8u63rEtqeFE435rjrUlVt7vPjPWIOoplscM
hUX3JBtdZgqKNnvFn7g9llWSmHlHPYYiCxs0k8YOnDHJ6avOjRqBLJHeOtrami3cTs0f3CzkytES
er/oTRfTcam4zbD8iHFL9q/CVKJ4JcnAiiAfgT164d91HH2us2VzOATsP8BBwD93zfqDZJd/uWyl
kQIlNbWtEkQPlb4IXQHbYbwYW3PYzLrxpwQgGS8PLm6N6tFS83fvu55vGiaf+Oy8s0GlJ6R/VRRX
eecqNPxhHIg6VO8/7utzZ6YIb0pPzYRXhHTyUgYPgwJHQSRNpKhR8I6lfvy5UMVjZDY9A0iBC7uW
6Z9EKvXb2hC1yZtqUV0xgQfI1EFfeDDdt7Dxv0dUt79e3bqRJJ3oA8dgELdmAAwlvHHqJMKLDO8O
+LwFv3qkeRw3LSXluI95VfNXUX3R0w8OzOnYDqFbLxp+fU8KO+/7iA3MzMsD49xvYkzR6zRwcB5L
jTBad5SsxQk4aAIGIRgqsmg4Gbi84wAyDBgKewSaxNf1v8+r4QIr5udHnYK6TtDziXT0yIoOP1q2
qNif6mks924FckGVoPZekM96W5USKfYgQDXEJnG2H0pG+NWDauLbeS1SuEmVvl1Wqv2nl0jLV3mi
+aHyG95Mk+IXFtyXqekMbxLfjnIVY99DehJdPcZQp4prR6EJEXD6aPwD6T5AFkrjdcUpAKAriiOK
JzZKICbsQOwx5Taqa1A/6DIh6PDupCH4mz1TAqgQ3nnMqknQzzXzXKoJL4u1j3jGv4PvsUdkaqsS
CEwe9yhS0naO4WVXoWY1GdSkdXqiYJaQuzY5dYrgF6nGKzVKNqNiXZeDgYWolWdeqAYTUsjlvwnZ
FnrD0QdNjVCwamVauWga4xT1g1iyRXbXCgg/An7aJW0D1KFj0VB4kGNWOjZf5fUYn84jdQNwAWR3
ZzWH78YutCDw0c7fyTT3wfKqlpB89KkVmv7Krg+tafsbcsnkHlskc7MnG3yy49f3TmNiyFYvXqC7
cxYL5f/momi5mwMsLO14GbuUSLoHLOK6vxwsdjJiG5xvErff8pY4pvt0YBiWKu4lchgJOj5j9SgL
Uu7r8eqj2d6h3O6D2swKBKW+uuAuVlmEeKkb6/jCyfRAD0zLiGdsqckYOU1qHVeS1CvZO+OWSu7x
Br6HxcNvc91yuHRHHnstUvin6E7PKlNOp/fFddRgHpVu47y2hV6beM/iM35V/Hl0ekhKN44rlvfS
Cz/cCmlWOi20zOb+9JqOTqgy7T5+DyTECHRsALZfNZkt4PRqazGglZDVanO3zw0WaUk/wgVMqwDZ
nWZTr6qliqbBsR+0QgiGjboRB9mQRxa50j8pBJPpGPxe1MbQMgG/N+Q2ug9VuSEu5OxBJPug/Kcd
SFZEKy/0yUq0B6+qZw9ptqbVgl86yPO8dCLeRUkMpaiFntcpAGyp7B11Hklfyfe5Xbc20GJp/d4S
pGcBb6EQvng/jqA0nZFwaFVyuXv77XFPveT081FLf3b6kjLocRtVNClVQynYmMHpXnGQdRWOnyf+
xdCsjV3e959iayiZ9RCirrD4aUz0RDYt2kY6nURNvF4le/ETfmN0H4koN6cnWu5aHhIE9IWnbrzU
3wggPiZKQXRTctGdQa/HQJ1LzaxOi12FYKD+AJtEunqtTxxDGxQrdZRjukPjhD2g5z7rf1k/MLNE
aCmEHmkT9v/hbNuregsDVsXj0MIGb5HA5r04A/hF0KTKywOTztgBVkXGxKVHqGxqS5+qS9JZy7kH
UZtzKI0RZ5xWEZaCiZr/l2fjxZMSZeVi7r30CuWC3gyQ0DJlVmgfb8q8K5Cd+BlpQsFhqRxIDHPu
AkRAtU4Lq+JtCtgdsue3WuSAeE97mkkzCmPA6dHfysSWOgNkvYz+8xQTNJXAbg88/brRfHCob3Ic
BrN7C8LPkcjT7QyBlKUC19TgeJKAEYbfHIpuCDZWkqOTs/JAvPxpt5wXvkAVp5FrK/zx+wglO4te
RwaZccm4v1bn0MsTrCWAtR5ZflxVbaE5CSsQAMO6wpx/przA1NjaF8b7Pl6gAq4O/Ohi0LO76Toz
mC4M+nnSgaMpo7UeAh7eZ4+sFWz3eYNpMLbZl64Gg9V3LcLP6BFY/AKLrfkjOwnGqrX0XaAW+GjN
qPZEiiB77WZY5KCJuYilu2scthJl5WsyotmVgwgeGpxvrG0aC2/xoZo4AH0og+9kK1ef85j88D3B
AtEPw6tI+5EWrcPlcqMngd+2cb3x/Rq977ZJdTo7FUJg7rj2PqixDyxD5yvFeobOkG0Qzp68KZs1
hP3HoEfby9O8hBzUfTgxt/SZ/WmJvHDG02t3Wj2GksEJr7fnAOvx3w9TcxRLG+uTr8MDcOumrWBA
peGTu7PVlDbQTEqQN+5OQCj83b9HoxvZYONjen4vcaCRWfRw1l78LNZFZ5y+UZTEWh6JiB1J11i4
x/n3uh41LQdGqRmX7N4WD+BadzdZVR2YGxMsZZBWg5LNrWwmk5pIIqJjL5ORX2UDi0dro4BlMngi
Mgv7JmwyYop6fumvMYT8qu/ga8RhwmDha6rMB0MNdoE6FWBoMd8CbglL6bU1X2BDgHSyiKSMmKZE
UrydF8YuSAw6bEXbbXDrogLwP/bfyP02Z06j029F5Gig40WjZ86YnPFy1K9S0M3DqVs2NYJCDhb/
+VoN2bOQ37J0HxA9+KjcYWx6fJck0tuLQYRmQL+6sglJPIGv3EgDvrZDvbBdF3KW7ZoJCeiHmNOJ
Wgf1tqICMYvgEg2ozpxvpALCLX0WP0hpPWY6koUv2NgemKQ0LYV2XGo/iqMCO3xfRlQ/b1qNqpj6
mVUgIiQwygN47mjssvMkdeFGBwIb3LBU1q4yPJw0mcNz9M2K9TrArhhkj4BpR22bQT3U/Wn/fWay
Tj+FW7TNqLQMVpLjh8tFvh20lOnWBxqN2r0+lQinhZXcj2pxTjCpr0BO8tcEflhGlx2/gF2I1pbM
irtkKPAQHjYT8BCWQFpWK4gXZJ0iXaMKbBXLtH89rYr1fO2w4DQy2nPYW4btEbmBdC52LoI7/aOM
qsCqcU6En4pHGApHBcIgKpWhAUV4azGCslEieFoGrQDKwvdsRBhaYWJmTqgCMRQKdeSgD7TItsaF
f/PZoeyUyloJ7TlKEA7heUR0KtZdPkLSJXFep3Ma++1Y6eqNOEInC1jGEIuf5DpZrpLz2p/vVZnf
49eTiNrVJIf8gA2WqVBzIa8bt3xc2tgf7PAqM0CY3nse2iBAqdg/KbfYJByLNc1e2qupj9PJjiU9
V4EBILA0o56P12292ZqPMv80AGTgytSLP5U4cr2E00unc232pYMNMJFS5ecJmBzkXoCSjwxZvrwg
EFU0SAOYW+a25yTvPq9DZFG7HO/DeGOHayl0K+TfbnLsh9Cfxvfw0NZvEZNFyvnoBxmuC4+/3aS5
7I7VdZ6kzgJXiluPqBsuVxZbyNM1aVrKTDf4nOjSjWgYR/0ZEcpryQ9mtTff91QJAN0ql+ZekkdD
ZdRXV00gdXxvMHz+oHeTqR78NcgAGIW/zxLd04HCdv4+cIZDhxcdmBDHH1oLw4jCDIXtmf4T74lv
ht4LAmweU5pqA5yrHq9XUaqRRBeUIl5vmUl+cW5trc5uahSSoHUNDg6/d9Rh5jVlcStrSw4g5wnq
GPRE7j233V2RkTpSkTgb0XvIqhrHYidiIZneRN2T/14mhgJuMOsIU7AYHfMajeBl65krilYRHsGL
CBuVukaXKciMDP4WKH/OVh+N4Ww1TC0GwceqwEpjhD6GI1wseW+vRUaPAmtmidP7OlXdDY07AljM
Lun2wxW6AvdsXwGAt3lg+/sTbNN9mcIL7kEEgt8QWQuA8b5BVTIz6nj0pl/WWUqk0eSin4NeiV68
cjLg0UruK6SS5nExb0zTPMSxPfBs7V6aY0/6UMRdFn2n0hgkOrBLgHZhgcwL52pkyUsP63Fffrlb
eDj9UQ47CYoiyjCuUWJ8utWPBMU03rw7MRNlSSIXwbPwdN7avhfEpUV9pC1WafMoccCeuOXu9P4Y
yClWuwskLV97ShCEE7zrZCiXhg/sk8uDSVmehUOKLfMZeqHGLlzO2xxTYGmiENa0Rr+SQbh7QCYM
YTzAfOLRy7ylboa7nUaW5GydBZMEATElHh14B+DKeWNwaXCiVC3sGj84so3SK7rEjh5anQBOw+Oa
1scYL9tACfKYcHNehre9t8z8zuzrq4wb38iqpYTfP5RS8hcxUDktkv2Kj5dZmUYm1GXqLOQdnng0
eSf3aXNbWRknnn+g7IyLi+V29QUfP+8tzm+ED0Hm+oouevQ2BV1J7Xm08luTf4lbnB94V7Rtchaf
WawMhbDQmwcILKL2eBlOamqgJk8x4uUKIm6zmV+RQjLopRNxdO6hmIIN4ETfaJ34vz9Vc6dbb7nJ
x8WP1ue5d9NbB55wl0aEnEFAYjca6D0GW9eMRJ4ShK4NDq9Gums5NKwK+XmZYrheQ8BpqUQrnRao
itnr+zo1+ALDXKVjS7hK3Ir73JvY8rLZPui0Zm/glua3UbM5tlVnE/XWs71BGaqIU+mkwJgEEgWC
WFkOy6+osLFNsc7bJWGi2zJUka8oo8foKQO0L++DgRhLi07FsjshO3e/E10EVeqEUyGCZPUsbZyB
TlHwV4Vkf+GT8At/EswHvaEoOM5kHuSRGUcsAJq+OX1TAQO2TJHR0Xxv698gDjy59KF1B+fhWPnw
+Dx1lbHD7biswcCQQyO5DzqUa9cU1IPe2lRVK+SR4kf4oTw8RllkfqlF9pwI6Lbp5msmlafh7h2f
97zcO1aeHz7n+k2DoaLxx31AoBdm/u/a31lMWro6fvEnUiPz9bDNeEErIP0Gr/gauPalvs+6rd+f
kgf2VzVGAEfWtge6YZvm0y43VHrRhxhbhAnhP9nn+eNctYYDEh2jo90rh7zPUdGuvoioYJcG1s6Z
wnV9YNYMlLBkvR+p4uXWfft7ie2HqJJFrKHQQo1ia6+YFV6lRmKumeuwz4Bc4loGmQbnFptCgffg
Y0ZLfsY6wIGnYSa3CkgkxKgKuUA1Attt7oCxYp43qmgWLgTrBCCGztpJC0i8NfZpG+rDXOKSXa3o
eyll71jzktsGT//fGeeUkRplHeQy8xlidhWjN4XCjkVJhu9EKGykl12gdCSvWF4amH3f+4Eg7XWk
GbuloPResEPS3/AYiOv5fnwVcm+H/bujSd3XNHRXA00NbaOyKpciRRzKWhDDkovHdzbQZSc1eJqS
lthvA6v/E2DE+DueljSAC+QZBrTCy3n/gceek5eFlRzh5FUUrMULY1mC/kXQ2jfgl7ylT9wwE4f2
R0KtuCd427xY/TZ2nH6fLri4mssYvQ7gBG16HKAI7j2A9+CBT82lKLCwC2xiKRPguRyotcKnof8o
FgZmNCUJtxnKwLEqlnCbPtK4wtCNeEtpJNk/zNwuWOCBJC1bTcMWxRk4/UEyVyJqhg6dIHO0hAZZ
3JCWhwdpIJ1JEjput05e8Ruv/Yi4ZBDJ86euzBAMoa4WJoW59bZ9MsMQ8oMNk4V3JG6KQBgWQcGL
ebYc2Aqz6Gm5wTF3NAM8F1s5SOYMwIjwSJ4QnoLFg7njVQt1qJvVPrg/iHkvXgum4+DvzuV4tvDk
33iTdRpELYFm+JustoZNDldwVQKQvz4HqTY3dDkv4s5Rlf+kjNTSpxy0Np+KjcDtXD3PuUBWr8cW
No6dHAj5BB92KCj4i20JuiH3zUXqrO5rGxD3uNawmkzvJgFCPxYjGQfeIxkUwVMQg8iww93mvUGF
HauzvPzjO/vDSO/EI7o8lm459bP/E5SnW0wNmwFMzvuO1EAhjSNFHCvIQm/PqwfHspQ6istxsr56
ZkW3tn5XKdHq1zZ8I1UUHaUpeibmRz08RwsjV5mSk8vhT49WD77zyk58ll9W8UR9GJcAhuCx14k4
tbzzpqFk67SwMQevWvjJ7y6VQqttMxY82tGYdM9g/McTDaYg/tFFRMPAvbQEJoMfGNCsR2uDPsOQ
jORPjqe6fTLmQHldZJtl+XKUb2J8ky7KiVumhiu7n2lo0r6Zup+J+9zcv2glrQqN2Yvfs9+5Jn6U
g9L69U066Pl/kGmEUNHRhq5qBpM/bjH1YX5i+y4MEVgcNiOSTxeIB8dMkqAe+CeTgPwBR0PrJATN
MV2AW34CIPDS8weaXxWseeOJiQhHf+7qPkSpYQNJGBzeDdpgfkjXMaYvOxIROFVswFCr8QD8tYQN
asF7ydr2SVaJA4Ikl4AmP1KSuvnv28iWhNzpD8mbjCyFaZzUApz1s2N2GJKKkXGhcZsf3efOOK2K
0oUqFWW1GGebc1BLdEfL9KYP7S1y3mQHDg1lcxeiv0Q3ifWub84mF8l5qlfNO19v9O680gUZ3WKg
0o70+zihZyI+JSdliiL3HPRqyX5/20Z/iqFYFnSDswaHzu6V3IsQZISGt3e9jjPtNwszmDqKX8Z8
7kKCUelsBtJfw0GG2jMqE9yX7RmTsxbEdbLqmR4xgmTGdQP0/KjNmjyc9tRzaFQtANAcPq5m4Pvu
SJyiJImxfTJ69Ve986mLyHUn00pqS3DFfKmeSoz0q6uhasStW1HFkxAdz7SL+kS9K3M4nmAlDz0I
GlbSSE1EfKPzjyN9Mt8u70LDlFuUMxqqI0szg+gV9ELquEwNOOK+LuRBIjo2ANU+o0EtC1gCjnuA
jy+pZjkB7O634RE4Ks3s7o04oWxK24AlUim3DAZwGvvWCQrjMrWe4bnYcHNh4nB/ChCkz1MLCNpw
49VdXVZngvJzhQAyROlwls7FNanegv+xYzpU7ifEKQXpzQfqoflXvJddMislTglMf3rmH1kuyBGg
jsjGOgfgLc54Kplg1/zenV4ewDtfYh1fZM1G2k4tQudtYFPMgDDmMvK9xovEe3Aj5ZTzst5fY1ii
01/KUEMF8On1sdyeYFqpuVXECd9aZ8Lwwq7/9JrRVF3ogBhh1xQmxm1ssAa1fPCcsZTito4YAyc2
1jXmLoUYIro476ufYETnUJ7A9utQMRtzkCHENrYslbUjBevkibRM9gcydlRmPxTY12n6KwwaAWNj
wjzHTFHPr8eXlTTksRITg1vjagsdiya5t1JI6plVcFirpKXoUnVUo8uHe/0+WWinxnElyhiXuFrE
P4LJPgINi0SCY+hD1TxcOJihbJ48d5CCmN3WKJ/62dNqD6HwDNAf+Qw/X/zFUDewUcAnRo5dNdq+
wD4oBBE2c0gMTJXEFcKpgZd5Uo3dXhzIjeAfMnN7A/6MObSIIcY/+O+0TJ74MHv8MXBkjH3Zsj6R
Eq8N8iPBX/Eu8hfUwufUUlV9w0mlEkLH1gvDfSt1VfQBjffvRIVCBkmgQRpkr/v7Uh6tfaDUCHTX
Bf7WwvwrFnviZWet5yb9Uj+MWv8G7h+6+e85PF6XR2XrMsbMX8e9sI5Qo8NuA6pqVNHMaHPeDv1u
yf+iAIZIiW6FD5crTjLPW57LJt811Rb45Vpe7XqKQJkavUQedFZHfNgdIsgrJNdGOi1k5N+tHTgb
00ix1HRSOYwZCetCcuHYKdmMTIOA0x9VHp7TdKWX/LeDleNdPRYXxMi5uNeqh1olFJjCTGt70AQs
yi4qXIN/+Va/Orr0XbBlQl1dSyw2Y+WW7DVdA9Aah+JYcgVLheFveBQj9gNZgSeKCzNqjmXP3Dv9
NRhQK808Xo21FTMUp57sA2WBS0LPQNGnN79EwlGQFApNsMniz26yeG+XmFZtHXIqzlGpn909fLDC
ShlGAwKlEcCKRX0tOg7Z84Zr2o6Rol6gvqKgsT8G+rCVLihhgEjmngzhflVMDzV9JwDDTXgIGQUC
a8yUHHWAtNYq8zMrp8ZLzdRTaSF+gjRZmjwasGKRjEIKfdBWzU5yHfJwAQsomsF4eforN/4bP/3P
gxDLYwtNp7aHS9kOF7V4dZQOooKgcZph/rJbIVDOgjZx+sQ70vNQHUFyFL1KoAJP9NlI+8gHWW9f
XS2iGoit2rQi/kOk/vpNPXTuAtszeUEpijLHuUPSS1gvI3y02rQKSq0Ex+BvXjw/Eeghe/ZZBf7e
9wiR6Nnc3GK5hrufRvCNjzmiJwqS8HIIbmtuRpQ/WfduJkJMXt6lmlKpaupQUnP6I4O1il2hF5M/
cRlLqoJHWWnqMt6MlMkGDGyYylvSbw1e7LcHk/OeVblDGj93THyIs3+XZojYkHx0xlqrBwL6dbrW
IICLmVTa3y28G0qmeCko6eaQ5Wuh5T/IVLqTkdun8cVhTHgoL7Z1t5AYrq4OHxR5n56oGh9kjxX8
28kRQtGWq45PiqvQKE7P5acLcw7krlwVilphaEbgj+/aIf8OC624FDemzOi19XtNfN47UiKqJE8f
jKskXGDsRqc73VpEYIqep+jn8GEE8Cs8ud91NqEwbWbPWxdtYIJ/HQIBLJvyTVUn/5BQ/rASocSO
dCCqD/4ibHuXKcSegVNLZ7DcAxwi52lyFCg1025cMPEu8gRJxh0SFKJkfqWUB1TeAjTqPdR2nma2
1IPm0d96R2K2ayZ1sGUoAmQ7Av0+kfqmBKw5mQCMAUC8xMPYncdrGTpUvuRVlDEzlPvRVZUpx2Fb
I9tHUvPnqxMoD50ZEKu/BQ9fabyRZKTD8IdyhfpC0No9iDpMsaLvycPkcB/VMt8a6QrsdbR3uU72
OTl80q36YG3ZcnZPl/TrGrlfJe3Wmfa7iGorzuAY09+IEz1PXDoy7FVvfK8Rcm/HrcE2fr6/9JXm
lJ+AdIVS0lBdGh2kdMqqUyM421gLWgiK/plUJL/ieMUOS90zyoceOxssV+oiaw4PwZpwdfYqijuX
232EnuRo75nxEYJxIKD/4oOX2j/njNnPpZXYp3x63Wm/UfURdliBe3tpg1waey2gZH16l8MhGvFr
0D9WHT3RCnfo1TIi+3NQed3vN6VyuWrKEUMPljzIfBzcoCUkGT4t7y/+2O8qr30R8ghUkRrb4Aqz
+nTUWCN7vM/9xby8MJ/xw8Ns9Ivk8+JxRTSs5dCGBXARi/rNZI1v3CZqf0/ugnZWGdX0ifQqu75h
Lo9C+GRtwMqwXtjcDgN+0s/mJBP7+PMYdfeppkp6diPAUgNk6PaxENiAotwfiBKoJ+WcBoCoz0iZ
zU7imCi3RvuJ5txoGM9syUzbN4kckulSKzWt7frMFcO9bVnL3k2aAo45dcBzrCrnxSf4Oe4yTZYj
iR/7t8+Gahuj5gHiMD9ZKUNR+HKoG6mZYpRmQch2mZjRFrFqug75MSuXgN1p5mbT4fUcaArHpP/l
uqRVqejM1XexQHjb8MhXevsGx95VSJIPxIiBbkHAxBFYaxNTwvqbMAMiGOsO3ewnbO/LqkxivuXS
UvAuCbDN0senbJnycIAZsCM3vcI53KyBTBXaoX1kHj+NyF3A7Ex18KxUTdLb/J3IsMyOjaluN9/l
IvTk6WhgtGiN9//l6c//WvP2V7rxeQwdpWpTUXTvBzV54kXMdgeawyE38lMDhZm2UKMth3IQ4Ue9
7frnE/hk+k4180L69nZmBqgv3uhAx4K5Y23jFgcdxQIwA9efL2/Og42y5SGPQUVffQgAykQ5HxOD
wD9px3I3I1/Hifq7dm3S5EZFZwWE9m/8hsfiehoblLwBSqZcbdE3gAyEP8xdj9UT2o3xxuzVPiy1
bkrV+9zfXJsrnRgM6AiLAZRs00RNmMSMihD3fYw4ZAIC5zHo9UDg3J+NuEkCiHJVC66EJ5W5R44c
TJnJrwDkY2XFx13CJXQM4htbeDSlGhId+lZ797d5WsIAmptdpe1emxgjiFYeBhPGXuEBoK9va5vM
KEUJiNzAt/5rz+A+R86jBM6klp/luj9Rop0knwqCRRh4up7pPaJaduaiZcC+cRHqmg/pqsJGMT8I
TnWlOlyyFOIiV4i4nTpAX6zaEm53UPr3PncooW+v47D2Rwg2ONcCdDjpAZDB+dtX0mJ6lmTSXpUB
vnm4hTZK1ckS89yRhSM3Kggb38qT7QfQxP3hm5jjWcxJWMM9INJxLBA7ieAWn/Yr8bglIp7WZuu4
s1rvA6BuXGkSjos4Zn+P10ju9lyFECfi2n5TLg1PwaihCyNtJJlXxELCt4NzUJ+g5mD8z1AY4KI0
tMpzQvwb6tVvgOOf779Gd05PDGKo/DFodG/4vrVNH4S1eEnG73yeVQJ5mp/4d6e8DCEtqRrwwTLY
HrBxVCn4Rmtq/w24r0frEksunv1hv2mpcTAy8GQN6LPy56dJE70IR8l1a4RVBvKJz3XLKX05ORfX
wgFVGzh+cIrnMXUTn+Z7CfVGwAURWmlLRJCLi/RvVNvamYU7D60I3A/HX9mJBj9F+lb5XAAICqoV
UEwXfFdnlf2JTvGq7sGYwqfdxhlWtIzZq7cj0I13cTDX3KUBeDBMyisXL9Pa+F5JkpV1eJAB6RRl
zh+tTAM+D0WYzUBWC5Z391MgdT0746/oZ0d4wKrRuuO0Buf9HeThv7U1Af0b97Zsr9Ac+pOtQ32B
SDvjNa28Q+auwK0P5xKNZUTccF5jEJQeje6zaQIVUG/ZtIV+TOcJLhwu7+Q5TKLfMmlyNy4X0SPH
aBqZfD6wXAKUY+816ICse1J+FtpRzRqJibEP8JZi4QU3QitcDFeG5DaER82C/4UjHtLwitoAstkC
KVBELMl4GlchpGI75HqqQF7Wu02wnyTXiqWCdns19Wr+oC0rJlK6cA1uxF8W7voZDy02XG48a4wp
LZDwnLoRui5Bqx3CwHd6Kp3nefYQl05Svu2GIvMLkuv3aRlUXnSNEYUFlK6z5thAv2eZ8Hx0RJXq
At2tUJWOnjts9+IY3jGYUOFKKFABDkDLn5SMPfYi173m9G7S8mOB6yphMt21+7V5ltZxb5Zt1dCa
sAGu3ztYh35vgNu6nPdSfG5IkkOLl6BKScT8uEUHWIrCEnX2w9QnuOrbQpVxYR+lXv9k8BEOPB8O
3VLysX0lK2gPRlH5GAymDIHSUd2xi64D9LclUzS0vGpyDJ4BNbR2qLPi68d0pFeHJ6D7EXPkpUlL
GjOEVzQpJEXEAxbm7ChNI1Eq/B4yeWLfM732kddBu3xUHvhYfy/xuDvoSe94pH/umKybAM8bmDND
/OcqWuDRN7oa48z6OzBXoGbgrjBIANEqtnyUmhbRLvcv5GaqPsbRWALxmIeElR0tCHngRxmK1Xop
7HJfrSIubzdo2XPK7DLyfYk/blv1NTY/KvaOvP4XIkZVch/9kS/8DXoJrDb2HPWqU/d7339Jy7/W
Trx6T30E8msl6JVWN4uU0n6MY7dMlK/PFEucW5ie4SrGG3TqrGhAWCmmixSIN3JJCNtZw41JtB5b
FE0jFioHedfBgu4l9rELbmlZJAU1yzRrov5QI2OzjtR8j6KJoE2zuf1dZ068BvQmDew9VVQ0EQdh
PRShnB0crqns5cnGYmaCUqjHuBZlZxY58fPDsguYO3P3oHqnzcfj2N2ckmIhfSYXkask1jHFKnG0
I/1ovsB4qPZBN2iHX5L0/lXcXx20qQKrcq72AoFERfWF7JmBOs4gyFDhQ0L70H4vVhovOjMecR1e
z6dW0ClRHw2N8TbClGlMxsEFWQddNzEAAzHWKbB/N/3zitJPX1DfB6ErkBy4JSjPw8FE3PqFMIds
rq6u3TDXasTjT9Sem7m2XvSzK+/uyJerRTNfv1FvdGcd5ZeD8XNs7XBqX6JUazZV611xLLQuAd7J
8PKjKRF07DkzrkMZgz6zGuhhU3/7er1ffJl7a2M+MwisjUvPKvFVHfqeBRWqdMqdVORypUScSYw1
/vClbgp8EjDc1eING87vbty5ZgJ/euzd3TCHQ6xDjdKO66SuEz5IjSt8mUWQVykSSOkSZGA3z9Re
MXpKpLmHXOQiimQSsi5YViRYmIoR8iRTxni5zXHZ5J2mpt6tEK9Y0NL2D6USMF97UDu2+tsqheRP
UBxfoJGTPpWIUz5xZJSnEXWS8bJx7ZzocqxNvmGATD2+O6N5JkNe52KnlbL9zsliPUPvKzDYFsI0
4E7iJEva6daej9xlTQp+ueFGFLbXcXpv3KmzEbWrps7jwPbBCCP0JR6v4Mx+WkuOk76ytm0w76Sl
TH8WabdNnTONt8Eisfdf8Bbm67PtNu+scxCVEKb7a86p+R0+/PIoGCzXymkLHJbxpgieEmY3Kgrh
bhKj+GMyLw9MB9WCoV3txKVPROSeRiz2lDwSqb2m9qUBKHCJQ7yTfcr3hN6n5TtfijD/DIPQ6ODf
gKmWvMMYjssLdygHCuHPQuZJ/fMLw2cFuNOiDH7CfZDr9avcEG4MPO9/7Ufe0rrJoN/HuQKMFZL/
aZE5RE2nAgyOfVxOuLpu1aE6NBfDyR43z8uwvAbXOTSpBbp7QBgEQ0w6UusIFnnlIiE4KoZQ1ZOZ
YFuwQV9wZ+RtfLjgFsRXAqXwIiCK40U1sHSQQIqqSYOJwsH9BR09Ft/8PCEeapdBcDfpQa7CEqdj
HDmZaBgbEq38TLgT3pmNKH0lIBXzLV+wRwI6mD1whai7Rpjg0dnKoYLubpGDNsinGIxmrAcRZwvE
GsT0DcZGE5YVvA+2ptbkcRjoY+LMxjpzu05i9WXh6cDnzqawrRJJjRvQtPVGwlvRv18s+D2OzMJT
NWsWYTKBCL+4rxiGAeD3gvP/YBmiOIgu+dFhJ/P4BfUE98CqtiYJpNypc2nDmUvCJi91Cvd3SP4+
pVI0X55ITcmCkNiWCihhU6O3K9GSK689w/v3J72M2l6HiKox66iS3yzOyvGglLIMKfIXve45N3dS
USzptA4ITwiZQDMfTwW5PZentfNH4nXXGhtpOpJgTr5eevLgN6KNb20pVpc0kUyZekPcwuYEIl+2
cb1ZOWSDckEQCacypkNZhvjkdt3+wWCt1dpfAnxdtOyj2iRcfRTUTcB1J6ak5m7x0NlYhUzFsAM2
I8s1UsD57bgjKMPBSvbFN36h494C7MJn577m++tXaRlZz+pomN5tJiQUvpiTQnxfyYgA/dk9xvfN
seuAZIRREgE5Tkbs/33dJ6t1cdfD9l+246sZO2/EbpzKbUkxDUcZJwjO2+U+tG14nXKIIya4VOVP
a5S3XK3+3dNju6dy3PK0rGmQn+LBQtIF0JXoAMbo6SJkU27r6qCAUVLMVizabuOPRR/vGnHiFm4c
RrTtjYxUpBjOAn93jzKRt5N6FyRAUqiwCXRyxYCn5j/LL8M9iEaC93lP7pSvBgao/vD1LnQyd7jY
vM/lm56F768zLfAawLcPCsrCCT9zdtEJmC5BvuxZKS4VyxnxNSvKVo0PEercXfTak+CWkVEZC0AW
ddxAUflw4OvRQf7Rhvb3XcGgHg9pUXzyPUJTanp2YMYP373X/8BIefhdyIOST3EEMufKfPPY8hjU
fqSQv4+7ogFEyfOuaG01Ca48LkePV9P1xSgRTeyiJePL6mO0ZLPWxqeeVB9Ktzwn3A/kyzF+IXnQ
x5nLc3Se+8FR9j1V/Li+YPxuxB8y3LG3nRZIj7WS9KQBusi8ZvNxly1lslTesZvl31jgj5rq502y
zl4h3HTULh8f1tPBoaEBcvLuMAAusMo+1MK4yg5IOXvdhYrNEJbcasrneGIO5/5M8gFFpkwjo//O
Jbjo0SR5i4JSXKMta7tLUqKjftTQ6MEFDXmcPiPwhe02xfDEGnHrwBhTAHqoOMuC87Ilq94erM2l
Ntt/uaF+zHzKBvqON75uqM+MXFeDcdacxaktVbnTLArUY6JjbX2Fqcc8drWRKgJMQeNyndebr8SM
GSw8uxVjAxGGnBe8MZvlfrOe5WRuFbIX+hXbbT0cciQBZEu6yDGXXzaGYvd+Ut8trpP3DsyB910q
E+m52CSGIN/ONS1tZysr2eHDhYmfqZLc5OCflAfdsVmovTTq2LQEBNwJ+6HBrnfBuigpK3LH+mu7
WoEOl8nfFO9MMZluKTkr6NfkA3mfz2vXx9Tea4uGLV030hDsmvYCaquSfaA75aeetEuYWtLLqD48
AFzd2jOTtrGqVjZl+Cm2JDqW6+M6+g+laXAsrO7YIfPjSZmvMVf9DrOmQKC7UCxpRUwrU2ZlJG+U
uq16Crv0KdSeCnd6mWPySnwtJbeNg9ngFe2hRDhU5NNk6wBM1KcbrY+6RtWwgzMj4VVWgNDtN9tQ
K/FqMSQvBxM5sdbqLMkAlJ5inYi3ZQyGF+NwXKNXykdGzfj/zZeddlf3E0U6Aq+T2GLdtwHz1xxn
U8ap9tlBbvDiaLKRTaAGDKdwJzR6OTKFdYOk9lywdDx4odLJ2A/YcQJirUEQr/u9DJEuc3Ypz5P3
TUiKvW9O+xDjBp0l0bt7PfushzWALPamRV+dzDuZYlWGw/xkxqQM/i9007M8rNvmNVNlwU3nJCwN
ObWRYEZDEdkZhksoX2t8xGQTwdtnpcywqMjBDk759NGf2xlidWsgbycf24r5Bw/IKO0fkmOhY7YF
D6RshJVXTDyf47AE8uvC9NaGdOkHnVFMkIa8B0dfETdN8XwL6Ws/TFGl3BpSRF2yw1ZdywY8d2gH
kY9myLyqGMvGqIdacJreFZ+wVe1PTaz9IXt4ccMfJIeA14uC0c3duMcgBPj7NEuCJ4RzZBZPP7s7
zskjgt9tXOBD4JkqFUQru91jNL7GCIPtfWcBB13JNfDfX2GABgG39n3RtOHCYtWbamL+qVuNrwfr
BJHA53NlDyd8bg1e7JpaAwuKjVkRBPsDWIm1tAsKlmCieFWrO9nY+cG2x5xsqATLxGbRmIWjRRW+
THdlvv8UIgJK0L6nY0ljUGZnhtaC64+qPUEozFO4Dkpxw2+IM1CvnDMbI/RfChAIE6nJ7d2Biyib
yLuRKG2oiLUMVlzbBkKulQUcEw0SYgPxqnBXUdpIEp4ZGx0MyFuDFeqmAVKJVZw8GBw22fdNHPyw
nd1INZpTR4TPBc7ViUTgj2elswcKQRqxiPoxlpiVKtymowyv2b7JAztmGTOQqOCYn/4RCQwmzB+x
csRvB80Tsg2UUCIyYNz76z7UYfqILoL6iE78XrRI8tH7cbfvAuHzcgzaZZ3wOSEnToK9ybUO4HyQ
UVwSDgAPUhcaBP0YdF+KkaUFZYcowh87Bu41t1jEofRhM/Ann8ow9NfxCrEdJHMbdNOqqHRdyz36
0iOLGMzK5voRx3y4kvpvh6Sy19a68otCFJtMugwSTX202eDSdV8gtALPAIdNyOvAH9g1nxPOhmUA
o2vEMntvCFaZEIv1BH7sIgJZe94t8n2Su3n7nIcPs3twAtToNcunm/xupC8CLqEUCXbUOio1NID+
/UAfaKfP6AiRQSDctzn9wpcSU4ynZplspATQxhmxv0dKyD1laISe8W80adeyJ4BXreqr6uXOM9S1
7WMYtgVeJLTJfaLr8aSRrElTJULZc0ykvx8unViXqnw9DLDw5y55uKZ9MJjuN2CYxBcx1jVhidIq
Mix1mYMLUcrbroSdNMmC01H1yx20Ak5AQupSKIR4i750SFeOuPOxGGuVV2kIuctAN+sxYh3MF5ae
PyBG/2G1D0omrlPqd+Wm9Pj2yj1PjzpCfBWb001zcy7OBpkRE5W3Mhwmk3GqJSEdjTS1RW1ZmK8I
UdM9jE42+SJyzGx1+JXf4QLWIeLuK/AmxHac/YKgAeMthOhyrIQF24XVfsTCoz44RoHG9hYF8RVX
uGgPzbtnVlpa2uz/LWycp1rMLzw9/3XOdcBnbO6dSmtsF8WW5tMlSkrknZrCnaAfWzdL165K7oE1
5QtA1WHS72AWLJxBUnMYKIRRm7sDLQcgegKdtigFNHQtZfY+009vk6iZ6u+pCk7dkS61IUdo9J6o
DJ4mA0ID1/SCN5fcOdVWtYvs6b7RlJnN44zBb9woxtFbQGYt5p0Zzi68pqSY4iGBKoXMKF//5hWr
BSvZ5fxv9NksAUy9grlFZyOQQwAIH4sSF3MBWvamQjyCxt/JiIJ/wXmqvi4l06NklMYPvbGKxZI3
8xcsNrITYPGSKztWSYTmMa1JfsScA35csO6OEevjAq0KFv3p9D7KRu+HQXW1r8ZEiIVt1QdjVAJp
POLsu38Krn+X4B6aTaEtQi0tPApGVOcnC/gMXEG1HgUwN42pI82MSSMAzNcg1Koa04aDoWMJWtNu
JHCJoz33FTSmeBIutNNCmGUwkdMfW51lb/4czcDiGInzJ/GqG8Okjmj5tUcIjQVo9+UoLWhk58Uy
iL2OY7DFxQUu947MZ/upWAA78c+d/1mjPNC0lMbDOpmrKAET8gt3lgkLwKrWesYyTieRaYAOK+Yc
Qc03nmnBjMKqJMxLs4jbOkbydB4tcHqcjiaGuzmMkwCyqz4Bs4gGABNb/pqEgpD/fgv9OreHRjRf
urBDgXKYFqWBPpeZY4Sf0FW5bhAiUulAL1ik8BniBTSeA4xNhs+QFo1iWJ8efAr9ADNLFTEB+wPs
kZFiqZcN+13lvgC2LvR8rG6cKD7r/1cnTpeOkZ6CQ/n+MjkGlJjECv3Lsenzxx+hPfxXq2MwtLxD
Icq1tIVFabjBkV67aBcJZo71UKWBpqUBrn2yKzpY/4Eiyglbqs9MJsibBsTf4LcaTc/x+PsfOq1L
hd14MJgBRiTNhPGJPLL1022sTQY0h/hKUQ1ldVfMipQKYNcDshxodm21o2Hpa5SSFfxX27mtHJRE
cj1nC4axz8CSo0uGY6pLdo5kviYS+aKaquLgW32dAJ4Dgj4RONdThxrd2dxcivM1mvcXcI/Sz1u3
fxsXRsGYcUTm4EB4XJcagB+FRs10EIdjCM9XMuDYPIBd4GwZlbMDevveQCv9T4+SWs0CFvRfRKTx
PumlXzrFZjpdnmvC9c0DNobGhOG0sJrwdBUPYkiQmMBNAgcuAfaVHVt/zQ6cnPMpc6p7eJpcW9Ve
j/8MzYQOGHHcMxJ/mlVUhS/QXOFSmQOk7LpSqlqoSQSxuwu+A5copwUn7URKZvgjGBrgsr3xB53W
fzd5rnS626iXn9U9u1PDta5i0GoqVt0Pl7XafPZYbmSErq3dMBBxD9S76JDkFBYtXI4H5RzgOy2g
jgufp3ON8XwshxfwM4ZtG/23m+h+6OmRqAWA9nNYaCYZ5BBck1CXRAqa+oajEO8uHk7L2VEedPny
H6Tsu4tjlOWGlnIiK5iKLXi9fQTZXpNdKhgPxWsYBxUm+eQYPqqfiP/ai8G8w7sEVu+n7ABUQyCY
Py6aPm0EpsMfd1xdi8nQpjMPF6qmLYPsD7Lhve2rpzfsZmhEJnTq6Eh5XJYn4TgF8rZQjKPtZHi+
6Gnfe0m0LP4LsNH14eRxB+DlwitdRHRpd46L1G9moEuwLDy5IrA812K/SjqazOyw/jHARXnWFq1P
xNYvfUUco3C4R5OlI7t2naX2SCczfZ9+dVXnHY/GU3TLgZk1AefieVmdiFNXaWFMBKaiXONzUFV4
WOCy7dI5kKkT3FJDPKqVlO1+iz3hzow43Gkhy4zFEFGLlscO6NAywnqK6m+G+9+AgdSY3d4lHqWC
c1UOCxk4TV8OvDCxuFgLkDtjKtfI3Pfl7CekhLMfHipVKBpzTaER8fyM1D9tL007FhP2qZD1YCn6
tbtcb7Bg0zhopOnzW2pvtw+2cFa9S3gxsUHcyIJhsdMrGaNJehiKXW2Rf6nRJF/yZYkmguC6dpNC
DdbhsRwerVRDdGxFZRxqDOA5lP8zT//RGC8Nn/gejJf7n4xl4vFpLPuKLDR7PKWbNPb6nEiEhDUc
EPKx7MMEFw4BP2tncLLkQ3Bdh8W5jFCXA0lra8lABmLbjjk3yqhnpzTy6wo0aSf6BvKq1sEYnk7u
7Gu/B8FbJ28dLm1cGu5LXbxK1iN+EPHdDerFCf/bTAbp9QVr8qMtfBRXbCAFU36Y3/4ZpLVQCR6C
GPU3NfuG26y6rg+WKkwF45cKgUlcw5aAXBKZANmpM4AKlv4+L7IjkKo1UUcWgKn/nLJC4evj53bo
Rw8+eX3E1Y6oAnQw0Jyphg/lu7aPRgi7F8yvTm53kwBQYN7UwDWl+mRioX4H7IzpHfWhfmFB5nOt
MmJSexlZ7QJqteB1CpgQbxF5hZUQ8KKufHpTbuYl/7rV42z3F6bpaEKvuruRzwS+HW6bzkXvt+3J
vs0/OLo64YWFZBz01CfdRJe5WxSqzhUbIVUzbdBbOYRl7jdhO/ZrkKws2tMRdlPgtd6SOoqdxx6p
SvPbgIR8ziXOKYm66R/djtXjsXikl+ilfNo3XCrWvUXvlAWkjWwXnfoEDNmgmFV8ovyb8MgHxXQ7
6mZ0QejJKXC5ttxEpaCHIGNMehP3FRe4AgfVWK9+lFO3FS30bcWodqRzMuARmy9ot1a1FJS3iKUq
nQdg3N4UP0tyJyybhW9CaZF619P79MwaSLMgz56leE4tsBqsy4AqCEL+t4Hmu064yHZH4q4GpJlx
Os/rM5TO8ZR1CefKdbxIKaJKTbnmn8PszUAZx21P3O8gRtr3AicK4XFmc45W1st97Wa+pRl3lJE7
nxyTrKrkmeH5ar4IcEgxpOF7v8CzF0Dg17gR6ICQCS/BAvZeOlduxPOmYMc6iGt9/WZljbEa5HPd
J6Sg3kUrOWIdpHMTFKWLrGVGi9ipW0lcKgkukQw2EuYkzcQIUSB8wLDpLnMTVVWd5/frkRL5UVBj
r1XCwzzEWbr9KFsOfhTq4o/ijSPlCnQUpU/nFR7c7szWbX4Xau2M+tubkdMw8GCt6w55Ev5enVzW
1sxQN5aF+3fotF/zFKN1FIpwGK7iL1GZTY+/xB1USLxnRDO8awMWR0XPM3Cx9eSKQ2bHQ7dhFiuV
uG2e4qlGD7GHApgZ7AYuGbeNAnQizUTVCcu+WKu71P1+KK/Qe4cAED/db3nSS4DiTDntAfvn9bi4
seRehg/+iPZApi+GIIRFJLixK0SRBAxWRROJ3TNY3HUpdkBIqFCUDLhWcHndEYVGmI3Iy6m/3JKD
gxM57HfX4o4VVCEWwUzBM2NFNJPB7FEfy7w7znr0t8omQ+v61mzJltJ0bokD81TqDR+Xse4aaTeT
bY0YZRJROc0Hk2u9xtu7ORg8ZsAVlEY+RyscIj1ktO0YTT9stbk1ccxuuizRjqtyAHS4fwUzf7dR
DY3pUjQfzFTb/vne6zdn6yON6rDIgAK9diKkpc5pufMk3xl8rlLMjHAYx/BU5m0ytBhig13EkL/v
WF+fAz6gXg9+KraZ3zgWmiZk/KtqHjBt+r2ZfV/qeC+1MRVUk9BY6wOSuo22RqbAiEhTNK7yA58d
uTd8YUu+4aEVe8IwuWDEwheysqicJQxy/6k1K4DmM8LS26TZrpmfKmZiHeQRpIyswJNsmw1JqJo0
hhXmgusA/1k4FHGm3omQIHZJPehikHnRw+Qb0dTRtuu5d2QncvgzEGTVRIUitYyD7C1vMJQZFPVy
eBswlA8IesLO93QM/7soWKzA6u/+wR1nqG0arYVsE0FpLUAzxyMhTmkS3NnrDAZIPMh5Db2W3uZ5
PKfan06qbm1BdHqG/DlzghKNMJw2cdWNj0upsyPPVWbvC9UtnJCG5rC93yiGhkKB1JDsK6BN69c4
agm2s8eAf6sapVaAYIFGGy0G6ErGXp5qgn96oKdpnWfGL+KfM8nBkg/svWAIElUtAp5WfUgcxrXk
ikrW23gq/YcwrAjRV0VpnCsq7knAVMsc50gDyOvZpjwlRvaWD6dnT1pojaH+Svp3iBfxdjB/KNPZ
+s8hF+qnX76NnUQhsMr0sKUM9N+xUkXJnJkWCjzzlblnExCG0Yp8S/fZfryCAlkS6RzQMTM2/+qK
gY5LXu4jAETzp6USAzm21oNCYTjdXKqXtLmrPft2InFagFjT/vaXDZh1ugpZsmgrxsEaiPOjLYci
SBXPtpAODtZsa0eexQURbhbeom1Hlg246tFNbUHDIqPLG7HPFgZVnX6NDIKV6PMb2gbQJF7OKo/U
7x3vZD9s2XNZ35eAPKF5SARTqjosscB01vwM2hpQtKHiaEj+4KQahX6s1ymWC/NxbEifGyGemq/7
Fz4pliiEdMl4mzgylsPdSNHXl2MZl717NBqdZu/v9ouQtuRzarlzP4jdzmeDHqm71rVbYcGI1LIy
fyfOrCpYwDqK/Y6kee+BZw6c+S1C757SualK8LHH/4Tulc17U4MHpM1vNBBMw4mrgoK+hVTpJK3n
EygJoBlepjX7hk2Rc1ggC1SF9y2C7CoMC850UrGkWYOcmj54ujRrpsodPXv23oAJEHBK0bq6KlG8
b4FM2aS9BrV7MnOAFR79wTvkcE1NmxQg2N+O3yshFvGHxFmq9NyBx2rMSkvT1wAhHr/CRhEOTuWQ
OknKRuArZ4aFdJu9TvB6Tdhgnjtd++n2aJ9+2c0SQrxO++xJm7etBOYEw+R6+V/PE6k3/6YFpEvc
F5XJVMGYKam+j/kG36uI9s0OmeNiZg0RwF1GEXJz/u13Y9bqSGbFWEp9Ee503BjX2Hi1fA/5UukR
X9pqJqw60EcQUI9regacv3QxfKokefCFzsT+cnUnBM428/2Ge6cyfkD/3xiQWJJTjXwIz+/EL5jG
/Rh//FnGuAVlcGwEfRTiyjPOtUvB0geHkRm799/JDlPCwwr/MFpFkQeNY8dGCaRbLq44bWA0vTNH
fFpx314CLmForZsjzwdLSh4COjEme2j4q4PB+pE9TOqoiF9IugB7xzwejpikW8AeXR1ybCSlygW3
ApbyZOfS++GKy0DJXI6YyuFLuhIqInoqfIGNVjxM8gMruBq0+1Ht6I49wo0l7RJHRHtHgp5ifGMK
eAJbxe9ETKujNzJQpMUQiPaFEox24w0a+Cm3zGkl61QZASTFnsVyWqZ+rGT89YfZOhFz94TDVsTx
NTlR+voddSlnNHvXEf6GRvqkFfO5FrLBB9pRphtz3SezfOlmc/Jm/2FJP6u5jCHS0vVrR+86z7yT
+wJf5MFH08uekUI7Ta7bwtqG/TMKG0rd49YK6ZDfX+t1F7Ie9+U6TbDCuBp25e1Bo1XMR8MChLRR
pk6jcenOp9vRnVSE3SbXlwOPGaZCEx2MTV9Qz4DAJ3XcTTjufYK73DYUjhMHKI41ty8clH5il8p0
RW8GN1ajNOxbWw+MX+jSpuGk2OMLzQLY8OamJop8tFy/smoa1i2Iwuj97nOP3czENHk3l8Z9vQRX
qJ7syU5rXMu/TJfkpDoZdhIjaO7R2aE1WjErp2gyPTEKP1XI8RC5u3vPSbwDpZlljqbpSwX+8kpF
3STFPxY7Tr2Zk8WbChNGyqnOg599Nkn8ZqIV88V0SPrbUp9pf9vaFUsS5Jkq5qGzHgwYhyTyXpmc
OiGHwfwl5Zt5TXFb0Zh4Lgh0leWylTGZLSD+mKCKI/vj8kndOzEI5QO4w0U++PrVDMca0vpVN6S/
bT0LQkafBwLxBXOidI0t/o8cqIyMBJYXHbalP+8/M4IYNDirfkgOnjrHBnGdkNaJG+i19C3JddlS
YRJjIa0kbgwI9z/1pxBjS6tpkq6bSMTIQnkRi5yCNh1aWrq0TvK5XHTjdVqs2HIVIQnDdYL1EowU
drf43g4Iz0JQ3hL0miohUnsfwbDqRTT9KmcsgfINjG2L31BzATz6cVlWlaPPcRxLuzyLhShUyuQz
dTYMS5rD4rZxWSXT9lFT6htlnjDol+ivla22h2qSTgOG5keaARjl8BPWGhht1WV9IgH/N3NDNxdz
wtcRrARPnD7SC3wRZOWxHMsc51RyulfwfpMpOtgahA+YRcE6j0wyO1R04VtIChwBypf8yuqMKx5I
Bv83qdJgsU5xNLNqvq26CDgEYbkXfoIFHsbQfnKmzTUP2/XRouk/C3nFhpjpJWNZ0ylG44hWjfAy
bOHNv4w7IVfhKb29c+3qQTtEUQ4DsGOzFkD97b+tLZRC/VDPcicK/DUjrnzDaQAs3OBSh9K4kdVG
V42G45Eek+rUHasIYFOOzGgws3qiGl2Gc0R50P2YG1Ft3MdotdwWw0VLuBm4u0w9VGZoZA0JxvaE
p8JzW7IHpMoFpyeQdFDQrJSC+vrS/yB27KpFtdcIztUSZoooGRZM3UyT2EdXi0Qc60YC6ldJZusC
Wq5DEvrm9hywKAyQmZO4BIX20AzqKDOtJRqlAhZdi7nOfOUkB4MvxeHfJjcvbfeyBXtCauCb23MI
ReoKQNA3gCAZ7AHthYyLkOQl4kTuUottz1HgHVp5D4iE2KfDcHKKZRfF9C8PNRnuwCvGr+TVfczM
b9Q5x3bxL4AsqQFtv1/Yj++/t9RTmFQbgsgmNS4wS/eF74yRXsToXY1GWEWraukxDH/aAtr2yG8f
GMxwJqKivYmO4CmeQYLqHKpaTxqExyn1uTShqFa469Ax9JjZkhstrb81U949COPomYqzgdF6di0a
6Zfk86t3fHUF2NkGAv1wDvRhGj+MdtXgccwCQ6ag6tja0H2H89gBoskgX/SpVpomKIZWMUUKKwR3
uZeYNUmp+lMSHq7UPZAblKrUnie+WHD2nd33o0WkRmeVbxkbQ0RlaF0Rczbe+lIWWx7/r09MX9yn
98OosYYWAizDbUQk34FXcCSx+IwKS2qhowfDQtY2Ysnk5LCEimBqI8sgB5eZRyOsq0aUeGxoKJ6S
GgTDiOTVKVUerodfyvW7sOB4qhCFKR9mDVbarFPuJ8YrlckUTim6KhfIMwbWnbjJlaYZuDFk/KY7
r0KW428Kz6obJRnlNyFPUaIG1z2g+JuTkBr1VeXBC2mxdK6vk7A3dM5olNt3L4tYMSsGchyji9A+
/C4XqtTXtH/WPyxqOP1xPm8hrsv7YocwrrM0WqdaLbYyDYm+HMaS9FcQ59kNc3VjV7IXWrONvGPS
wPBXheV99NHPP1is4ing0Ux2OqK54MIonEh6CtmdCxCCTLhf3MpeUrBvzCJzenI/NKtHUe0JbyPZ
V1W0WLqqvzVcwfejsZbJ6tLEL1sRh8c8/hI+4tmsjX5bIJGzWkzdKZuHE48yD2gWc5h3BCg2NvOZ
uj5foODmHUVj8qhN00KbanVo1krKX5uBkKfK6TiGAkdQZ9v63Mx76Hj2FaLDh6RYp3cvGsS1ODW8
ZRyw4buqnGVCZCS+Q66IE+sJYiRoJN3TpKq9eEETa9lX+W9lO+zyhBKUfCg5KrxvlKnzPYT4eXxK
EIu0i3WeH7nq5jmOrIWYySjMleUZTXpdyp1XDQzPyb9f5k/3IOvVOdrFC8Rw/VrwVAJGFZ37MGxO
y7gvzJ/NlOV5J0agn/1CpK0bs7fMT9QjuQooslW9PHoIMLa5/CgNSpsa/CEO3W2/fusk73g3lYb9
K68HC1hyIGlMrZIcTUJMeM/49LWZzFpHuzcpfffFkVeaDNdv+ldAVdYy5qIC4+j982a46qho1U+x
Ro4OGSvA+XoNkLEzoLJjCUAjma4hcABkOgJOg2hANGB+qwD/Opa6n37P6Yaq3swAE9yhAWBvGODu
uhvA3eutgsDUQiYVbARg0ePSeTha9rtSRGHJbZAnuGGm9vSaUs9n3x84+DZXr/QybjVRaSGhYWOr
P9KyrOENkVgsP5qRWvIOEnr80vVvXMTgKx3gDDfRwn8Mfd4BFEyBYWOjE4rqzTUzd7+jJeS/Ds0u
unKx4Cf0u06TDjCnXd32MCFkaN64iJFTfAg4x3NmPwbK+PyfkB2ITcdGchtsXunRPXhkL+2wZ8hX
zEJu37GCRdqcdCGxBRsU1JIiPTeAUfbruVCO5une6UZ3sUGuR4LsQuqmJx++u2HNCZwIbPRf4Tp1
nUPfCtPDTVCIlu+nmyRTnC7KcJzdLcVvk/Uu6VXejkuaetEkA5CRt3XtgtnFsjrncsp+hjM6F85K
Qa+l2ARW2JNX9Kc1mlC/swVxUsViCXXp46876SHGEr2TGr07BMfE4wvU170Xp6KxyaZPPUag8VGX
Khf2C9S6PWDqxAjuy14rwNzPftg+u9SyeGJE4aGJcek5YU+AjqlwqCue4TmogjJfN9l957HK8sx0
ZYUxMXQj9zKbmrNmmhyjjJMV4OkwIkohc2Maq40ueMGO7fSQyASHY9Ln3DgATmbFqOih6gPzJp9F
CEF/k15g0h2QWkP8uta2+oeZQJmawILQn97N+gPL7evu8awjDHYQgELwsX7l4j1amWk01AF12FVX
PuYl7gKxEiApN8EsDB3aISGE3JW3rLEzOqx3o8g78AQeox1wT/oNkVXgEULQlJSi/moATRG0+c3m
dBT/xi5D3n/LudLAzErV+Xl3qvx6IdD1gXuDfWRXPqfAJo5N2YQqs1vb0bNtlI3kbKr1BqSWwNCE
LTOBDlNIF3Hl93Ek0xUhT7fySCq/MfyOB1rNIgZFQ+XPNIRlKxcgg+gBR2kMEFbWov8qSoXC12ai
PtMz4VviqImnU893EgVdO7TcoNodATbTxLhbc4/rBxTVSKP+ywjKCp++Ea6Mjhvo1aSDM+tOkEWH
TubAgZy1ZAi58W9jMm/Pumfd6Ey096niSIqMrFuXfj646CMy9625SnIJrDyVCc6XZcqg+evHMFz+
ceU+cjPmA1GWTKEqAYyghFGeSATaQ6yfHdvqj+y2b2z6ZjNcPoQhvFIA/MBIKGMEDqVquvEWExI8
Tf1G1RNqB3mHkKyzmAn/ur8N7g8krtPoF6Ky/k6Q4cZxCL1wafODxVnZhSlLpjRWatiphBLBER73
72HJK4rEm04nQ6QYNNckiGLk5Y/r7gdi1KEIoZv2zagFNxXJ8yEH3ZomfiDenBX2tvNbMqrJaL7X
aQGCpNy4jksdy7NXr8B11UfsHidsXnrFSs52WBwEDyfY9UolnfzCKUcpfn0OeIpiRBNlSmO0XdaW
BlFrSMyV/j6Na/4uZlMebt/Br4Q1QrPuW742Irh80c7gqVPrrPAglA4p0TZcIC+Hzoq4MJNOrkSU
JcvTT+Xr+T18tNEMMyKCM7/7aPjuNKpa/NWWYQjCXNx0M/6zNx2UjzOyPBeluuM39XVgoAUQltic
lv9Fs166K032vNV+Kd1+9N1zAgqxXAz7gtPa35mimXC9y8d+eq8vWdbGgwmK1F9dxEx7qArYkPJy
GUsQDzUv0yjlENJiL0UArOGxqETi6gk022lF+R34/mW5U8745JjKKfp8v/xa70ZDFlqgfnEOnkPO
VmmxdMs3JgZQ+Itp0i2OxuA/R2Hw8khQF3Lo3ZrkraG+8bqT24QBLikXw/OdaXEAE6KIJKY6I59A
XstRaXZfLOK2j4jaKPrdLkBnmL8+Uqquic8Pt1dZNhryAU4CZjYlhCYjP0hCmjHKRUPFRI/6mQPN
WdAb46CzcEOW+nb1zBRnV/mP14PlDM0DQyW6mQblRxKZXGizLCt0Ozc+gOsCHo1UW7uflMrLL2uw
I+hHbdNmOEowkNKUPC+MVuQ6WTYQVhdjDLHnvYXlKT9j82MffLwyzD/qKQFSJb3By9JAwARS/C1K
wjps8IKvFv5ZJvWLhWGJQtlEyBT2fbBFU9LgbnyDs5sevUlYs1BJvHufuvrClznQiq36gqOazBr1
dJuYNM+kuf3mU3rcwql3NqzUea3W+wtN8QFlrsQHX76DgXuzO0+1PFMwtKqQ10Sks++20pqFzM4K
z8586Vm/0a+Fa+nX6jIGyUeup6258CGYAr46BOlPBo+DpWk9sHOSMjUkYIc2p4tIyEzimkaMLta5
HAMk3glThGwESXw1FzPV16BPIfzEw47uICXKnI3hk6e7Ij743QxFpG/ox5oWClFhKqJ278VHPJwD
tCqnEqSPEPFar8DmON3IxwJdgEtp0NlnxYQmdAy37HKnUN9MnAPuqzpnabfGFND0dpu+bRtN7o6t
dI/SlClOMxsDQIcroyIBauHK8kv1+uO6HCa01bKRfVv8GNoa6QKrGs9QzKfY4Be6tBhUArdMOPs/
lfJ37SETUZFOhHGLQd5gOkfSNqDttq7IChAwxnkc6r/5KP24o1wvft9vo2Iw5hOq2hp2kCM/yfuI
uXF4pRBFdsUxc9tn10jPMaITEnkib5J2vRGHA/C+ogBJxpfvvlkqxg2sgRE0rDvfUM54MrX2Yq5J
4KUts5IWCa7jVTlu15YpPNBq4pRkfY25NsrnWfKVgj+I8/tNOUSMYKBdimuW38ILRK/QarqcFFPs
xXUwo01FrQaD5PLiVJmeBv7wtyjme8WRjdU7ByvQk0APhkIeiKs8yKMJM/AUsrDykkBYWdJJ3HVI
QmSG98wpo4Ycrqy31zmvBzVKC3PCdEg3N71LvyTPptYO3k1j67ZI6XQIyjLJh92EE27Qlt5nBtT4
Aak7uDnk76gFKVhyvuN9C1XgBL+yBEQJiYeUvq/ip6IzXpQC9P2//bj0WEn971cwbU+KqL678gjW
N0WSIMYwKYbm1ql9cZENZ8V7LJq6sbfOR6LX+DEDvOhEABKFHDpWyaA4YbDeMvlnZAnUQR2Bc+Z4
6GB67bbxpUaP+SNjZ8PDTOx9lXNf//EGnG1bz0J9wtwdz6OI2Xf8TUhppk3BvW9CfdUdQ0mGKxyo
JVWO+Jm9Au0yaMqReITC2oxLFwX00HXH6vhLnGxQabylrv2e/w/7pcICMLXZJtBp19qF4GsMlVeu
yKIflI/OJL+FaHnZdHK8Y1KTsGXkV6cdHxbMHaMsKafDgG0bCCeTmcirFpq3IcqDY0slkYwIr8Oi
EDHk8nygRi4qSNa6P1E0nWEpyIWDq1+jQXezLd1CmLuJKZ5e9x8O9B/jnSo1yeAWKCCXwH7NfECn
PCjpbeTw+HwBWR0VN0+vx6llbVJQqvWdHS/D9S4zohSzAF7HMH/Titf4ruEmL6Nz5nkByyLIrb9l
BLWHThK5u/JY0qWYamEDvXS52AniEOyXu82NcHyte2qD0yNKrIvrsC8i5KEYfWn+Im/JusIwpewz
j+wNcADxBbJdHZCCK02SGfHlt5Pe7ADiyOFDMQ8z0eQ3AD6qSlb8bN7oKYjG8bcDxvzgZsvJvaJs
C3GcDpmT4uDmus1wqhyoat4UZv/Ez9Rbel7dD6MDBmInPdypV8XYD3HSXJvrYXmdR4XWsaiLfhkz
Nt/r4p34NUZmRl1DvCBboqz/uPZALjXieLGWG+z6CpjQF1gVqFeR/ow+bopRkADPMYNhe0hV5Etb
ItlAEqVQQbtoqnWIzE7UWSLdZn/PUUbrELr3yqDo+csovnL36P8jTYxdh9Pizc3HpAgsi6k5TNKo
WS4qKqKDFsa3pfJ66mUo7xddHdsaYfelGu3xLma5RLgLu+MQbMcT0PPYEUuZtO+C1xuTNBEhlLvv
H2X940jOR/gkG0ECiIiE9uxUZpLp34HMAfq62ERwqmPakLetc1klOnjR1EQQlhFZjiWxCfyQrGj9
SgiojiY4zp1a2RhhTX6UnU14FHhBpsSZ6Nq3FFIajuGppSyHIHLUGHwdDpaKcK8HdGae0SInjJ/c
Q3aaYzbFzYZ9wsGDbvNPN82vPYnTYjGqQBTm0aT0X6vUfrYoSKWp+oXdCd50VqOcQ5XN0OMrin81
W+e7XVPo6BWc00J7u5ZFtkuUDRFXfpgNQUm0ZB8bast+hM9aI+Cru0XMZvTYNszYuZp0LZNM4Ysf
MVK7VV0xXbV/GmJsAMZSSXCACmF524vP5a4Eex/YKRxPJ2IPT97rsU4NfYOrMVUiOkhP9u63LDup
iw4dh1w17+KzM6Cvyaec+eAg3MMyuUW5nmRiE2ypbTHU+8NAcrDAOD4kTu1Rykd9ENdqesJ+i7DZ
LoH+5ZYrYZ1fmZvJJdu2VkqCBJcCGh0QYwmIY60eIP8B+EfYtALsE96EICVxtCbI+zWY0645dZci
EXBlo0oc1ldfDmjhxVOBKTjK6Go6N0N7Kldf1srXZJ4iH9aq4rdlNgM/CStepmci/VOnM7Mu4Rsc
K9MPQundGoddN4iIaoa+UZBvhrg9dhwUN+27t1Dfpr1WKaIlFgYGZGpIFJm21mmFmZSiHwuleQzu
eZdDSYLFU7N5j0CwYJBZxkNebZpKO5ALZKSzJOvAFqQBiC9GujbPGtlKG+MQENbNdKpvLpzgvLg5
1UJqgXFsfNt0IQ3EhUuXwaSGB0NhmSOmQ2dXcoGLp5Bq9hYo/XdX24975KqC8STrlmRmwhGpvBt3
ZJA/aFg+byDhaea1feeACFlgantOSs0ddk4ti8BhfOfNMk5RbWR2jn1Dbv6DIxWoMaotf0rxFzN7
WD2znHLYsl8shobqN8ly49WaZS8KJlLXwr2BoMgehT+Bhyj3/ZwDwSS8DlJgYYWHduDNvh1j2LQe
SbUHWHQ4gNVvZH4xYDlNB4qYhqUd9zQ8QBW5XtGJ5ipbppafJWDd/JF2bfSrcT6805lQVqPFpkpx
qFRfs0zPu0b4JoHvfNZjBxh92HCqk3r/yUK9K+uQp3odnwkDh6QrERVkdk+EHrR7R2BO6AqC7JiO
Bgr5bKBDYj7BrlSTzYXenr3ziBJlhuAM7iNbOWnji37bbbQhbQlNCMNVE7CNT6sJXxM3PxlsZRwF
VUW6gqQkg1c7xV11hjN1S0cYbsltB3BeGV/4SH4ADaMpSKPeeM60Byi8pu5tXR33dDRM9Z6oqRBm
X9wDesoF1QstCA/kJsCJWm1pN+HTb5JyK+yzUMH5TTPmyN8yfeKKMRF31jav18ILGw+Ge3bwSLuS
DXGV7hDsTiA1J2ppw5nDEVl855bsy/3ik/wKQ/pVOhCotJlwGz0pRLtmL2GMjcif+5QDw7vQnod1
NMwoMg3E5/V/+BcGkdDfenZgzH/H32dStwb793pEh55zjGHy5IGHuHy660oq8Vk/vg+zzbRu4KiS
ZKne6DwIwzMMQK8BuhITNUKdhvS0s7mMIO7D/BqlZipFxL3imPt6JGSJ6gEwgHnm4xAiDRZEt2dj
0+IRdcSen89q7Bvp+x+2hV/dXvqm6gGwSoKrQHbLtaxZC5yXAp16UCwDYbV71kd51xuwmvHtvaIx
6H0W3iUig+AyqGebkZ4SC0eQJ/pj1x7CO4HAG2ne7p9YB53znKzdQwhEkX45K1z+N02jeM8iXZp0
M7/MMDeMpOZ/T55RGpNeBYDxJGjoHB0swPaBJb6AL9GK8nZw6S0/khYDij4P3imlj6SmzzN/23uS
LzEkxXvzn9x88i2qsXxFP5v4q0R5d3/eMb5Q212Y/QnORDPXmKnjVPw7kgCBTGizqqCaGofPAZyS
qzYItNhyx83Lhuwnjxrbz+X/y20Tn5sWGY9fZvnIrGyCA9f647WLENap+JDEszZJrMYIH92WLfE9
rlCo8a5b1IUbd20ZL7oIWPzwKWjFMAg3SZzxTqSxDg5zPgrArttQRtXSH/DlyRW7O7dA5jp6iwbo
osEyOb5BJzVvDOhkHpNBq2bMnYD6H6Hyh+v7XcUg5d7lqUg9qkJQEUDz1btNleVf745uxgLelnAK
3KkGuKqfs7QzxuqIHHREFiDXvUtSWgkZqkDv1nwoN/wFD/JOUUzncxfpMuwC8Wry8PAuA6YnkE+Q
WPO62eQ+B2gtCSUL6VEjP7LOU1OjpLpexg21MBLbkWl16h5mLyDl3b9vA2I7OKTFrpSIxeYAU0rW
3UfDJFJp4/Jv9sK3Sy7ZE4UZqynTBur4x6CDH+/Yflu6v/T+geBJrhZaiELtOUh6Ese6E5LGF8oU
iE2hcyRZTrCvLDjviOAx53amvdH6zS+/s7dDYWqTdke7ppl/5Cdq2GQLr1kmK0Wl+ovQR3WXWy0a
44U/uLBbUIQET5xe3jVDrK3r4kJhEoX5qDdgB3Kgnp1OGrZmvVPGzezG+88DH1ZQ2JiT6psT7jkh
dhfPvg2/gwEMSzz13Ul9AORSV5a+ppM4KCJI1eiSwUCzJ2vRof42ymE5l1crpyQ0TWWsSJGhjHUc
G5gbGU+kv6wgZsyhiHQAvxAszWMtKRE9Jl6O9n37FIrDo3dr57p7hS6A6HkEo7XDXJnCmjD+gbIy
BVwJfEAS4zHuXZVamAL/nehrto7enqYkjMt4chXsTD2ur+KADtuiF7FxgaTCQ3H6n0zw+yzMsoiK
3Vo3YN8bw+mDHiKEH0aUOI7dI1M8VjFO1LBPHqHJV+DKbmDmDISLGTmitIu+KvYOuVte2rctnggw
8GcFOaI=
`protect end_protected
