`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BzuthAdvDfdl0CCII/61pOeCXEfAmiupSv76BNYf+PWzobdufoomH8RelIunxtMCiFzOICRuNZuc
N412B+mB3Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PCdWclX+uYbZBFUDCLEPUu46oVtWJVHPtZmBwbf9UqAdVoddWYMCr6mbN9WePG/UTj7jutr61WHG
JswyX2MMzGO2XK/FB1JHrBc/DNPEjgLO+MagihzDULC7T2BhyVjtFVoQdoTy+liSDYdbyPV+IJcV
Xw2AjxEeepkPGhCFbLY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Hbi8nlq8tOlmmsjmL0/mmwiLaCRJLOHW/B+TYpo+WM8AdPCxCZ0gjPITfuysAWxNnGEQAsVBek2p
XLypOkVe/CNAU/76lNsK+jSsYu2eSxez6J5yVNU22O6FlSNlYQAn/LzABXBwlloxMGZU4KS2sFlX
sxZi/fyaBuDfIh2SzwMrQaG2e9cNSS4a9mui9XB+mfgGxC9L7IgSDf1znr+L64hzOWdzeh9+a2MW
7fet60JIUlE4zPH4S1MRKB2WQKxWGFBOeYmpYphAXbHQlC0WneOo8p79hkXeZAcc/q7QcXlE+dgD
oQz/NCidJvgVcWMQ8ZU0+7Pk58GYgkX3/hI3MA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
v4rKGni41hGtCcrqBHzUnhnhlHoyneZpm2LARA9S8WbFbYw71jLKketgUnRYRQjgDESn6bWmKgjV
wUZ5wDJ8WqqjWYpRd5cKNN4DSBzOvMAp3pRw/NFtAj6ZBYakAYBS7WADERIofrw4QstdTOoerMFQ
4G/cmlHllgpOCjKLFT4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZS/WpN2gAWLRgBZeVIapoSrAbYdLnzm+M9hZz3e9S7jsqdjHu3KDnjbSQIiGv4HMtMJt3oHAWb8c
4r4QfsovlQ9SmsIaCdIq8TnJN9fWMjHWZinhcW5ebhE13aJYHK5l7GX1faaXMRhFsLJf0u7Ladvz
Oq2r2HXn6d/56HqtFTiutRDoSh3bY+OF/mkbfFqQ91C98cM7mm0TLixidwqRDDOJbJVRQ/fljrXO
+ZwMA0s0gPpEYti2M2hkSLPMMydjlXBl8mYzMf024RcIysi9NhGbUHr1MkMyuJ7dpZpimN1DNH+M
KoO7JwDf/4OlAcwIDsVK9QT3OiCXEvCG+yChvQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54512)
`protect data_block
9T+ZB7gGAF0l/S1Fbw1xPe37pvvfE2Z5k3BpvXeEWvcZozM1kvDiS734gjYciTQPuAwcbJNICSOE
wdsSdLxKp9Crr4zqe1+9JLRjnmxOlSQpEfziZEMrsLXpngywuJcmS5ln9yTzBml45vr+xKiwIdS/
CK6HkX62HS8PPd8Bjp9bKiKEmDep9Q+i0f8STErB/u67BaY8x552tL2+1IdAhYdJKAPZS7nTaVAb
7xTuL7t6nhZLR6DBUMsqWu75v5JVOTc4vPPikRSMpNiL5l8cUeMkqOy7nWea4/XUjd7n5IT/6oOl
FUWt1LjtYztGMyFLHscuYWBycSwlYReAzEBc67yMOxU45y8eY/knzsJpA3p7pNAyX8Nr1HQtOUZT
hLUbzJmow3XpIV+oVY0q9SRwh0sb2Wpnd+fT9Ugvl8RnM74dVXRfNBTKTEQVNT9tGWaK0JvYqDWq
GvRdcD7LOBJZLdMtdHZhW+Fby4qDXM9Be6kGrMD8oSaZeK+NgeWEszTXLoiO66NKe8xFVkiV+LZh
/OGaDyLwq/ZDT/Yh9xsvRXIRnGruyqtw8kqsiQ8cHyNvi509pER64mTgrFMV7tp/fyk82IHhIQAL
8NSIxaCnq7V2bGzUUmblG0z72hy5TZBjtKYKOpHjSjgt8cG7eXawRfKHkY6BlPKDhqAJ4u9E9IAP
edlumy5/3UzbaWdcyFpYbWdGFNtC7AaKW0m7fYl/1bkh18K7XZu6rM9Zcs/B2TYV1xafmuUmdfA2
9dZxzmV7gjOj+jzZc+RaylxNzbrHQNqoU6NuxlYkr+izXptupux0FDTd1Isjx+r83LM/iWFtuNVJ
Joa404f3XtXkPYDI2Mt/awtSTCRQ7P/EMdYvVPUOFziH0hlsyvMPS11TdBrMyH9Ch6NdBXQVHf7g
3bbesktS/68LRCAj2gV8/p3Lq28+sf8YU3XFdGwYkbjaI2G5c5KDXIz/hreLOgXM4h9ChDlVfD5v
xxqnenrh0WcKzQmpV32kmscQWs3Bc7m5AWpxv7fcvhYPv14fcc5jke9bicqkT72iIGn/xZ2VXMEs
6i8PPjX06/5Aul096QEtHUeaGLcIHuSzBReqKthqOp23r7DrcMIebf42ECeWf3KupcdDqSIeoI7n
32hXLQeVsYFPB5fbUAGIKBhxQN2J7hZ0b66VN9qOtZnxb8M+tod9ab65MCYqyhpKyQABzJYbKyHh
tqpfaC7NrgOih8fhXeWeB/aBKoZNkNS7VioEd/tNI39gW+jPxiTcqfLUxiVI31HhOERqWDlq7cmC
BHFIJMWRgDSrCew2DE8YZQRtSeA0EnlkKDTNp2AY3L3+xzxzWGgaOxZlVE450IMuXACu4WkMmotC
+FiQ+FMLkVpBhqdB5U9KEeOFpNwvjESFtlVgv6RSP7svbWS+TgN2HypdS9wbYe19jE5265U3hPt7
egV0yx2ZEuEUM6uA4LhVGkPTLELHzas4Lc+xqn1TA5DV2OF/2O5OleuIhPQ8h8hGxvV6bIoiPVec
enEO88PdJunlHXfysFc3BSu09lNqXXwO99h4AibU9Ui9aTLc7Jyy7UHKj6XIlx8oEXgPEY4BdULQ
qYTosZPsWznttC7FgPRnW7RwkR40B9oP65ajL3LYC4u44FWwTcldjt+VZh6c1w8gn9pSpIb7X0q5
FFNkI1rBY98XiVj6GiYB+2nDP3NVsx7oFOqYsNHqHUH10hv5oi7EF0J/20qh/T6eknWrMQB5XYR3
VVq8lXy35AHZGFxDo3A2uLcQVccblTuS69B4Hc/qn2lFNXjepQ/aoXG0fQurClUKZjPB10cwAN4D
a89Nym4xU8oslv0Esd1m0iZIywbSPp7HF0R38tcoxL+wQ7D1mJOCMnIDMvRkBGbO//0Kysktw9OD
AfxfH5FC/E+fL03O88TNml6gWD6UbhqOnvfb3nl3QHAz3mSknayBJGgkeM4NrGR2BFWscfBhk+u5
n+wEnKr5BQeMBEztCBUa8/x3kv/Mg9/vmm5YweuFLDnL7yOdAPZy9SbFLY0k/sH6oIB5Grutfmdb
LjLwZgsCgnlYWbdDZ7YMVkyrnwEguiBEuEvJUFl4fWbKrtLzqohtWAcn+NzoElAXDydZGeYQ81DG
tlCf4rT1z0iQkieO3cZzLZog2A7IGcyqiKznvhmIYfUv+wSHzxmio1I8udqaT1Wn+sKc2SmLX6fU
upr3mLlAiqkmKa6PIiQC2RHyQY/j9b3L2B1+9rpfTg4/BMFtHDyrlxKs4sUvL2pf4LkZPumRWNLK
XMRs99iYhuO1cyFPt+Iiwm910GXlHoX/AG4WctVAnvRKKP6HIo5EFrdRLD1eH9eV5XFFdos9hm9x
5s39K9lmGEFZsH7DtiF7LxO+fB0gDDf1UXFfioWWcGsE8aMbC3c9+mNDcciOasXevpX4Tcxu6I7X
0uDpNkIXlZGkgC2tfhDSmAsFH7IN1UKhGpoP0u48yaQde+GZi8cQ7QFNaP8DmjPnpVnWZ1olxO23
5JLE+DsKtsH47xCivA0mEI185qcfTBAMkKt1+tY5gBNlslNU1G4dRZSd4uQaD3fETgyunFyfJlHp
OUQlxJyLr5Qcvf6QCcIH2Dg2OZbEZaF4zAKGiPT+dW1qG63CD1ct/vw5dGXnAZ6ZatbVRHLwPk4n
R9j/ZLMwR7Iq4gIUWtLaTte7PfHlXE05IBu1Cz6k5HcTIjHTeFD8qhI3YpP9mc8hCydClUdJPTpd
v0+1WU6ZmXieblS3GIcur0TDSVijB4XbFh51C6av9C1N/3zDIqffJLZxudEC8eY5UrGGYWRq8dez
ujlPbNUp95a8IOBtdffUsqH19DbC4T8sjR8/gfO3huRr2vJojN5vcJ+DlXC7M1qjpi5KyCAQiF0Y
obf9kBHw95UvEwvx5Ag9Tu5fBf1+llkVAmR9rU6XZ1wQW3xBeNapBbTrSuT3dnmKc114MGYIZn5G
H7RyabnpTs3WMbiR8IdTWJ9Wz4kJ4vq2RYOaf908QaG3SOC6ny91ToyHjMVaZh5F2G7s7zt6WXJC
sbbNOr8ubb6cbX1ZK1SrZMGsGzhHdbZKdPed8r5+79LJuuyNa9uyUu6d49TpbhnE9YDQ1o8ZDh5D
edeucKRmzmMvC4bOWilcB3wkA/BiBxbGHH59aSvojpB5vq1Z5YtErof9eTAj8rHXzpunCMBmoutr
MaN3SUYlV75ktXi8S4lrJSx9ocpPXUMnqk8DRaVkiNCURWxlVJ8jQ/BwaI++2Tk7oyfBmqtHbw9O
bO1oK23Zm+ocIkLEGBnPGfERlRQQozV3AmRpyeAATc54CLTHfjP+Pa0T1eSVa54A3pMCQKsn/EDA
NUsI76wRSr/gn56t+mXFutd2a392q6+5L48B1DVAX/F/4d1456VJ8wUcZL3ZgxWjl4jZAB8fUNX8
J8cT5AJJq54rXqm6HUzYKcEJSVH9Tpf6Zzj1tze6y6r3UNlS6IVQ8PgBPNkBrNVxFP4X1qCw9tj0
/I3B6et4V8N8YonR46F+AafGuzzgMDfr222/WybS4P5nwbZ174i58GacxJZWouVZhsH62m86B1lZ
lWFnodxBsvplVp/mdvXSc7LDyvjDQRLNoQAk5xc9LnJaQ+bY23sVQXB/njU0VW00txI8y1i23aMh
ZOi4qIgLfJTa7cvnygw+Q+49XZ/IvX6ggtzywWQvXvVTQj9AE34KYROddWbVvtkjWInYOo0h0p/e
xZRyrm5GwEf4dxRVkVF2N1/lCe++v2vZmc5FXw1fXPHeURQ4bGySjYjcV6R+uxoZyMkK0SnM8qOj
LDr02kqHvDxzClYuf0jVTGjHIqiPRUJ8sXm4ooA/FhLf7KQsBGnKQMozr1aghrjTmsH4g/o7pgsZ
SgYmfN/QHJtB2xHPpiyWWH5lEDqJbaz4aaNaZm54R78X2eFac790WOccChqVc+quNQfMfavH/Lrx
YHXYWpUrKUDPaj3RoeGkwtKjxUjxAkWRSH4DJYElltmHVgaQTuOlV8U9H9EXFp7FN5cwCfdP7qVN
8YaTpv9jfu/1J1tg/VBegVbVTO7ru0A0vrdknf3gmioRskzN1BYcpXU2OME4RWLpHigkAWgReDOM
3HtsyRRU6uVmd4I240y4v+fZXCZL+w8DvIx3XjRTThE8a+y4J2aPHpa3YaELpPZ0PhnPKJwiRV5s
E35QQfRsGqQTjrzd3nKj7JciwB+6vuvYOWxxoCC9acbeaXO4i7hMsY7WDge9C7efSqaxpGukrtNu
Id34JoLuheWjrggwvkUEAR2QX9LRGfuiQ2FKT7cNIG8/9FYGxjBvYNbnRUIqOfC/S5KAaSNt3L+5
F+zgBEISiGquEEG7sdvSiKp7xa/vHwPYPvN/aP+mOtMu8+MRhf80XsIVEph3Eyo5tkSZqqMlLxHw
GdsKWacVwgmsw8k2RlK0p77fziI0M20O9f+mBR+q55xj7TnjQvqdMAVmRV1to6P+24gSt6jFs6x+
QoVArGqi7EmDSTxi5psI61A25XaoOj72lsPPbuBdcydMs0N/cmmTjIGJ+pDWJy20gnlwsED1E2DP
PoXdMnx8MOLjsJrWR8ZXWMZVsO8ZSkO+Z6iCDLKrk+ChAXfHIqmilsPIpEyQLx0w4fycBeuqsoUs
cW8fHGa+N+/JSFP3N34uz7ZaksVz9Xx7f+KI8unPewF4uyePCGs5i93XF/y6yxin89K0SVd9OyoP
OhPHLWsgEdVYGhbw0RdOonFd3EGYxJfbY0AX5cDTgpmopvFy35OvK6xjw6Zjpr/8gzb3KROEuc5p
BJCim0HHwgUeYZQD6b38UCRx5t6onOrGeNpJTBM3nQX6O/ub7FrhV0mOEVwa0CH2A3WqZCAt+kgf
8AwIJrBeRZ3Vo98nm6wrj5npB1CHHtstm3PP7cVfqDmjAEEjLpiGOvqI3oJdHtt0a+ILOxrokJQs
ahhP034jHqygdgbPC8Z2VffNrK1TLEeNvPNJBGNRcHTDgDRY9dO16uv7K6tlb17xta/RGGTEhL1x
zp4kscLw5YYkAwChlbLZb/ejdPfzRjwsVJBbyhZe3bo0+lQS+9MNcdJNIyqaz6OsNmPTJlAbAxhd
vhYd+C0sQllcyHlCP52YF2Vd1BJ+ucOz8STi5JEnfK1CafgU7AEKuoZc92Crpa8x3NCCwyj/er8r
g5ymQfV9DMbVUzs24rzd0ue2fW5Bqv+q6rHBGjBYkqQVIFhumr88GkJz7uFiDh1SpRTAmLJHoCxX
Ly62uIaWn9cLObETvhRDiNaWfCVULLrzdtNOemC/3scJJ5TWcFBD0CG7Zf0dLxdLxIUbY5Lc9B/0
TN4o8uJHn5mn4OKl+HMzh9gA1gZUHhA93kIyd98HGi+5VYDF+IXA7CTmAq670Da/GIcTT4mfCTX5
ALJ0CAGKwjyN1Fvcz46KfaP74Oi9Usb8GMW7V0rz5r97+eo+2NmQPp7dCxItoM0kvUmOjXGxznr2
hO3qNi+QapwJl3TamoCv5iFwCaC1hYYiy7gNpMA+sp0QksC0zn7UXaTDcIMQDxVPfMhI5+RROvfP
Rq/ppkvQ4auApJ75Moy4EJmVke0ry61FIui+9m+vT7Ds6rMKOPEtbhk18w3/FgBobplozvaGhnvR
NjZ03XpD79yO6wiSf8TuAXOTFwpHvfaY49u1YnYYP+G4vgnx/LFBbObGJtsBbEBzDzqEzxzbiPb/
tkkjtNbOvGF0ZOPJiKJshKz8tZz/ZHI6L5C1AxRBfk6mq/tQCpFArroknwMnEWTX/ECvRd4Y9oP7
RQLmntBMEYpgFhThJ+Dje36r/mBsq0kN+EVAB+xwKuV42TcrMmYWRCw6rCJunji7pakFVKIDPI4r
HPjeOAXJHgaoGBrwOuNX4+CB5W/ywDLjqBmW31tbsilyC1mt55kZwQfK9EOKKMm9jDU0v2lozFMI
aJEQlVjT0is7ZeulcdtF4sNRxCtxbHgGNnmP/34oQJepQT40MmYs+HaPepIHDBrrQBVhRUxQrKuY
CQsw4Gi9tfKlDBh2LBmZqjZElO/1fb8+McKjaas3LiWS8klFoAN24Y8HOmjXENo1Ugvh9S7kpV4G
wkvspkVOu4+WBeja+ngB3/bJlUGSNRPZ0s9BcQ1P4nIVKYHCTD4Ey17GUvRZUwewqaClJJ1Nywi5
okq5j05LHiNCaI5Y5DR8rOFo16B87v/rnvhME9vh6VM0qfNmNDUuW7eGXR9mNRA/cNJkt1tkFNT5
qm9KTG+tWxZib/LwrL11IQMltmo2y/ENHPbkO0BLcXvJ7x5LIP+aTNOu38UitL1nFvZRZy3lsbMr
BsLHLAT9wgCacG2Aj3agRqQntz04rkQnoVAsgK/iiV1kBINikMNB6x8FI9vr0spo6LRJGxuI22ZG
Ajfl17yr7DM8K3WNLqLpaw43d8Q3cSewjW+d3sxcoUBMJD7oiwbzC5iEQTrepj2zYPd3ySvCSZCA
IfGgBPWFlBOqVPZRFCBj2LdUzPJgRbZtGx991u+JDdjGsCJclyD73pZjnfI0DqmozZw6tC9rrdNU
wItneHa2UXcZDt3o75Ww6rU0OwcXyWbcp4u2JoIJZtIJ4rJ4phbFcbvg9CpOqpQDyL8r2PocdPoa
XRdtub1FKWcTa0GBzN1b9TvpWLph1JHZvb8byaF2a5paixU8hRRPAIc3GGCmC0ROnKSoP7YrPu4k
RlpqadmbcTGNByUahNsCiTYO8+rYAzms3VNQ+xpCWswmJw6tmfDSWocn5H8A7OPWM+lyu03VBWy+
ly1eK99lGSMonWYp+jiJ5gh/7VqXHSL0C3ZMqDVAUWepjPotKiPINWPIB7uTu2rg/gqN98ZBAm7E
gHBtdF5hUaVEHFl/5f3mzvhmOVSAspkMz2cG594Alc3vR20z2xCh8w7OUHmPjLGAPa2QKFzMO/O3
4rt4j5lqdYOmB8qlo+gOsKDjxezCU89qLWByDcVSuzNAX+Q8jeKEzMh6E8paHRn4gd0NA2f8jS3w
hNS094u/LjD6nELaV9IgTox9PJOeKdkcaLXC1szskmRFrI6fS30iCE0OH4Lf/Zm3QyeQSQcWLu80
581y2tWGDom38UXneGgPgLZAVms79nzur/JJ7uhdI4alvgJUA4liGRVtYSXmdlx5P+IFt7ZmO6/m
0JSRiV8R4L7CDsYPQKQQxQkZjyGO08CATL8xFcbBr0UpU+/OVe2kqbiU0cB4YLdD/C5+zgPDe2rZ
BW+hehbdF1rolbhCSn6auVgDBtZFaDR8b+9G40j1A05YyVpsxInFm5ccyASy8YcbIJdTH0XAEizi
S2D4Hpt7g4WzPzyluUCA+fDd8api4AXiLwH7SrJXpz6phdYsfsALkCN0f5He6b2B42uDk6vY+tZ3
pVyprBDJ7437DjKzD7NqmhI2EoaugDhy9euwvwLbltcfOUCliDo0euWo9xdTIn2nQ45E39DMx+eT
31V1pCCtNZDX97RdeTyZNhJ2vHo3gHvDg2k5rR0ONFRejR5Lp2xTLQF9SW9tz1gqb0OzUQdDbmon
8+W61jVuIfD9qYytjmAkHDoI6np5ycz9H1S2GuFeS3oBv6wtycbzpPbeF1puwKL7KJcXwtWf52TG
RaoaJ+JW3fk7CpHEH4T/PatB2ttcNmPptNVSLLBl12bJXxFXEx9ZTXE2hhQuJWRM0FaFut3QrP83
0jU0ttnVcB8X/Uyu3Lv+Lh7ttSt2+igd65n5aO9wba3CYlq+dNGbz9lSAWVA2PSbIgTONxxSlXXi
wzh5z46EDF7PiMVM+N//v5dSVFAcgQECj8cQ83IFtHbmELTFBNHw/7p+5DD2k/0qkdAPeMMzBhGq
2YiCgpQbURxUY271zA1PA1u5bxW+f3WIchYBZz6bWEFFYBvnlB44aq1oUrPCvXs+GZj6YlbengD+
n3UMoFZUoT5u+Dko3M0dpeZoinE4CKoruz7u3HqfyFPaD76sk6/2T7xR8fHkjSVS1pu4tRVw/T/+
QIYdNg/TibbUNmoCToH+h11eD5gS3e8kIBuY3c3fIHOHDD2UxT7YwCFztmpTn+hCrSINNymis4th
xZLLmjD7c1Duq1mLfR7AJ5jWeWfdAU/hrYJwCPLdOU/oZtULvZ/MtHbOMw/8ATI3AJtCCU3GLzgX
/OEfob+HX3P05O0HFD7u2Meo8y7a8iUiZTXzw9C/JEL0nX4npI1D9B3qf7e6Ca5atISp8L4ZAXBQ
eq8ygBqOGI42VKbb5vxtBR8WTHXSSfmES8Eg4bFHPWMC68tBtkyAYY4Fea0Vqb3E0FGSPHD/3/bF
w5IFs+DPe64EP2dTaAkM4X5GHsdCumsdm6zQ/ONBPnAc0RRYtY23igBNNXNLfCjJwjfadSxI4wN3
H9UOcxaHFt+mDFqqoPchk/dAvYeD716L+oabsAPCWe80+alkE+t6Uv4yE0cVLnrKdtTRy+eH7iE4
XVFqldAnL3Cie66ThtT2FwAqUJN2nBXddI8yZ/YlnlDeEQ1DAj/IRBigxZBLykmpTDWwwwtsp6HK
4jPQGocQ5pMW+EUklQ1SFF03UQweDH8lTKa7lkKKPg7nOYTk4n6QypxL596p6QDa9ZYfn32gKxTa
gSq6QfJ/Uwfp3q2tJ1Wr6IIYigV5DifNiMXYZJjNuu6BOAI5/r9r1ME8dXXONJ/FUOZrbFzltrBX
/8ZuhoE96SF4LWU6Yx3IVkuLo2zvTX3nBgeVS+lWPCjTRzQ60Rr7jiAMg4uXVr7z5L5L+eIxKElt
iH0nJqv4rwG/lqYydmeKMMJcngjkITCqI+aNlsbqcYsjvOETZJQMsRcaGunxfEUMACqz7BtjfVgz
JvChHDJgUvrWdIWqsBGEBP5UOHfv0QQGWzkmHgqeK3L1T6OZqYcfiCuPSrixCdF14jUG/ilXIr5b
XuNQwzFTnIq46DuEM9VJ21Zm7MDwyxAR/5IDYuhCUqLtnnSeL/azwcYeKULwowaXZCsl6RC4UQZY
JGX/IAuFL12DQ0uTuDORAyx5JTqMh4LujqU/P7g5wF7SfwedO1etXBUGnEnN7Qc8A1OLa8B4uaxH
p7FK3WPxCjfIvRvpCLqhMF0uZtl0/fWGaNggj1jWcHd51iPtv1/LuV+l1Kebw0fHLBTogsbhk29l
r/BkC4hpH8gdvjnwvBp5tHuK5lASIWTfU1w8HlrGbJ1FdK6FKgWQZMOtgOQPD5+OmFRq+KkQS+Yt
A4ulyhFGPQAYBvkGAHNmPUdSxHYxfHteuqm4z7p8cel3L/FRfBifu1rBspR1D4ClEmRbFKfYknwg
oC0PX6jvvDWDarqAKN2AGuKcUU6muSq08GIkFLXm22jc4QUAlJD1L6EuQpjTQh7kOaFNeZ6sNx84
3RORO7Kt/GYyCtdWlZWqY/KuTUs9R0uaFknHI9aOeHInTOXI9RLbIll6fc7NaLvrzUz8A5g2b/ZQ
OKMatrnNGZUdaHctvyFASiAQu1XIHFn6bNsCVitLOMZtcz293223U0HJngp+PKmPT9Ta/s4AnbRs
Zn0MjSQU6eJZ1pKu07VqvL4vy0tqcjzluxRNI/0X5wvYvHkF2SJKZ3xv0Jro0gd5AG75huxRwGxf
D9MbZX1O7b6BaUO26j6hk3bM6ogf46KbPew1wPIKWBeq6nmtFu+mLnDt5tkfYWWdLjS/JUNmAxvR
niPc607apkQ1gfx/sBIt6zWhxBsgk1WYk7/IDwg0ZticUSXjCYGKcWefzizYF1h2uRJoDNrwJa5R
gBRIhxQTfvrpMLPOzY9e44Et2yYOP9aH2B1Z9VdCzfdxTFkEBVhv/dDmqo2Xdh1BTJzfslwgZpmZ
HZ16mH1pyhuT1MGg/daIcWH+averS2vUMkZ3MYalbcTuWUTXOPntPE4dq1jXeCxacO78A5TKLo0D
QMqw3ZS7z9S3DF66EOxjvG+u0CHfhG5UhjLvCeck0KUfQ3S7rTG+xSTM9WVL83YMan4o8WaMUt/j
ZpC5SoRBT6Bl/dJmqk8VlnYJsfeGc5YpKIRscD2MkrhfXjdXMUxWgN0f04Byg1Rks0pKwBaMxwwC
V5SLtC1LGFRloM9d7nKtGubMUbmZlKCMwhoZDwGoh6uMs23+fRlL6wEDkMaM4edA5XAWgzT16neQ
MfcO0MKGJ5kdnPvMWhXIOtd0x4csnRiQKCjzAL0lF6ibf2uVJg692FuGb/M0REd6bcvd3Czqf43w
8+kmKzHi24Qry19vo6YzrWX2ALC1RWjqz0rCpuCx59umsq1whl7VgXIJh3M0m42WuSabSDGq/96C
ohJ4WnRL6hXR0Zug6yN5QnSqKGa7hGGR/OOMq8/jLFo5/ohKiqQyU+oNYD+P1v4LRf7so/QcZ+dZ
sXHEJ8/8fSEbgBFIHec7lLujGKSdXNt6EL7/PAnPXkK7OtdpGuSuig+6xaYwgb8gY9FQF6saSJkv
TRbGd3qtWV4wdpGwQKQVsJk17SGyUskbLZE9cL8BbluntGyGa0OTHXZuRLi2wpLRIdjKAtXSKlfH
QCdXH4XEqCj3uwGl3j11aq1pMUy4pLlm50p67hyVd1nKTBGUqKLmD42Gc6gZ1UTckQOhuSHHWImD
Y3KZ9DIe8Vej80mJ51uFq6r6WFZkYroDejQe2w0rkFCPdECpaR3FY9YsmgVp7CUHZGYcHKVq5emg
h+J47nuYsaMjYG4nkykz5xxLGY9l+y4adlkDaEwIbKsNDpQ96hn1xg0AGTT9u/gBgH4Ks6O/RYzW
cT0DKB3o0KnniyzOJcaqlhqmHma+8xnfPFWo6io1GcFWtmCKzCC3qG9X5lw1OsEbOXW9tsr6ekGq
j+Mthqqa7hQuKBT552SnPFf0QKwslN98c3zEBi0DBlSIpMm6kIT8qYkAbbK+h//peK99Rvg9vI6r
ujaZzi5pAvH4vhXgMakZ14roMpv+sQ6z2pS9BgNG+7qCaYN+hd4+85sR2E8bG+nqAQFnsCSavu7n
1hnhyD0dN0VkMRujE9vGlL7qp9THYG9SBHWDrk4qY8SD/fAVplfMKIoLTZO8CvTskBsc7hJ2XDBZ
tE0+pk18F1sINuy+W6xhOoIWL7NJRTgdyS4VBMkJ/woqM/syBZkItUJJ9Om+xAf9kQyBzoNY9y1U
tT9Bm0pRdvXBxlLw3vIMzNPH1d69BHcoDUZTqayZLurVvMAPtF1bg3hiK3QPFoao6ejW98VJ21i0
EMwSEN913kMAf5uo6Qvh39Rp6sUw8Pn0NiXrx1x8g4yuBY7Zb21ntgvvVbPzlVxi3AEPaqyY7CVd
TeOAyGxkabYA8736v1HO64aDLSulozcMr/N33Z2+zS7efMbwLNMkbxPydco9KhuTqgBp9voxmdVl
6GPOJru5/wU2poWXohmI+O1eK+4a0poVkHsTjlhvpP3uRvnWYbrvXX6G6oCGvda0sRsBybSnA4mB
UWQZHAucpOC0+Upq2I3WpFmBfWCxAUDWB1crf3RF2y0Up6dXv7t9XrSrqEmTUGP/fPsqoZyVftRg
fjs+mxw8w0UU+yb/TWa/2c3dRH7GiPBXY+Ai+W9nZFPbBZJsFD3eTLXrqCmPXeyUkxwTrkM07Ijw
CvaKm60nlxZeNKzjg3+x6eWMiXQdvSPkikA07siZZhDpN+CO7hZdMl71EmCLJzDiHx34EnioQp7A
GTsOJcHqm7owfy+/yB5Msv/lIuehmfKFSBhPCQjB1OIYQ5Xwk7c/gYjweTZi6AG4UpzioNJ8NNFY
SZXsof7txEyPMAUyyAcLdI13oss/Zw6WzPNg7fmSuWaMRVOB8ms/statvDk/Tl0YR7JeRSTykIdC
IL87HJ6GdKqle3uf71qzojjtvoM6fJ3zGtyx7CdcwdRSVilY1w/NBIWG1xacZ1OXuf2qfe0Mj+ir
fd1RG80Bvrx6Y0rl3/XavkvNfcXCiAkOkVuSo1VxiGq4o6bL0KkYhug8c5rmNzR2fdrhR2yopfBa
WBgtHypoRt6dsz4xuhWElYZPpYMfnpJKvAy+JfT7gM7YriA+ZCJI5VNtAQ9wbLsM1BQl+3+7ZP6a
/uCA38tLLaju5+FudPSYop772y0VTJBWsSInxfv7E+8xhbLU0YfbQGJBApKxDhwVeP6cWg0GWni3
Jm+jjWFDukANHZVvls+kjiINurb8a9Y2LAVoAB3h87V01DlN6g7LKNsvIO4E/WGdZH5CzoetZLoq
WNeKcIuOFmOobsju5cwWPzWd8WSRO2NbXzwAVC2HREx0jpIxdSbedO6Xvcu4+9MdCK7CKCtNpYB4
yi67fGwj+ZzdSgHGNpfuM+uO5RBkUzqD5hNSHeNnicXciUfRMGTIBvMD6exONsYnYOt+UYC4Yd7F
ZiE/kJmgubGKM2/XDqyhvFTT0CHQvxhE3bBKYD+ZKkGOtIRmtldik+Vq2HmvCrz8PjjEZlpIfN5e
dHr7v26/eXSucb1RjA8SwYsCHglc4yL5CKnGiS4ZoyCr+VUMg59TwwBL2VrRxcir/tquS+k9dX71
4efKFHmawM9sQn9DcBn22qHm5Of2v1YuBFzLdrlukqCGL0Ut2YmzijuU82wVxJ7+I68iQYS02j+o
UmrllcJNKihp+cm2teihgPz6QB81HBIG3VFM3/kmPD1vS3H3q2n/IZQHmq8nkCWSlODmc8VNwK0k
uMQfCJoTvMm7XwblszDgMTh8ULZzHMTnAWEmTQYpuc9YgyJFkCfLF2+XMj8VL34LCxGq++eVb/Vi
DOE6RO/56AGOJbc9JN9cBq2oVLEQcmMobeA/W1EjF2yKwdIn6/NbOP1k/20XLRyVSgwzHAuE6ou7
CmuzJNYNp9XehybF7P0sol0WfNFh6QOzRGqYuV4J0o/blI3DiQy46iQP4uXdbZTjjaomDkONn1ww
kmMWfK1cwGhfGzqMCXkH5c188zDLSUFpf1wWF/COfhzuTcrVtV2fRaGuM/+r0WrsUza8uRQDmIV8
PMbqjIcnfu32GQTJTScStc2mVPNhjADrd32ZEW2aZP4hl2sRCEmBB1q1LpRK/R6Ja9p1ydbVVmif
W7KddDAVhpc18nBXNLGrbQQETU7SB1amxcTzDSTQfN+IXMuX1/JEJLJt3emCB2HzD5kgpSUmx1Ad
yTA7sbH+9eTqCn5xBSDWF52douDe5Brsl9oAK/BSUG0Orj7veZ7UFrVQ4ANW/Axyf832hspX3YUX
bCOe7J8q/oQ3z2E8OnZ60rO63gPAr19pC4Qq0YMlzwEnc3lnlDS4fFSsjjy4xTtvJcUY4vt+MHXI
lBC2r+F8JsTUHnVAvo2hfGxfuuoA1teHnJnfVfzBMa2cCky0GfdYqqDgMKJqpP3AMe3ezwz1n1W2
3HxjxrKPl6RYSS84fWsXKS89bBTV14346weOeEK9e2+Mt0Enf0fNBxgqEkUrtKbSfnUvuSsuW5gV
pJo+yfU50IUX1Egat5rsEy5WmM1NjcL5QBNDXkYF2/AFKzt3wvQAh/nsiNhOWMGTzPJ2m4nx1pjA
J/sPSnMnaQC/QfyijcbDH0AvsLr2l6GmhBqmw9+OEWU708J6cNxX+HsyU82ESlKoIl9XI5GMIwYE
i7rBjVNwvLjwmKWfEt16re12tw+fBCqt7se+XRqzpr7jaXRW6RZg/xsYe1or2zKzN5Ub28VvsDtX
pobZN4qFYKgxckAaI6RAXfhaHtCc+Eoiqp0FhNHa+pq4siyA3p3l6NEzo2j1QByHDWPl1uSxYlDM
P0qmz/8zxSKilM3YdGMkB3k8Uo9yCxOM5cPrOEs83W5MfcoP+6nnOhmtS7dXhNc1UeGSH+efO9Zn
R4NcOfkQcGWDO0nq9CPIiaaGwavyhZCiHDFpdfHuwnIeO9yB/R2rGFTzn5+u85/oRPwk8/J7YAQs
ZguwqgBAYbH99LWsc8Tsg00LJMsUH6EasQqiw7/LQ4e8bibEF9QIimV8ACNYzJeISzdrqacbgKoG
fVtD7W+ONINNj3vuLs/BGP5xkZgBaCQKMsPa0h2CCQgtfA5GbeFgXh2a338CJ9qkZjpwmkqquW3G
ujsB4mB7ECXNVoGZt4+Gj81kS0su4qAUsmOO/i4mKWILUaQ2M0JoURVxTWdrUG02QgbJ+w9apl/T
Og4SJ6CZeeV5f61dGldkjd6kZdSgQ9SwYnQ6oH4A+CbS2WW0gVKcWnlVfBMipJ6PjKtJu2btSigT
nh5Ou2IKajVNMkkAKRHJNOP8sOZVXGp25tYSZQt6whU6K0z7of6xDmlrQgvT2ZfdKJex6uGB8XID
PGNdIGLL/FkzztwncyRrxgE4Lld4FnnPuXEOR4z+e7TZVNSb6z/uG9b3GTvnp54gpTHpFclonDCm
qfMtmJdxNYDY1vtSoGOiD4KcFC46CKlEbtwtmykAphrDu3a7vag9Y7tuq5/TahouD5dY8JSah2hg
UI5nEOB3VR3Nzq8lFvIVB73dFPZhjmqwkwAC9ABPuXIZ0d/wWKeXI2akuZUfRi7UAiJAA0CobNoL
TCHD1towKGiwUjIPYbDVDFiMCV/wAYc2jpXhznmPcVP0Riy07brEizC8ZTuSJpj6mSIJouj4RXKh
lPVze/UdZJ60XopcIA0nW4RV8uygL2TGEGmARfdyt+skYDDkXRe4OeIBEogSWAaPgQ8kbbqRZNzm
5rKy2anmpwZfv6k520Cym8xxHDxMN/eRtY4fMoI3gVhbmkTlQTPeL1/59w1HWRCH50sD4/eDcy/w
MWOPOiXC027pERHBGFcvXx5u2UrAsevWn4fK461cwHj/fPSNKqYhEZWR0TyiXvlYqCNFGc2EmHnG
kMhgWrhRFMOT3W1scHzob/IxGeasfVGd69niLPfJWps0G9gvTuTOLB8m5WmCME4J2NTviZA3JLuh
JFEJvkR0wkSUeaokFRtPokwXKX1JkhefbGcXmnCAt+5z2d539yoy113yrc3EqLAOk/iF0HUjFeMF
D5q9HK9hE4qxzRj0EdTcKgAqa+M8qY7Pd38Ve4a/8jhj9bQOUdm+E1UHa/tKH/1EPq4T2Svrqmx2
Nxd6NslQK95kkbb1z+SV01crG/gOvUvcLo853OBo/TyxHt6u5Hzg7O83a9JavxHb4eqvX6znArkx
8y2lDa3RbmI64Q7o+OmtxLXrHobCOHV5ddQPqxS8YK1x8LQKoWl43UsoUUUo9NoGH58gLLliedLD
ZRZLC9RFE0QvADpsNpfR/m59bT1MK6c1kK5MzHdVoQKWYv7fnJFKcgaw6HRUxUGC22twIJDWVY8A
7RdS8uIfBJ7cAX/j9ymiBJfIoNvfs1UVhGeFAFWRdieGnpRB9g/HSk9ngF812IaVptFt1cnO92cM
f6acQbUsqciOcmY8V+QYGEla4ua8YeiUdntclpTq4Bbwi60oDzcvC/tmHHPtGEJnT/9aTMwLt9li
mJI/B8ywzMaPxHkEVMYaEHqtoxQUVevmOm56/9/Ch5pZaWfch5z09th8YaFn55rnpqwGhW/FEhGV
DXocDzeHnR0cAclMH3aVwjqkZswO0NjF3BL2kSfYoWbODxy0vALxwXYcGvq9wHUxWxoYPhKC4qpq
UFM7/CKJxMOh6oLmUgBL9Zmy7RNWGOR+NP8v47YNz8BkYQVpGFg2TLnDlXQozPpVixSEfGzbPSZt
af/mB2UYa3snili2vKOdOmd+ADPLnb7QMbcxen7nC0+VpJBsbkQSpe/MQxYcTqZ6rrUEZ9nANtra
6lYf6AlP0O4uXkKO4Dk8Jk2NkzWde5YqwrndSRgD5I3j+cUA/kRdddafJ8FPXTFQIq8SWpnPNRaU
GzYi9B4xGS0f4IW0C8tblgx2UB+6aP9CBQIrrJSZKSJcfk94nR4c7FE9MkO488LTNq7M7VWU9J4g
cSTcVYAsAI42N+eLO7jpnfX7ILnXqYUALUQQqXRep3vRrbsKiYfwGiOTfesZYTr8mADYyAa6tyKS
V44wHbXY438gC81412evWZaN/keg1x/dJHRi9Qq9GXgjcQ5sX7PI5obsl2BOBjlEZOSa1eKZozVz
jQjKnxMm0g0TeNdbkKySZrtDZdd60jnfNgcBUCv/yDPQ8TwlYPbj3LpYV+qNCjL/T8bGMtPu9vOy
LimCi0c/yrVki+Y0NIR3hGJjt2TTf0oTtL8r+oB6fw8syqTdMY3DYk2bUqwQ/qJQs6d8e/B+qadV
wde8qAalHNN8PQc7zrufP/yT9eK3gdIzeXQnp+OiBE2krmzRN7jAbNxg0GSMuchl6zcsz1BW/MZ4
StmVrIjxS4xaReSiOidGZfCk4ZlaZASXosPcxfLOSSNpg05ruT1CQbgBpgA6bB0bmM/HVtaX80M0
AogVppq0nmskJZp1gzW/6QpRfZJfu6ABQdAo1kAA5aPA8q+BUcD7gl9xn7tE3sNx05n27PvqX0+5
ESLS/hwyf4kuQEkrPLaSjc2aWN8eDswZ+C3ndmP3TtoG2dtBtHR6vc+/Yy1pcj4D6qJM24821BTs
FR2zK6qnvgfuvARnTZ9PR2sJTv1hmxXAwFsCxs/36cUwXTNISRa+EFzC3+RnvUIB+v801zuMY097
0UyoyZnqXa7xirWbZH4jQpQQSmQgrIul34DlCXPDZUD84Ow45ThvzyVGP1/hdwvvrlJxC+ukZgNv
N59P1jtwNKe9nBXu42uavcdJ3J9RD4Umy91VHbXV4HDHTlvjKdp0v5VszzaI/xQrG4lteOcJWpzJ
wZ91aL+oWAve18BRoCot4zSCfbLmzxh0YJP2DgZaAuDlUeMWMb4TMOnYYZ6jdUalfG137GVuxECV
KhG3ywTWRpwA/U1LZsFNUHsq7TMvT716GBcBUyXSLDdeWK+/hF4VWAiwWv5B6q6DoMt0w6HDhpNt
h+qlaT3ILDY0I1WDezTX0ri6zYEYOV9gWsARZQg1vKEFrakfn5UXkhvw8/jbiLd4HSoSKGO7MPTa
S1Uj0jNgJ5zIIBD1dqKj8r6EXOTJG1yyong18nXbvk3r8ScnK11Q3T3jA6yqnyUAJ5j4SEOl9Eay
YVLBozcVwVoPJ2riyyov3dAXO0NMsv5dfW3cRKVwK9goHhjPV9djCnoK32K2WFOLH1bAG7yGrqDy
aav5OE3wdZ/DXzatqWyRgg9wYnAjZj8z16QbbIlo3GzQqCXL0A/wiNb+2SMdo0KK2Zge6kuR3Mf2
xxnJQ9e36V4BE8Bn4WGHA54LX0XWzTvQs7dZxr3ELTF+ah7sUJ+HIvfq9x5uMxFXrGRYQdJbNwYp
IX97vkfi5Mq1UkDf9nSc/ifo3QUav8hxlEQLte9ruIkiVvj1TBLzMDZtfmYIkw8wu1mW0rXHl/vj
bwQIRIPnnMs346fHTKZFZShylIqAxBpB9UATIRzAXTVseu2nSIgK/KTOkX69pCqbHmPPKM93bRjb
XYtQt5Gehi+n/bMvrjxCPBb3HKzZ8tvhE8lToWH6cbESoXPOdlLrwmQSkOThHJnXWMYf4mFZjTVc
KFi9MCV9sCKRMHpciHv1xD6Z5yWADGIPkGA4Zrid2I0buZCRPGLA/Tt1c8nSW+C1k9S6G4UEZPur
dAdElrI8nHJede80Lq0PPK+pIQviRMvUC6FIkc910hJBHAH5N40jYaqpFgSmJh//JMnS0hOa5hQZ
CvVvN107GWCsSaAZl6LAbn+quPIRUFbtgl0tcuqANackvdhDvoEg5CsI/zrsvKhZgQR8TqktGRSJ
2Yav8+r//nrBT4bvZ0n7UIsWPO7DRrPvEJlgFAhxHwpGGa3+4zxI+c6NsQ74Eg3lIfD1hOlVQuGf
3kwwwt6ljec/Bf4L63Q6mlh/NEi47BgT8gkVp7kPJJrnTSJsYIA5S2OSPlHqqjTv+sWQ5KFFBlKH
p5e5ngBgnq2R0lB0uku89obWf25EdF3q8E3rhujXH20lx60VptgzJLIbtlw0VwsQGAn3W5gok1QN
KjqQBJ2ErxLOvTMwoJG4XiyRmtw46FX1loQsafZRTwXfCoxVgFWSB656gH0JYFbKnEVwrZ/ztXQ4
eZ5RuH+SMGXNaFUD0DGBk5Nnyw2I7CTP1Dm+fCJGJhTircZzuaT9jlmhUY6OVaFFeaXZF2mLxuZH
/0A6PbTgDpAcn2VEm7mm7Ub4lCbCmzQvWcjzuDpcdOwMQ2yo5Jnh52pCRw1qsD0ISkIQ2yeBIbSt
F3X5/zSd5RfRUbexFIrJF0Vo3isA/t7gQiWHKTVn9/T4M1gnd+bT0+PkqM1eDDJ8/uBR2PLqaDzA
LL4wityuu7MSEhXQe+cKpiE7IC90fophTaXIk7YI4juh3ThPc/wuW7ALlmi85OyBT8OPrAc7B8Xh
fYuwlWLTWvwbHlBs2wJpM3XzKv4lvlEcCS0QSyGt/kQJvrI72eLiY4UXoESmlf8lc/ceSuV34vbv
6moO8uEjHVLh7NSY1Q474N4rBvhB+sY1qqQGCN/tE2+cJQwaGzsCdtcPQbhSBu3dPzTaNKoQ3LKL
gu1AGD9uZP5+Rgr3VWAAIKafYGSAxGJIiDgiQEqb+VAen5KKjh/CMfEXmOC37BvtIeSqLQkd7xT2
mCUl3Rv6YkwZ5UIf4cVQwC3JVfS5otWWo88veJWY0wvWj1MjqzTvKxc/7krLY08h41czZQA7qPrt
9VXpokoGHUyheQHszpuGaY5Xcfl/aAjEQdVPeoSPN1FHbVp21mQUBRKa/e2yrTNBfetA532UyBWG
XR40JJz57AfdqFGIIMqaKzysoOLaUw87InrTrvMv3SDWnCACobW5q6dVDX5R2OhFkrvS3ONy5JKh
k/L48UrpqC2hELl0S/LDZnCumcriqIe8XQ2Pt8Tu84SHWjjRmt2gyWDyMeL7ckjYn1Qm/mTXmUMM
sX3oIlmaA00/qmb7OLs32ryVMgP5QHUMBejUPfkf+cbpXqrCmmt1G2fHqnis2NyQo0ymqSQ6M6KC
4xbQcSlFn2LrwFPx2zFtnkROLa7kBg1HRsxtk4lmRmzDHcl0sDW6YydVTBnqp9Xog9f02yjThvjg
3fGD8ElkAs0GUkhlv5yIXG6HAJiVNztMUqFt7Na1TY3OHeNHVB86CZ6buKhod+tx74ezxokCSQ6D
PEEQzEfcsMH1H2gE+DeOngDMSTrXHNVlam/GiiWU9fb2RKUoZvQNyPQdyV3KDvnrvh+v65GT3Ur3
9+6qYhu9wzu5in69pjAi4vWEFpkbjn8tMoCPxMS2yZfZDZ0Uo8BUUq008F1a2vqWA6J6orQbRtj6
VBTe6REMOVsbsHcsPUvVczUIQy3vB6r8WKO/I0tDuqRo9Cjvq44RiHH9prZH2GIQ6UOiUW8oj0/7
GKIWxTHJpbUYn9HnunFYOeaVlAgDGbGLRp2Nr8Um2/wT/oebnTXp96nGQ7inWRX4tG8HvG50/7X8
4W/4JwKTNg3TvvMtDDEGaJnS1zfXAlu/5pRL9UR5varoo7OIoxaSkorpZLz4BuEw4+S0nKPIC+HM
R/DnWGOWmW4s7tuXFzno30fF+HFz0PYqnC9MPaS50JUdWcABtcNRFg7XoTSHx4gls6dLL2A0ZB5N
GKz3JzCP9aXgKmsjk2I75uwDf9VjrLCnn4kEih94KEMCjA+3/Onc5yEALzU2pdTrEENv+eHKCbv/
Zi6b7t3FgG4ETqU4EbSDL+QYM3YpF6JunnoRZAtDWVDLeL6ujKDJdIhOFevYl14y+42iOubjHgX3
mJvJQPNo5d1grPzJ/YQzScO1JgqlLIvl1FXQ1+PUNul+5OrLEfdmt5wO/imSd+1eWRZ1T/iF0Ked
TiURjw/0nl84IvYHTOxbDxxQV0jE9mjuCF15s8Dm0aKNkPX6lK6n8A/pbLY/RJOAWJsxji5cjzt5
yfTc0GTpoAGEvCEV8bp0c/nS+S3LhsvbiQjKBRhTVxPy/vsmoh3ycF5rqC7dwgKz+SCS+wxyTdh2
noDF6y756NkvgesVBp1UWqjD5EHsHKWGjP302qfk/ANsDFBbMjTGz2300A7frz6nnEFlos5aOuMw
xo+2k4gM0EmksDmhLxahoRNVC/m643dCtT3xiKqYK7htRJGlALX1FXtWj4HOYhWM2x1rSfHL5jCf
RcULRteeTCXrjnOcxIXSl5CAmmP3MpjozOml4n6Nb2JzpIckAmNs4dnhewqprIzUnaEtdpYuod7F
+yVmULWa63f6kkVbJljPIOSwv2rjbtw0aDNJTpU7G3ZQ+Vz5ULjeDU/2cTScNfjrwPbgoBOQT1iX
OZjfhbn59dKpidzejnXCq/cd+m3uaJgaIL0CA46WpQS838V7wzKtJ7v+d0QQHp/HtdyfduhcOpPe
J3Q5Eoh22un/M/qhEjk7THc9qLplnNN4r7fGeZgxIu2aerWySPQcVfhH7PV4PMjx+wo/IGIz2o7E
J56E99jLlhVVqzUqXswlnazVn62rwtpIY63AVEJZnoYRdHd4g2x/BZlPRpVYhuKXbsOikeunpGu8
YzM9sS73mTK5A8ACnZrWcksv0YBiC6aQtnlQuHTEhJCvphZ83sKqjlzqB/8Mc6o6tjb6hXJ9T+CM
V8aIZRCpC8auic7JamXTNBQmF7VauxbBMlgqzljS3GsqTetdJywDZWPCbVuXzKfSjGAgApj2RI9L
YA82i+TzfW/CI2bgwOl3BZzwwElTQgxUHkusJLIo1phQ3BlINmjOlvLKoESl4+sMBd54rWZPH7AB
wamye57IuYYQH+YTbVCmkoVySAn9mBLIG2MbCC9JUZ34QfbHSU1Itw2WDacffKTFzCZg9CY5qa5E
/xI0r8Dqt8E/YFky18cpb7+46euw76aiO9MbD49tNsZYykh2zjuRkJ/oXv86YCwaLrPIm9BprYoV
LYY3T3bsonxWNM3PRXm3KcahnmInLZUIOjwrLaziX2CsvdPZbmsQa0jApPbNAmyiSqt8dF/lTobW
ZpU2il+lVgT/3GIF7IFg/c0OzjwqIXTRCYy2MC9UUXHv9IOlPwuieoeS2Kn/4QxXNtCinSpgLW/r
F50XZ+wt9kZp7SzCWrhhzDe4b5xZe3zHEUzCFdpVBZcirxcbyqM75p82oR6hZMoOEsKNlM3Af7tr
VKQbH5QNzMAJhTo8AflyFWD80VnJmeQEyp/3Hoj7Yedi+kiCYzBuPnG41Vch2ecNGwABfvvzmh3f
VMQL4TFcgedcbJ4ckwOzDBhoOwaRHHsuRCmPi+r+94WJb4vrFcbpvyjwq5MYgDUd9WZyCDwX+p+T
V2p+3M+lg9qTyBqWKtbgCBRPn+cseFmBIAJxzDl7D7RYUqv7z7Lg8B+SjWOoGfBuF91YMZ63x34D
b2897x9hR6qcLx9kksitwiNM1wJ5YjiKNVpJKYHts5xf3bLnUD3aMHJKpSIrqhD8t+BMK3fAELAG
fLGq4sOpvDaYcoz1AAYygLejUlNbhujF9OUK7HfEXQYDiJU1L0vvNkdkNTpWT1y8HbABQ79X8tiZ
eEjNPAK81A9yRGq9D/UuOYRm/N7vCrpD4YqZlifpU95X3aPFSBsQyjIz/iWiEGOIoMh9NBS52Vwm
NeCK1wXTjSY8QgTySzkfQuUh7x9A8uKTFj8mfnI0eXMWp0aQmUZsz9oh8a0VXU7qqg/UjoDEQwEM
XvY8hsEmqIGjiuKQyQ/fDho7G/wMMg7Ce1OYA5yG8NSe3AW6aDufR+sqW/4opzxII7qDI7JSCORv
za/V1xZ2AtxLSmAyvC/vt3bOWWcJiuyGRoyBFW5SATQgnt43r1jWq8PvlcISwUInWqjcGK9qyGYF
aaJkzNdzmJL8bo/37+qMTNuW4yWO8jv09G+RtJJNupEJ5f4yUXIbfG5f3WQ/B63i+qu+eF0qOjic
0cny51psoXEnoX9P+3hKV1EHhtrJNV0zS5LMVRxq3NtY1AIeZB9ywSwxICxj8lmfGorEzyno6R8r
eYJ1l15NlIA0ccZ/KULOYhNH7u0rfi260346EEySCN9U13XpLoPZkVNJ9ZMUpsvT6SewWUfpalex
wVrqWyzpy0KbXMu9OzAn0h6WSNEi4oc1Bhbr53SzLr3Av+uP1EQH4jopDSzXetDRkK8Bs7RwlvpP
/wcLbXYKCFZ5JOQL3mlQ/aCEPO+tXop7lJY2Xyf56+F/bkQpbKOGnzidFxWzS42Zjew4ZPE0XRjP
RksCebrdeNE/2IsbJssqQcT7Ppzr1d/i1b3X6u5Ncrxs2uigDbkeO46SyHJAuShrEaeMZaZEvA6f
dUDZGBDZSSXAvpvT6gQ4+C3rADkmdxaWg02ozUJ2KJMQakIhSQ+t7cwBSzbi1oyRG7Pxk6dKKtEh
VS312zFLPmxQptDdsZqPm9L8fqi/Q1whInJYvKec5EUx5Qrmtq6sWBKS/D1M9Z32IeLW2SWEg2Pn
g1038SGeJeBYrfyBQIRWj1DgNCY9SE5j0AdX0iUqLtGN4BZHB7tFWx9a/1SA7UU+7l731EE2onXp
gODgIn96RJTJfyt0Qgup0kYw9KEMCTt/MiRyqS5Vk/8bgEa2N57DHxKdqLq7lSx5CRz6gfH51e/O
CiPG8MGc2pdOGk0hmKW2SSHQ7BWEnAOnBvaeVX598VMgqjxSxLTdXMiMgAqDBjZ9FcSQcBGzrLpK
QF4fvw8oTTzqxV/vrIdmStlD0stcutR3MVDWacKIAv2SWQcx9Ytc4vmk3DDeKTNOjEq0VxUHnmHX
aWYWSRtI3uNoLZW7Qr3DZWD55V24LP4UfB0eCWw75JQ7/XB51EtM/gL8ySGZ1H8rYkWbPuaZo8Mh
kNKH/QLWgTcpeOITjmryLr8S3CtouIe2b0uwSiBwFfv+w1u2S4vBOJD/iq2M/nQp83eu0OKgPUMB
cdmZjR5dzT21y+SbaClYW3bPF7Fn7lAZiqzSEMThLcLRPZvt7l03JniJyllncpXHHZ4XBiIpbprl
ZfzSpJ1hhnIBuCkISTGRCWdu8gcpB0NUqx44Mx6fplziyIM34Ab6rwUkYjPmD8F3qpR8i80XV3+U
hhPHPKqABul4C1kK2KTY6uTKL5hI3yPZVHtNSE9sfzoPquxHlEjdMuAB/LBwmNXwFOLMgeEcJa7u
pEXu+ufhiWjkl9Jg+jX0OBBvCrwHxG7z3OoPHCXrTm3y4AlcOaws4B4WzsUxZEqA80pHiOynT/0M
GC/PBgq47AeCeFwOvH6u1AzJAcKa+UF2P3/nZH2blP+CufoiAO0nVD/ePVa6rH60XKSqqeUZhRd3
++TYkS1LVyYgXORyY1NtGIyfpYN1fBf2E5KInvq/HNtGXbSD7qoTVM+Gve6mW/74AX2YaSBCOG0J
sFBMlkAnJHdWdRZe+uhqcKCCENMGWu4rg4PwftUoA3/bRN/KO30gnoSKuy8F6cRYvxEOzGVfXjvK
rdkB3Hk21708c2SOxFbx6yCx/By8rob6GAcXUPc32M5KZk3YT55jCzDYeQ4r8/VtBqBO5iYfnnkg
qIZEXoJxNnMitGbROF+AWmygjP6mmRexclleIwppYExzqot5WhvwOwTb8/OaWCvDGzEJCv7VKeSB
E+KGJFcTHZgLBRCS8oP+6R2bgY41pyV0YYR4WAIDTes7rU4vpWWrOfliImt52GYBZCcwmahXIbGX
zy/3vqYSWCiMcq3rH6CKF85bU3sQBQI0UPPRwtjKedvx83nE8Ekb+6XZM79MeJq09TxduEIoGiIk
Y/4glmv5qIcqpTOVTgz/5lz24I6czyF6wos2RN5LFbNA5SF+RmDBszZBnN4crCttXzUPiK+DR1w+
M49aCNvEU8od0KEIdjva/A/Cxp2Wnt2bCt1wyIrZFoq23RpI/0qIMxd/iBi0fXOaON5Av643IxEd
FoPxy0HMlskYIeYZFhhCcnWz/aPlm0Lat38FT3M9sYjVs01uXol0ReDIGn03p/zIOb6Ty11kqzwq
ZlXg7FogMh4ymeOs2Yd0QXzLjs/ccnmz44UJtWbot6C3NlRtnOL4NQycdiPO4MHxRsD8jwXu427w
ITJu8iop/TcPxoh+hhp4xXnKAbqEUVeHsej8p2/tIlPEN1U+v48yJlvin4rATdarFuN4QtkEw0an
o8TrBuRwbNuDQfLHXF9dNSlQj1aUwb2m2vMRZKdyp/0BkTGCKQLEg552tCPQRk+dt2kom0jbodZl
g3P1g8CALqSQmj5kA4zmp8oMfDb0uTt84h8tNwHRjhXqYFvfGEOhAmlzxKtAzFIxp8HnpFH6s52s
DYw2B32eCAw0MPwew6z7z2pyvpwp26rvpUsbhcWBBD5XwP6EdX1MixUCvK/AkuiBbb2g3Vti28D8
nR7+D38WHhGzGt4psZVRGlfPs7RfaDRqRc2L4Bu+OqvdO5LMN8OzBH6O75TDY4Xiy3coNEwQCDXh
1fxvlDIJ+1j29D1f+fx9n9fQAk1nv3BGJc23Vp6QYOQT3LVHfMB8hmCGaaz2aOTdhuhckDaCcE72
c41qFwJN2pIznrJrH286rZnKh3mNuA9HBoQjH5xZdLxiSAyvkzYmGrhemMq6CfTH84C2n7m6jT6L
IxUg34vvicjd0BXR5usDmJZmMrs/vq9GL1h78omx6RkBpiOGlcK70m3HLKvsDsmSUz+RNYPqrFon
VOaCL0A3wbISLqsY6AuO8yshEqGgUjbiLy3qjHNFq5bUA05hgTGbDKg5T39tE8Z2K7b1aNq6p2Rf
185wLfXw9Eo84p/d4OEA64adB5rIFGDiKe9r8OeFNq/J478nN4nl1GY5VULxDoB4JfNuWuq6Yy+w
HrUc8Q+sseGyi2mNy0c9leXYxo4EAm+D0uMq2n/s9qUW8UW3i0s/zSKtR/iDiMlZjQFT5OQMjN1W
f2XPpRWZcnInKa8SF5KmGe9OOZmVpbqD4v2KEbBe9cDdz0OkrScsk2BriroR7J+HAcHLZ+yDa9Qc
ZHu+FIcsNNLMlmQcowGhWxCHBR3G7yEyt9I0ffO2BBdTcbFYEodTnN2IPkoOaXT7QDecql/s/pgW
S16cJjxUcL55IFg8XzjfkiKUn+EX6741eorGu4B/37Es01pUspNxPwDOi7hYu13bl6DFqgKw+x3n
K0AR/F9YsWWCWoKTGRRfffmgZ7qOhfyE36YuYN88YYfB1iVpkZexqOkLawaIZ8Ad24Rvi4XOP3E4
4WhD6bDiRqoCCu4ommx9UdGwVZ19lFidw82ogcH11cnR28rpTUof2AYkt8WmpfRyOddjAeSRZiFW
oVNHmtOErErVNr3F+TUnOB6xBFWCZlCjbbw3usEf8g1masd/eJiqMyZlFW37pgxWWKuww7nKCukU
Diwj01LCCWkgXvb8KuP0CpnbFQi6wHQ5cciEEbjZmhFIjb0RxwqD5ARudyAfWbagSmisZ7HQMjTR
nomKI6RbiHrNpWBDcsPsbugd5snPLh1AnO+uM619H9g/ylnzo/TXz3OHADxnFN3wFUBpQm4gCNkC
rdH+5IAN6MqOEdsQHauLAHM8pEe7tAsGvs5XZ8uwXKZtN3zdXlpMCN8tDyIzI3JdedKkko/iap80
komGiiIFRYrHXYZMVXk+B6Z9iRsNIojcO2hFFsd+1TQ1eLT7mio9dvQjQbLlgJio0FRRgvR+pJrr
qAokoNa2XoIQfvVAOq1DNZxX9n3XudyuaKVUevf9xPMsIB10sngvlWoPz/HT1Y5moO4QtYnF7GvV
Pfl2G5PlqY4ZzDjWGKsgFIEkDRrJuPTP5iVdA3BDAbgPvBZvHOYbOrql0kdeaUPTBqKY7aAFAdp6
D0Bo7Uzj88IKeYIFaEc9vaHMIjBkuLuhpaRpSL+MyKiVds2ZqLooQxGvji4DggrrIh92oSb1tERc
VHS4p+YwnXHmYW1vqf8j0UBAh/e9f5IWG0uvkfsu3oJzPLUqvSv5kwQo25G7U/16j2Nqfo64hrPp
OnSO9QanMnnvFtyVCC9Vg3yqYk+PHk1dr8K07VeZb6RLFV0ueUTInF7SswsW7o0+QbI4wjNU/tuw
h11ZfgbFDj7gPVQyNQV6MHu64ie8xlGPDW2HF0C9hjB/jw8mzelHWpLe1yB15tCwAq6ID7TcRB04
Fu8pVBUkD7oLZ13gZ211hSK2RpMOrdSncR9o2/BQKa9JizqxkcIiXM8IsiUHcSM9am0ydfGhk3fU
Ai+ZWJjZ5T/xBUKshxzOsLkI6Om8sDX9aSyRnCRNBj+2RDrRk0U4cSy9U2nyyPwPs+kMNz33M1uL
Ezq3ul4wlM/C0Grl7laRzlkyEflgVtK3Z2uMQnKg0RyE4K7QvZqcTpyDLPE4rRb946LSElAHeT/G
9fuZeDDL0fyyqSW4z24+U7AZiZLCKtDL+EABDh0pL7bYrBWZ3E3quE0Yu/ZwVjmMMRAmNJRAviGA
nwD20XF4GQcIi9T/OfRthUwBGdtZ1UDQ1SHGnVc3+XBmSmJLa2BsT+FA9Dc+fVvSJdat1fn22wsM
IwcnFWkBXV1kvyDP+F+03MDzAyUPbd9ueOfDwf8ut0lhIZ6lgJxwte35VYIStJj8aIvaKU6B6Rp3
XZ3UZrP+MrJ3htZCj6hY+uEfVP1QIS/AbbVqX9BxrPSlOO2k1gTLGcbsMmU6i1152TFTO3CqxuOS
QhIyy3qz1nXbsABMEezaJoVAsn1dLw4cpswnD6XRuI4KnFizZeoN2yMTHIP3knU08z4//skFuhLK
QwIf9Pt633ezXTJiFZ252MwV1OY6jbRDDZxPd0eq+D/Kc4OcuOgbbdBtkMIt7CY6hpAP6pciA9Cn
ko824ioAGwafs6ELV2AKzC/bwzsMZqY5Mx9Rchxp4tzpIGQZsqM0N+FuRLlr2SyZJB11Ns0IlJFk
87Z7stbxm0pQ2uzpSg5Fxe3vUv5NvawOe4Q3e4s5GkFmCk2+vXB4v+oD4G+5sPjFjHxFX7iVEeNZ
qpROT+4Bjh8jauNC1rUogmGhAaKhJuNUMH0GBineRnYIbx7P8YpQWG2BNoVIvM7BA6RBh7OsO+5d
GnRWd/C4/ePsdM/WnaN9Z3yiDEe7VSsCI3ltbPNdc9s5J1i3mn9LCt9OHonNXbgfZKiQfSN51mhI
SAaSdx63yCs+Jnv4NYKcx4+a5qfyLOLw10a13WewiVVOo162f2Yalu1r4AkgfquNQFTlzQiLMNA6
RdO1/XelXB4kED6/drc7N9EsktplPWfE3BHhVY+T7UO1X/toKJx8qirKiF6IEs+6ZACR2um7htyM
O00L1UTn6Q6A5QsmpTSHnHK5IQKowRk6DuKpjALZMDDvOwByAQMWYK4t2yE0+bQeSpfEL0mqQ6KS
O5EuMiYvzyEKOTKvHLP+OAHjKMVMt1/zxzxf0EAvevwij7grtRjtavdF9uVR0cm10cWvoj9GHPkU
CjvZ9OPVN6+gxIfgV3jN4+phlFfylIYi+b/7jfKp2QAwCloTw1sFS3NxkByyyFdJf3q3CQey2OJ+
CIvjVywRyJubLleEXnVEGpScseV37RJCDXD6YZQMor36BUStIy7lFwqFkP8ZksqIjWKJorTUXSNv
ipP7DZgoVPeI9FjaldTLE0N/zh8j54YDuvI2l3Xdn6OTPOOUD9C7ZK+wBEEdG0vutxTd4Ry/Lgc7
esShKjeSZrVB2riY5uyaQX1NaVijNZhXKo5XMx2Sk+hecKJ4V1/xi1RVGvBd/VTe6sFpDNUGUnj3
qG55ixluRmznGg+vLKp0+pz5jG8EYrP0ma8KADZWSGqYWJbXFj9m10bv64OZdN6rLFsTGRdN8sxS
58TwFH98hpyg9WhDWNBrJ++yNuQHW6PaT/p9dkAXHezt4NMlVYiFO0Y330a7m6ZO7Qprm1JMlg8y
HmDP0ap/Vmhdog1sJa9zCLDejwEWVTwn+ywlAlCb+VHqX5OlXKh05Zah4XRQtK1gk2qdlsuEKDrL
m037v7j0ZFWv/kcosm7BJRHWdpI8t/MA4TcezFKMzSKmxxV5JsIBnWo0qQLjJP07VwGXsdNIggVA
OejuDojwmujZruNnwCbixDfNlnbFxRT0zBqeDGs65ROIreDaJUCxL+PdPKvNiO8ZweeVUH7Qry0B
8DTiHJs4N9AB4SZPpUonachbcQQHwuiPGpho+cxSAOLwWxF2Sa2bVpxfkdGOiVrE2WF4tdqYuzgH
1R8ZequkNwxL0cXoxNBkLosvzz5TKhCF7EzoGJ64jpXRI/iPdTaGhWBT2OlRipLtzkVEGMBfCTfq
OkOZxO8Sfc7J7BrOaMWcbuEX8OKeZrFJpMdjNF89PCeL83rwB9X0dZIwziBd4xScVkny21KaVcHJ
BaRe5nDfqKKBTF0jV+KKFfzfm0DnpYSEcu1QDF/V0f0//PspDWT5cHoKSGyMj+g05qfzDCykixe+
AwExpIjg75rIUTT12GS9QSk8QfWUNmIrFPsuSg+TeH1e7xtgeFUsR9NfqsjPK3ALu43U9VV1RkOH
VZsaRAY1suzwdTEwRl52FdQzTyArYU+KFqijr8Qe2GukXjuwndRXelmYN/qtx8UuWwkBFexM5lTG
ae/0OpCf2JMIQ1htzmtkh5p+2U65aHCwjuSuBFKoTwJwenveqc8TNyn99N4OOrGjY+Kg9GEL9xE4
LhySMEZUCGvaHmLg110q5S0Eb1jgh/snX2wznmibG+OSBpqIL/NCmUH+YUMmzLntNDlZCHRwxr8W
HfFFyLYcIgZU/mNrV6tpy/NVOGEjgUw0SrM2kvgMB8tMEVG1GMULMs73laCrC8PsNp/+6gPtg1j7
Q7MCgpvMtx86BlZ4Q+X59F97obGGsEXRhZMqYKgA6JRvd2Q7+BQY1ADqOJLCUaIqzlwFXLLiDRPj
2wduTgzj4sDOJSwKLX7yWPjjzCUiU85R9QzSyfcutREXGAYkVeagJpD93LgKV/hb/+oPOZ6HI2Xo
mYBx8d+LKpRGdYqfJDjqJ6aLK3jKkMZzy2Q5Pe9p6Rl6krBYewTnWxVopqgdtDmaoKRluYMORWCv
GhOCNQITKjrVg0cgh43FG/HqP2rMf3LU4LA5Qpeel4QIQsZfbWTayKgX4kfYFuym1EIsPi3LxMIy
+C7Wx1yK/bxfBB2svhvwZ5oWIoEYbYr7jw053GbtRZY7VOZZ0LNa1dCdaquxgwCvjbuAatrSb1GJ
x5pNuO3UZILed6HyZuPMzIbuMRrdS3TtL+HhTRoEa8d9nDFcClD0eTkb7h2CHlcoab4LfNGhstiL
l42HUrx3T6b/DHUWGVckWqY/Dk94JV4EJPN+Zd6P9CVzIv+bE1YpTnUERF5HCYAXMIGoqUG2Dn6c
ZiugPDTiNVGJG2LMez47gl6XwW/ersQwj6JGlax6LrfTzzwWtatdMsZIWWSwkf3K/o3BEDLv6AHH
8nXfaf6O4z6huvT96je2KGTRt7tnZDC+q8nvJ+IbRl+48Fhes8HW872BJ2SwfWt8woHO9rlMZtau
+tPeZDTJp7hdiCx3kUZGHOqJXB7kgifiA4WzKIzXMhAGheCSw465RR4mOe6NeFW6swJPMn2JMIJk
UELChMJ0RG8oYVx862eZDGDMmLrpuZKxVv9BswybI8ykIqHbYeqzfZ+OTP+IeQLp9ECGPe2RVJaU
aQijYeKcWmG5RMiScuG246uir37KFyIRzfgOaCEAPzeMaRiZd9LvAElBw2uYiHiRL11pZV6/wzBr
Px1lbH9x3m4tsRwjWJbu6y5mbexCVFhL+gO5tD33S5irTPVpzRPPtFW/nPJzctCvearLs9A1+yf0
/Oz/LidZi6z1cnfMPG79v8SJ4fbTp8A4+hbNJtLTlkO8RFPdbpivu7NiVlYPh0J6FuDReQLB+cWh
cXz+KNFefzaTQ6nulJakynByHpLicEi1L7sLhQkar2BIgbMtcQ2HnCU2SSN21D8EU6ZaSHCa78VH
yI5RgAPQ4NWzRZ+3/RFMitx0eQN2QANrFbVucQAsn5ua9/PPCKWxsIaJNY42XYiwLd1MNqidszTp
wQy180KtM7dO02xHbV3bvAfTXBxaECUy+mEEkudygbr07GT3vByz/avzdrt4EZQq3gsimZQenIOU
m6aEq8gVVnHyGXRVh00Lori7TpQFInRNPd336qHMA7pnxfk1ILvRiIh2cVffrbAuSj5QHVGmjdDi
+rgOtOgCgeOG4IhHLFxEHuXPLgXdKAl5RNK8ChDI1C5ZuIePUz2pQhQJSlQ7u12P6hG83hY+PNGn
wpHZ5nB7AOGFUKfA5enMo/kDUObDE69LASziBt+iAO0cOC7LDyzfYPZhpBXpA70ee7uKwvCG7+rz
2XTK7IOJr9XSOX5+YbHfQYicLSPeqMaDP/VPg1lWJgyUz9OKBYdscRPS7nyYhUR9SEtoI/Kk6KoD
P1drCvv42MXKbXKWh6x8J9+yeAejnLy8fsepeVgJrUejqv9llQKBvwgueKXBa/c8+ldOqxyRekcR
oVhzNmn12c93rAgXHM8NbFIrQlDBjXxt4KxWpi3o5c8BANpVcyOl9RYbqFShwyU/gy63zS1XQbb8
evGs6Ti9xBu7QY85NNG74lBKO2GPcsI4TCc95Ic/hWn7dLbzUnZ4CsdNRVU/uw3fL/R91iUSV6Sm
EtMoxNFYnho+LGoulFII8ldqij09j+aaAiaQUb+zWbJ1NTRzwYE/Zrk0A5n423Ezna25vucx/m10
EjyTLw294/MPEtExQp4fJl34XKO9jQicxM6MjohBKnrvKK1K7WxT1wANYd+dx8TOnCj3qTc2FQm/
n8MgOC+xo06MiiJLvg9tYtrc1Fmf+8/fnBtqMrAsdzTGUjZQblwj0zF7PEc3xzj5JFQUBFWPOkMf
N+VAFUMVW97/v/MpD4g1KQdiqvXHYdQ5A2It7zRxNc2W5IQ5eVxL8Nvtn1DbVzmg2xrq3YcMnqfG
SYE1c7B4bmSXq/F0egjTOkeg2N6nP+RpZW6rR32f8Imfx5HfmyKTLVZQ4O8GkpKwjA1h1FoggKpL
EkoDoM0krn6lNV8oxsse56q+gXBwyZt2O8qtps7PMEfoP6HjT4CoP1ZPUfAoU/Th1nvDUIA7oRfl
cSrOxBmiIjhugoNJ+DKoD1kNj8eJERKO/OzMo/kWyYqzwwXd5HYrzBQneC4MLYP6Gf6nvizXw19U
K+V4/qSNlH/3OF5OMmcnvySSOn9TDUCckEB9/amKKYIprMUHhIPeLnkrAhggx7UT3Gg04tbdgvpY
vG+IaQ+Y8m/YikKUdlRrbwqF9cyyhEaJHUcgMw22k8vytqwag8nzkl8+JU3yPY8V5tMvfW82V80I
fHfx+O4eo/jcu3obZerHbWBhaqJAI2BwQFmKI6AIAIxjoMxu9jE78xON5C7c+JcDZRsKx3qN05gw
sJdVwK4WYpiaLx2v8s0gGiCQS09orXbapdaPXmNxEVx9mBWAB/5T3COPvQl+6UvTeznYyoK8LNfv
gu4itVMkY9xuryyM8fSq2MhsI16KTxcgUiZqPeRvsrvGlhV4ZsoLv4YfLtv9sd1pHDkTEjFKVYBf
GGn57wKfUkn4cn16oFFIr13+JGc1O3x+KzECpMD7FspU5rwR5B+53Vq3MHPIDLjRZrF6MrpwnAr5
vPwYzjoUeR/LyrCU+kc7aHJgvbETThE5TRmxBglMGXv1KG7juw/8dKPRB8ezEmZVKWqJFghxztrT
Ph4fvGSyJijeAK1xNU66LUx7HJgfxc12vEVr17KIkWjCKRyTycmkBs2hJjFo8sjhses1rorgPobV
ufh3b6q/ZjI2vmmqMxr7o82wucW/b7D13EqORuXuP9ggwZvyaSmPoGbez2OJAjM4Gu2TYkjRBGLr
LTJPQaV1D3a5213GqYzfZMdXXkNcxOUuKuWo0ZGTM+CMahQ8/UTVQ2qimu3r629NaOR+MW+rL2Xw
R213Pq2D8Yij+TvaZOvqZ2KK4kg5xoc36TppPCtadKLzVzBpRPyl9Uzqwpmv6gF1pHme1k0wT9yM
UJ8aDDq4XIoPcL9q2Wfpjr2UEFiyWosqDIrZfJt2v0HVF8rkzdLIm2D24qv0KBVJZzYTDULbanVi
MN9ZhFCzV6QcrUYHPLXCo1I970+xmCVRknwrvZNibhiy+HLHUwXaYR9+Df3BI10X1NXt3VmDAby0
OuUA476R0HRse1vjx8sCo4ieEUzLv0apy5sa6WhtE+0c/CUDB8ZFdJQJI+G2II0GGWFp1Yl2OBza
MYapY8xEsgGayyXZw3lQWOxKrtqI4MffffaUnxrABk1972u1N4WH7yb83KB0UKY4zFyXNHoBKUiR
JdWHftm9NqFHXb+ncmtnUM3Ul91/eCVbeNZxZkxKRE81FS4QsFXcEbk3Tx/5mVzLFsql5+T+X8U6
3moMD2keLiB1+a87N5nS1qSjGbwXwLxsX9Qb40aJeYgmDdv4z+mm+C4DyLf+3bDPwtjHc2UNfRNp
B91hlEi02c91ryfIB+zUlQtCkT6sx4vbHCldP819KknZ3OzJw/IWIoKbneM4xUA4dXoHlq5Nj7g6
q35ofnRz70yt3yaeuheWs3ZjJL+lvxLsRHwWmLU8IZ6hfj3+g+lfJNhM/GbesZn7gkdqfwY9txdv
AEm9CNtNzr5R5u38ZeCkJaO/Wsw2k1qxREdC9dLxqtTRTPsOWnFKfDkY5h8DWXiZREtI5KMcuYW9
XLwZeqS4SGjH9BAxnPfXRbeMWy8gXZAqtIEH/3sfXF0yYqxbQ1BmmDwwVB/FslH3zRAhuq3JuFwm
jtUAK3QmZbEEU1WqSqOqmbMKo3xBWMHoIHDCM3BtM841RVXgoJeFlsXUdDPT8TNqyH6MdGG6uYU3
JO5KLq8HO9S1vZtVq/6YaFLZkK5OjxEucuh2qTyYmCAJpYgPD8vyV4w4RUCX1oSYgxuKbget5N+C
eKDO7VwXWt3hifuWDkE+jeOtijuP28bp/tQTU0sMNri0sdDOxkwpzWJVYs5ucEUzrlP2webKNy8j
vwI3B/kWo27434G3EBQvwygdJM+J/HlPL72np5PnAwWdkBTQcJmPB03HW9dKQPkTX5b8sJT2kQDq
MeUQQqH2YP4Jrv/WrScF41VMGYliLYRY3IJWAaS/jYEmamn3G+2pnB2u+Q6hQMCgd+CdTwmIDD09
sqkE25O2ZAShtJfxJ2Vs36ZYeqxO+NjGMttoOPo7nw7/o1Xdkow/wSWUoPlTqVInHpGz5O8EN0uJ
5gZ0DwhD5iKuoZQbUlfK0eC/OaAl6oYOiKqZWZnkQAgexXRrxKWpru1jDLIYZZ3xtNvmd8cE8aPt
+uTfBH7+pwc4w4gwqX9lWgMIQkhEv133CtzciUF5S9H+t/jLsVr7iOokJCgXZTRyX+xko9OyXLKX
5ssEobKZ2vNmWKSOD6y0q6m+9VrUFFdFpZTyQsk+8PLC9ZdStjnIxd0sk1gOlOhfc3kHHCL4mHiF
m5+5Z1diuNUONdUitFx8wimX9kTirSCP/bzARaBBP/vIOIQBHqfxSjlc1FtmzPok/9pTWQLy4WOz
+QKJTkiCIExv0J+3P5NbcVVeg5vNCfkT0fat5g+Ifc03iqdfkBlPSjTfytUcblXmMn73v3P59gfI
cwChe/T8r2qamMvJ9FOkKFv09ODVr3jllTAdeX5Muam548TVNdacW3SmLn63i044rqUHr8YqBg3E
PCkKFdyeshRFzLAO/o4BQYteKgc5OOhh/PkNtFp9cIQoUsk+zXOuIrlapVyu7SwdybBWINIZ1Gia
H/7MidfoakAiaIbWZUlTLfo0SLsaKxpTfIJxFZjn3MRGeplRI4cqdAa3REE7pO67NPqEQGnnc92/
K0kawE6Sy1UQp6V3HquaMtQyKFQrCfC7FP8NNauA2diRiktdgCB4IQlMjGwvYpwkd2Wpslikr8lH
5o9kD6+Ekm8RPhiYx/2y5s+vRcw8YVJn/UJq19DPpveX0fkIzhjTPH8KKQmOfjmB62WWSphioElW
pXwNJ/18oZeOAA1j2Pwod31I9iyVEoGNepFWOa4I3BhD/sK3CvcJeQ5zc7QsVLON84cDhSukGvyR
tNPuPWQ7LkeDoP6iXuMj0DLemRXEZguK2RAY0OfEvdvNx9l62WLcTdFlN+2gOEptOzdkIPN8Zvy/
uJz+ZWGGuur1esrJZx3m9QTEWKmn1zSVu3Pw+BEeRfRSUFpPyp4nrA0rHwqlNKftvQ4mXsg5FL5V
SZf7NT0oQ7UThFxJVxyBHrTM90N9TS8uZKYE1vx3gB1Zg9JesapCrMYEWIaDQP5G+9TIhGltJ6uT
ktOH4XCy/Q0cNPC2OyktpXckPedlxPr5OS/KBKcMYBv+DJZGx0kJ6SdYUMl6EGRhkfLXqt4k6UUL
7Ou7+qVbI+78lqUa4lYczl5DqhUtOYkvZW6X138ZDhHpeNQDjm/ltR8Wk+nkeknox6dyiVwVD4fa
LbKTdtzO/YmHGwnp+kP3qE/BK0WUZJGk5tfoyJpbb0YPWDTulMCCakfZoaxq83JPcoOqQ682soXm
Zxf4omjFR77I0SkmgOp6COEmWv+sl1kD2tZmrtLfoEL/gqITOlUzVllLTiDGoDemV2o1mF/BcCcf
VkqKt6KrFDYrZmdwpLBPTgpMhqpTXKKPNqvicH1dmE0mMhj0wf34SqRDYT6g3mIBgpq8BHbFfRYe
SSxZAdRYUijIDd0HMAO2eKwxV3kIyFf7MVtvg/8K5kkPrQrfJ3kQTYhPES8puDrU/rcqKgW9RzsG
qsSC0SFOhX3nAiHdSsO1HrkQZmRHuN8b5pkCW5DSX1Yq69m74nwqJ3vq9lBthcsIzTwDij3kECsQ
trkvUnhC2RJJa1Qbs+atmIVEu/+x+KtUSz22QJSQydiRSa48es13YX/HzuBnbHYInzX5IhxdOBO4
Eu4a30huELdEtxsFQlX8qkLzsYag4vImW+Rf1q7GoaPWfOe5BA432VO2xUeN2rqv3JirBu4AS8R9
3mapkKQfFuQzUJiRJwDgW9tURCcRnQdLMXmTviY2m915Heb3UOWABQIf/gpJZC6vEZPh4ftwnhYZ
Y5RuRiYL3edA3qUWY0Drz/VY1A9nMS6QT7E6NMEu4xXTveFEjDf0KcgvvdHTgrZWReBkpiRGmdnK
yJsvZplmzqqZleLtYIkSteoRPDcry1hs1bm3cMT3TgPHMaCVfHzDq94wIs84Pnhz3vs0aFmo5mFE
lIQE+1AXGZQOUf12LqI85QX4vLM+WvjaECwpjFuDgy5ZAaBm8Um2Su8sQ4g8KP7pRVcL+cLoCp8p
nQ6dmPYVd587ET7Rhknm5hOtCLLRZ324q7GkWzlxRYuyX+HgrMk84OC3jO4YfUnp/to7sCk39xt5
/aQy2QxKVCW6wbTpZE1bNgRqeXPe3pOC5kQNAU1IVX3/xpSN/Lihd9DIh3GJYZUG8VCbbrR4OAb3
FBQmoxqpP52QqVR/PO6+4BlzJ6+QysK9TaVS7j7ipu3EwQ6v7Kr+BYRG6/+VaQUdkcB5h8lkS23l
qGrWUAw7j2tJ7MT50aeiOateHdCPyES9oaE6/jh5xW0l9QOccpjK+Pseg/++6J9inJlONie+qkd1
u3xfXNoZMWQ9YzCvyIV3WoNuD4MNny2+0EyeeUkjbO1aHGVyBpBOJy7P4C3d06QlYWoH9xZi2MHv
9DRlfVjz3vAwk5zla4YdblCbVhGy/uRxH7pMj4rERJybjKXgqwwYw01u6Y4gUDUA2KBZT08eex4V
eKRpwM6WcCwc5y3Tiax+ZmWiBHdx/HyKQNPiIkJwOcf8Iwn7R03ZEJphohRlgrkZhyka9uoZWcoi
JzD3S1JgQKc63QBDiPfF/RQpgA4x0i3hEvjRnJnx09wUAlgj5v+bBvI9kvMTjXGvC4NVQ5o+boZt
ju5FmWR17g3bZpf9nqiZgnCHuLVkDEwk9Dm1DcNRnGv87srmP2emk0ce/810grj1f/+Yrp4dxmYu
ixnMa5Waevch7fpxvmF0sVjzP6y4WyaCr3EqSCtDpZrAE2TC7eIxbRhKw0ERaftCJIXGwgv4k9tb
TOAg6pvmtq8uyIKtUqOyKYvxkh6j7xAMC7nXWP72xjieUJs3eoh61BEH7z3CUhApdjyRm7T9d6cC
25CuW9uL2LJpzosPM2nr7/TOxCglS2AkTR5P28Bne2eLKapQTzuWOE3sQ6fSdgGM4TDLFgmjiHKN
Y3utm9guVEhhnkhjYk/lc/H+BbO2/FZArKbytPCbxAwDpJj2Q9UVhrOC+oBLKJHi7+TkDzaTWNn0
RCWvClu2gQQrPe5600+pSE2BSG5ays9uo9r3jK7vVsPPo9a58TZrIdQ2MWpGIaI0Mdll+1twpzQw
GBhjC93weBK5tyVo5Aj+fRRUx8BqXytZQ4VNQkrwZqIYFWM87S6ueyh7BuPOisNFBmKSeqTuoHZ+
VvFy0ldNwIrDGAeC2tWj/RdGTg16K8t70MDLtEhqVVxPyvV0I+5HRqRUZvpA/pm63PHGp2bgIs7n
HyN45p/rYU9hNvDv635l6bunq57I2X3rLw0WN9zb7bd0MwJ/FozKUBuZQJexmr/nyybJaNoI30Ky
DQPaKU4orz8emAdokSFjlNmD9PCEkLiHJJCtCZ69feAmsFPcQW77HdaAQxj7WwoUpC079HZCnjmw
byyJugB3DKb4aFVt8axkmVCSPyCrh6ImZEXYOn30JiOCweizsBJm5m/9P/eu5QTnJWj1skrOeb54
R9g38YeV+l+nlXoX74SVFLMc3ARYLp6NjUAnPYiluxygHQIgMFn4bfk+AjQzsx4oVNg1rf2Ytpi2
vqBBBrRnGLAUsJOyVlNVeDNE+YUUJ6jKetc9SKIclqmS5R0jyap1r2mkRmbTTBOpWcP33sQEBex2
DdoeLTLegJZFrEIlUecJhqedS6Q6qYZj4e4R9+RFuOQH8JOl6z9UdTYlBBap16Gg/CSJJYmV4fbo
TxwEMv0kO7D/F0FrAM6NIl4ia/wCaf44npa1a39c4sMw5yEE4+tgN9++J/Osy3EWvuRtzTooOmOk
uK7NP1ARggRAkmxoT5E4PgxdcUXuPzqZknDCp5mxYafn283+BOD8/iVcopiqRotbDQpQPGOm1YrN
GHJAdFvuUYzEPJgWxaKM7MPoAmNwlqR0/QARz9UCn/zAjKstcGXHjrs6CwpR8vQ3ujdNdKmuY+2B
27o0Rpz4CUgLSyQBfTGHFqugYWJJzkoO682HChEsXCpYDKOgtJSnGK01FZ5aUdtruiGF6tyyKcCp
hyhMHobPKVBX7jkfv+hixmYLDZOVaW7/Q2Xug5G+9TDO3oN2tGots73s7z2kqOuL0vmx6TImkZuu
JZ0PgZk2Fg4XriZe2UMF/HGdtSeTjtZ33/pdKgT8h7Frusujk1PRF3T8l13ZlM9kEPi8VGOcr/sm
Znzmi4y6w7Ccd4I2oDXlFI3iauounZUB4A6f+wUw1hwkaWUcGkjawWqt7UJFr6ZrXbcbljf9Fj3R
CTQDlp3NretJbA4uPQ+ZKT0IDJnbcKeN1XuZfoOvDUl5sFKkc9MKU0AaOT4dtpRWR3hPsE0vzWMX
WFWcZVBqX8UqAcX9Fp2VRHT6SOm8ni3270ntN91LoFDB9wEHhJa4dzSWnlcy6G9W7VbFODoNJP16
DlFkksE8Z97e3EHZc9F6/1gEH5ZPaPx2ZcZIVy1tIiYra012Kf/wqgXu7o3Pyu+KmdP8zCy+KbxZ
nZ6FzlEEMd3jspEOI3GGfhEGqre7CRrQaN0NsXISv4WE3QdqVyRdMO7wFbwuPK+X+ggt2RIqwofc
jPMO9ZWYUSGVcP7sjArj6oR3xl7F5lJAKsPb4+nEyXhYaR0N7HdQ1AU6NTYzmLTWfem29oKqgJ2U
2eIhEalt15nIjIiVAz4iljbKgSGcLtb3/qSsrBq1WFYGV3rkj6nY9eAVhlLOIHTA98y1nMZnwjyi
taAyLYOURD38k77NJ/u9LMNk6BVkVrFnvRaETJQVE34LkuTUSH3PTNgJ/xfmtDTfXnhy4+VK6g54
JWTJ8XnDWcQGcrCHiU0gDY6vChzuAA5Xw84LyXber2NiDSYnX9jFZbjAPWkXxReyxpZPMhE9sbjW
1o9kxwsoJZJprFrjGehcqvBkkeHvAGh9kE3YWeaUW7EcdB5QP7mfjqHLhEB5UGPHLUfHwcLAGeVb
5jh3J78smDRshAVcw8UONU82jX6Sgnkz9QhcZ/CIGInAQIoPc7FowsIq8m/x8exVnr1Qr5ZR7eca
jzYaU9yks4de0Bni0qP6+i2lKck26m3Ks9etWB/FKQbnT42OdHUyepdNpkszq4l9eC7OWpCWp06X
HNo2GvR4mmmqINUdDFQgg64OdLtMAk2NI/XKbBcJUOOGLBuLvAxFLW1P/NyuI4w4uc0rcaMcZtAG
iJvxF5au2oOLWSyJ2SyO/Hd6tKT1hHf4Tqu26imhy/Y3iqiN/fe0QsryobDppiJRqiyYSevoQFdp
6N+ZQjMJ3EAq6FCwcJpnCzwtkloMroScDk19PnjXvOgIUeZ6BoQuiC43hpXkogXqpOopDcjP63CQ
lkwALuPR1oKi5GwzATPqRpyDIzEegeLYL1IHSwLGqyij5K8CccKACTYJqw+s3WEoodp/OQziYc+l
3kOlsvPCwIMlsqYxC7a/OBpWKawIZWgb/TMM6yKGvK86DnNNBz31L4W7gVgNeWiCe6U7FimtZdEf
1cyVgGifS9PrqI3ycDjqxMoD+2hTzWatgMCEhrOnAebotxyoWppEKIdSb39H+OpIz78vGR0zmTw+
3nCwHFQOx3/KGEdlwbymeEDe5P5KLLf8TZODOdHzrTTjCHhiCUmBMiTT2FVEOWtyZ4IrqJk18BPb
KoPSFmZ29+8UO3b3CiYPeYYeQU3mjW7XcyHIV/w6gjGNN9uAU1pvuPAoIoaRH/3IoMvMfVJx4wdl
FXjQdeMwqVO28tdNGVREWI52ga1pjnHtr7oYgG2Hc4sVo28ZVWTI6cIbnEwR5Ad7kuZ/ED3WGYTl
DNxYDuRNsBCw12xlgOtnJA+C5KOYNNyfDVCJDx7mlflhBYFTzhGEXmsfGnEZ4rd88WU6PJyJldhc
Rhphbub8MG9EXqEkoUlCkH2BGlJwk4063X1hrjjWsLgAVk+TNkbf4rbv9Iux5r7NNclJ4S8LfgbQ
mbxdjLOoHzBs2m6WZA9tAl1++BkiTgW4FXJj3yJ2/6eWVxIHpG4TZ5dr8oy+U9UDAFi5cpAQQUX/
XPfNcBB7CmHShKDxhegr/v3rQkzwe+12k4tRZwdZcovxLsSViHb02EWUPYvD3/+gdtCqnaixTjwk
UDD0r62nakyHSwb+9Bgs/9WzgxXfOY271OlmqbFz5y30U75rXq0FpbVU0taRq6OeWemzUF5bvzsW
7nmM0MB7rNivwSmIDIhPVeZdkAKDtDBVoNKC85gltNYNZ/yA4PVUz4J6h/CrgCDitHahdRbFd4FQ
obCC0xuzB+I7B+fVYMOUqPywY8g5HciY8VAigBjkZbGVTkVJ0WdhV/iDYn+PqG/Li6Ty9tTCgS8m
oJogFusseNrn+XiCJlyRSO6gGj9pSCZmde7yMaTxLguWcydxq6VaFqhkohg5TXlMqnCHTKNjh03/
v1BPGyZBj5OuAjecw3IEkiXwad5+FQl7gm73dhoP+4F0/Bet98+Uh66udk0OBuyk1GW5bNhoS0s4
hKIezLlTSvXuLpG/bSybgQxs+KR8lR9fMd2Zh66JC2hfHes/ZmblE5Gn8cHoU8vukbsZmhWLqxMc
DWgvF3DD3HfQf35W+COL2ZCdvGHdDA63MYjPd+m9aSgM5d1lVJIVofroGYyHQxc/TXf5Bn3/218H
4RNZQUWqIU0GriOznEuHji+kBkn+x7RFQWmySs+XGbu4Vi+4guNFO7eM0pL3reWhjphGg/5fRiWa
wh7edw+CJt7lsgTQapUXmsDWZcC4TETrBmuYs49/BHmj7LgSumC7EQFyCCKfGSHONGvQ8IeAOqJe
E8Wz6mwWgKP1I7gCsquZRy95dATCLc+lWmtCnSH9kMCZD9p70WJ585R2EoFUuuyadESzgv87uUSy
0LbQW2qz2dSmCwXahL1VbhEr5hS+qBDdEluIfNS2FruysjHsf1leePkj19urR2XHvO6h0NT0xumr
UA3/0RPLQXHVkSXfPHKp/O7YmnWAnkCOq8ED2ynGHOIBIb4UAhP/vNBuLaluOo+qtmC0F+4HexDL
6+/EdLm4XdUc0m6uqQtx6FvetmtoAFgBZGhfC9xKJOahNpQ7NbOmjZ44ZyVGnGpb2r0Rh3d6YeHR
sxW2chh0Zn5PzmTEMf+0Wx9+lfYO6PIKZQwmrupnp1e3CHk52TfDGBJvXDSL34NLliQ40bC9J6Vm
ZXPNqbpYeowv/fe3I+KgOfTULPW1IBJbmIm5zOnYXtndXDYBU3zDuZD3JXNH8/l8KpouXO+LtvUn
qvOsIRYZ5i7wvZulp39ZSbeJj4Q7r6MUClqaT0oat/HZqH70EuJzVMMzwmwhTnbEgW2QEVM0aAdw
4hu+w/l6yKbl972ueA565GHS1iA9MaRUQimCwW8fDaqmDRGVii2SP0o/FfFT0/bEzRwitLPq/l3S
pN5DtIqQ5H7SM01d/NQf23rQxRikB/LMKtZPpox4L+3Y/e3eMil57YIKR0XLJGeUJaoLAUCgbjMP
nMkiuuLtNuVJDVASncV9sOHTDXV65TPzIQPQTrhHhI6bG5oNAJA8K7yss8fAM1d2ZhagRMJH7fQK
NHWBmFEu+A3kK98hMQFFjZbELb0ApljOJrZ8acVNLiss+6XjEeGMC6dmofbc35GAnUXxGvDj/5CR
sTbVhczf8H6Sf05n6EMN1egV6fjR+wYvEZsfKwdIZwgK2xdhzCq/jy19ErHWW9npXNQJcMSVKhPN
XwFr4Z53cfiyd/6qx4ZE3eSMswDdFZXDsxx3wDQVqKziHxb3XduqL1EzFEVMZxQWJoM5/pms+bIz
jzuEwHrqq3gl1vGPYaNoHwgn7KEo09VB65FfuPX2V7tjivpTWejk9K9GH805ENoBA023bybThr5a
CgTd31DN6fjzBq9jwj3cyCZ9Yguv3JxLDffcQxSKoGoPKdYMTpkUYxYp6ecTR0bz4UoNrG7XCmKQ
Jg+FesS0kp2QYPAmoKjCjk24jQQ2loErSrJj+jwA8eyUCUSWkgkQH/PqQeoY+S0EfXDA8H7RjGsa
LOKvBJ26FrhZMjTKVgJ8mH2Icq7AHb/CM9mYjIvxAO8KO7rwSZS7HBDhzMSTWobtOFxOORxjzbTF
+ntm69QO+Ev7X2wJF/EqDDtGmxk9+m2g7GuPWByCurmN17ze+b6E91clERwb7qobBosbvwJYRPkC
gzDXJmI3VVDF1I4+nJWgG9j2nHp7vc2ZVIpE9SG5UcQ0VEad9zHxyUwuG+CDvk+FuBe7USg2xLbz
9bYRLDFFGm5/yVWjkADtxfxpqmJaCUhwXzyRexpl2eYV6XMM2XJsJ/RgSLriorMD0LDh5L3RCKZu
xeKqmjHmP1mAZotilS2wTxXkyoodK5yI/O/nrScOLsxHfmgquRDVl29//E209MbJ0Kj+W61OEgti
7OILePPE8o9si9fcmR4iRjy9IUFGePLO2heTu5HlaNQ4TI7JEaBGd53sN/k5XwN19MhPhGgtWvMD
Sy4w3d2sYlpkObFhwClmdpyZiNOOh+WvW73K80/zpC/burH/8E8ZlPVLLyfJuns1O7XpvIUxb3FH
3I0hQmZJEf8Oqv85febNXvHE9yswIdArPoSPatJX1SuYieA7f1H6uoTvlh3R23jrWLvknBEcl+Gw
K79WVtjmIbYxWMrpaC89KW8imTz0i7T2VvXai3BaLYT6Pux1sF35jgf8Gic8WrF2Vwj5ZcclbpJc
7BlaHGnXnR33NQvGq2rB9L8rGbktf5AYCYLLD1MekASHI4kWrel7BTPOkb300z2ffRMKOu5vB3Q2
bV9V2bVT9DwJLG7n+0Y4kaaTAYwq8VyXN/My6j1jYQVleBoNvxcY61p9IHfmy8bXUX8zhvYegG4h
BuF3Mikod2zm0lF5vjij6//6WebkVBAfuJT2IJaHCiCFPlAvfub1dM1E9B5QH854+pCa2fLpOuW9
boUv/zbXiYW00CQMTgVj5E0oyeN66xziC8mXCZj5rzBMs1pE1v+EYf9sBBVUOowLhXkEqme38LOm
FVDAGUk2cHjlVnq5W+bwDfv7UjgfZ+EdhQlvAFSMbs6/E6NxE1q8671AuIfduW2gZZUgWAg9Pl6+
+PIm527wR9bUHRIvoiqixn59yBZxsCmIhWtYZihQ8MUSxUA46egrBKnF1AYRX2iKoJ5e9xRYstOC
BdNs8enREOfZWOT5KXNU44u66ZfVNcYb+6D6z0kn7kh3DP3jJwHfHFiM3kt82zQ/HiGmW8c8/9c0
zpdTNDyN+C0HMeffRPNNC+NLYx71+XZ5urOPbmR1DmGwaFtBDD5VTIxkNI0KTxzoLNjbNQR/hZT9
qPDoL/pCxKNwzyaDmy46Q3LVrioUgf4j3sD3fh3E4/BCMtHIwT+FtE9h0bNk6ilCnfs0CPqZdStT
gfplsgOKRjyYwk70a1KjTVG2m2BUQLhHorsbsUNgeODyROlVtstUitFoyO58LwfjuH+s3x09/xwO
ujU6vupDfnh5TyoXv/KhiQuzY29DFQ4Vc4yd81vJw39L92ajlprBDNbLJv4oHJaBShx0edQfUi2K
6/NU0cg1pdUDSHi4clYn6K5JMcl2OTFAByhY0GWmFOg5s6u4taO8R9HGe/wCScc/oUwIZditUEwd
zExJ2XvDZPmUuuxNZHyfBtJzdWLL3XVtITA2XYT5F8iA9xikqOrf5IcUASwRTqw+qbtTxErjeEsI
12M4tSslZRE0nEPaymjdWOzgwlYTm18iCHkXUPuvAfxPwRR4p4sQik993eJBqGhAa6RV8RllQF82
O2WippOOcp42FUGBBg1bLI3DBl9tkot6S82tn+dzR5VrUhtveEmqSbwynPCEAQn1/K0ZgODTD1ZY
GZ55Q1i2+7SJvpLwenJZolxT32fuIOO8RJeYJP8q769NU15PNnnQyjrrInkEOtH5rb8D1X1z31i7
uQkAlHMFYj2zhlNSlGxvcOfZzF91vurtKd38O9OLV5T9hehuXRzDnYvIygL9u8p9XOZ7p5lq/KQl
+fiaAFyvw1NS2kis5gb4kLcnNGpc4QbSJbfqZFNfKXPisyQ+H+YWJoQX34eWXh8e0o2yW0+SgU48
Uzrn1xyj61wgBjQpVxy6VenY33Ng5DED2CfIrcCd0/QEw2g13UnVpr7kRE5TTakCd6GWOHuMnigA
Wt3gv7KDvXCs7qY9E9mufgbLfrXVSybZTscKgoY7ygdFF5pAGU+I5lNtWcdTk6JhDSiECHMI1GF3
V5EzNzLzisNZj0janiuVxmSdPusnlacziPAtmnsnXBqWaNwC5Oz1KfnNHlSxx+jZC5nYNd9Wnyb9
BFugxWYg5RcYkprvP7xtb2IsqrKpc21AbbvRN0aSr2/Wj0wYi3TJx0iSQVoI4eZ7dZJG0K8GXMuM
qMk8GvOpCs0jtlhMy1gL29fcZUAKiCJqjfiA8EtFfKqxjG8TtgQv6nF+NQeFJ7mmzv6PuIZEvmhc
GRGCvx9sYhiN8IYkxU2jvy3GNdnZRsEM8ZQbbTux7RbppfYQB/MXGWk8bzwDdkb46uxg0ncJGKlZ
vajEVLgYQDVfA+9ihYAqroDzgrs4XeVoljI2AkCQC0TVZ3W8j9xmns09QMh9EOABdncf3V4VfDT1
ZwSNFfG2u+Wz/172RWiZMEqwdcOpnh21J7nC2Q20IcHEt9EZrG0VABpDnRB7DZEui4OKw9ijuXmf
AMjGD8qOVMcib7/SXEfx2aqx4T2novv0lHqPiZaey7AtYeig7bqJfZ6qmMwViUnMn5yp7kSbFO34
LrV5tbedFTYcw00Fa9uv/ectT22XViM2DTHAGbOSle2Cij+TAflAvCHzFcET76r23eUbaZrC9QmD
MLnIHszKDsOptN4WVRmfvRo6G2sfr7bE1mxL7TCNqYb6JfVXM2sP83zRV77rTZXdi3LJoT6fc0/v
7LtzpRCBGOUxwSmF4Af5bHxmYBPKSyssuGKLbwvvEn2fqoMhL8yM/8F/6/EpSskG3C6XDLYEAuxa
hEfzh0kzh48XGq9qT7COOu8zyTOLBXPb2JGaMvGSbD03uYLmOBQ/Jybm3vJXD/kRAwa7p5Dd6Mrp
F4+j9rc+mwlXmRjTGedUITU9ZstxzbCjUEGMxfMpvhfso2B9O15b6A3f4Nt3myDE8WJ/RZWEqCf6
TmdmNE6uSWNRWq4Rg39vTkM3RfXp8GtpdKzrEsBWyeoNHBZJ9pmLy/mkgxG8+rz+8+3FA01Ziazz
klfl7zGZ2fS302CHMjAEnbRmLjymZw5Ahexo7FaLrj/XbNB1MLZ4Mqg82lheQ9mH480XjrDeftMf
NQi5ah6o3uIizTV58awbFsj6wgKGURem+KuJOePQhKXle94mYKKethtQJ9mQ3EJFEe01hAbTTmMc
fNhMJT9p0Un9Madoq005GRcISAfOJAZhZdb07Sqqo/Is9w3LB7nxLZAvT2k7RCKLGFHEsJ/JYbtw
vZynOwkLI8P1pppTLPKbT+EoGWtfutmGCCOz7vL9lnn8pp3eWDkqmvb3bUr8TdkucjAA4YcLhyRj
TImiPWNPXsNtmdm/ZkzJd0qRiDlA1tNHv2/BYD4W3vir05RRVbnhYXr0Jb4h9aZ+Ndk1UergfAow
BBihXexIEfUJmcaQpA46l9kJtA24ovnYasZZxAFkTkBObHJrj8od13nW2SI5NyUYVJJfSjniTOlh
UoCUNxzW0Dfn+aZQekAyMkHUOFEpUOWhbmRTZo6hoc5T/SJNVrq+48LhGan8EPwILf1345dJE0hR
xEGQbZi4rBH/4g0O8WiDCq9B5Ax4wJ66WePyAjQJFl4JPAz6xKjzlev5NmKOyq/20wJsddZGK7RZ
+Ppu29Ku0of5bHM1mU1AkEvOMWiCiK8ZjoVyIRfZ8oo28emgz1dDyNDoB2nl8XF7uWmPrhkckVGA
Sqhd9jcwDQE771ytAHNrYIYF6rywe5xFEOwXpjqd7xwK0RZ5kj4Mn8VDXQZimu9qDQXLsGp9pO2n
N9103kE6aH6syP4dbZrSFjm4/UgUZ7q4tH2Bhu4UWb1pG6dNxBdKiK8P1UxDl8ZgGZ+MYbZN9zIR
FWbw4n26Plnw/oWPj1s9rC2LFXafx6MPALhdyfAbrbMAMxP0MDTpcVLWblDz25jOY5ZTItGa6rIm
6J1KUpZWDbmMUvOaeL/nNNCkdKwA3xjRiKRVqhqF/EUJljDjbtac35v1AGgF9SICKpYYyigX6oBS
7Nb/hSKDvce93wsZqzxN165uvETVeRgYovXvRnabIUbREoTBxeF5Jcffz0mxH6X1M5sKFvElk5RO
8MwHILW1M33tECSZIhJIuW6H0RtRpUKt2TtKuuVSvMxSFH1zQc9jpWPXZ5e8Ol6ZjcfriBhgtfk7
bVLabtCrAYEw/hhx0vKSDki5gCqKqhb2un7dEiwr0g7JA5VdCF5uHK5ZRULXVG/uKYp7YtcwEtI6
Ds20JpXVRyDpm6s9y+48/6rhbdx55sUsEgdCK+jEcIepQmY27QyJBrCAMyYSk59V2JVgfgmRql5e
a3wObxqyz1xYK3ObINbtlVYfyvy8NDvz6fGuH5tBpPCNN/E/ANGLdDptj3Fj6ic7NVeNR9nTQTvW
CJntnxrFAP1OPO/Qy4Wm7KLGxg3uWTJ7RYAobdR1WHlCnQOUQPPKNfIW0+9cbrGf387zcjtXVGVS
+K8Rd4J+sYaEC6a60lduMr4RcyrANjak8aiMWVGAJqdL/q6FeFkaCO+SRwgRQqUQW9QahCO8Buuf
UXpAukYsN4cHPsQpHGdumXJzlwgWG0PymsNdJBVqwM9RxodQN5dnq9uLZtLxDGno0rO92Rri+C8c
Ska2X0s3AvlG3NDES3SRYhQt8fFGzXocnYXYD7djmZPRHmxO2IGEtKpdSqiaVnPMXRe5hBl+1cNs
VdQi7UybE6SXYagZ3lsLgQ1n5IaIKsrvfaegG2yXNiUxFSUVO/x0DF78qoNejrHxFEf4fd823gip
NvDfP6JrFome5/aT2iPvVKxtPESybD2EewYoe6C4Au3jB2FiYLiWonGztjSB4fRBxgOLSnuYPBs9
fJXVcZJQqP3ORwjr3pNld0cIPffpWLuceJvN8x6hgUzOajm8TqjDRpstOCFXn3YeJXQbYZvWBJBy
bx1jGx7VPjHPA8bDgzVAe6Ww1EcaJINsQaBjP989ltyBkSWwCU5X5t7r7JxNrFK7PRL40brrbg9m
BalU/TpOrRy3mTOlYwRvVwbvoO9nRjPgQcUYTtA4fkVuf+GG7U93H9qRvhcuH5hvTFUUo2cWaUqt
Vtp7kRL3TF5YYcOm6zA9kRiy7OCgfgF3ABS+7vrIqVQ85zMevQ53+3aiuOSXYGB9BEIg14s2syyL
hpZ95d19PPMYmo/ED77jVf+E0T9ICQjgSJEQIyHadsRt/wWI97JrnUU6kxPo2xMTijDKhWwNU4sk
u/C3dELGILyAuahHziCJDPZYOKXkKgZF/V+Ni88sD64z0NwPCmPuR4honeOqFynjrban3Hh35+f2
u6a1banyPaffHkTUdEifeeHwnnmPaLqgVkc+dQ/npqAi7eWI3R08kQ8nh9MoQ8lxVCvjJiowfHCU
uf4aSIZ5sVWtlqz5HBn1w/0WzjlLF6AMSuZNWXXwIlx99sI4yY7TUljOBEmoN6nmDCen//G586G9
bQfJ5zAU5mUbbQQY2WxJmgYf0DvQrX3Z+f7hkrqtj25hcbbRr5ARTnErl50OtTXf+5NkBCImD4Xe
xuH+Bs2x/NivANMDJ6EqQsCL1X+HLHJ0PnZ77WuPi6TNtSGCq3fmD5OcX7/PjetRYGcume4N+4+9
ks08056G1MKTg10XuLxrlH36VBcjQ1DggHF4N9fRq8vfGTyqnimFpNZi2FvWuXQnQw+Q6eAAS/Iw
d64o6NTgbPIE+fppUkjUfzN7/5MY+y+3Xx8T/0zoSlCD/2UUEicYWpjA51ekskWnS5jeFWPAAkpv
QFrCbXTXCOe5cJ4C5z5C4/fxPL47m4WI0MoGq6zwX8z0s7c6s2EJglreW5yjq7IcauPrjTIkhsmT
/hZDJ5lvhkyDyZilmtlfE/i6YV+IiqCSAvhPvh2QwLCYYPHGu2/3TDqSip51cO3spM1L5JHem9JU
aOqvhnLoCoHlyBlPG7W+BOrI7P+LG3xsAMT97ldgYrebQCxLGyyhS9DBD5HfbICSbWS7a53UCbcu
L4e0slQCWi8Tf3SBuh13ZN7iRd1rqUebUlCsVPUdQ2n2z5iO2AoFwARMoPA/5+3su6MWa1d+lDaD
ANil7estdIcjsSzUDW9RdR+Qy4SdbW87aKaJII7prICdkxGExeXLFoF7vH5Hd7FDZd4lVM7Okod2
tPFBvx4QAwWDMTXY71VIzg6CRvsqd1JK+ugeRS2Vkfy8eht9P15r3gHOqUchmh9c2AZN01FlDUTC
aakZFbdyh/08UBacosI66vPApgEgSk02BLLELh8mH5THKT9tzrqjdsDSWJNpR3LFx6gO4hZpqGr4
k+/6DUrgtKeokzKXOTDwXP6cblFJrzHjR0/LO3zlCedWm90q1au68ux6ws6kxJRZ7zkhnHgY/4hg
pmi0fOiWO95esLsvd/f1Vpq66sT/hgDkwc+NaDYXhYEMYCf0ahrtupjFfFV51qr84w/S1nKygOZD
1vUGDd+AsDLzbY6bpRcYdegIckznPWITddsBRC0f7GZ0qkxuqcdVx5y2tDNDUiYyCR6MO29WidQt
+BqbVTo304jtdSlYWXs/EyTRMgXFxEdZ8tzVpLflarvUUsI4AfjmF91zz2JiO19twl51YptSmSv0
A9GES0aewj5CseaulctZl8huvLUZtrqYXQGNYgZjjeg6PrdhQpcQirkeiJHYjxtlbtIJM1WlpkZ1
/7R+mdbKIjST9FeGyMkU+WToEDEvzdZQpgC+x+KMyFlZaPeinfq4vd5kNZIF6G0Xme826ecOAwhg
dy6xSuz8x9byTmexoiwlIU1h7L1pytROmg37qCBTBm100P2TY+lJSoD9jYEeXHHIbf+Ms/DWsHWf
9iZxAUCg9fKFrLT0tgohKWC3HPPua4RmVgHDxjOGMNLKkGI2rTq8GcEiz8ycf+7k7trIzUb389Xm
v90lR4GTGu7cJiEJ3xQgR8QS7Jds+pt5M5kTZr9aSJLt18M3/Zmwd57fKGEqiX9+BeCk1b35YzSQ
WJpiqmhGe6QR64V36O5wA6pdoSg64SOUiCDaEQBu6/0F7YI/yNE1ny7GLbpumTrsWkG8BF57ehMt
aA9dWE3YfM3W/V8C+/W+/sfT3ihGh1ZSeWn+up7zCMRizifwp4dypH2fvKLujGqfb0bU1bQHpEZA
C9jBYWjMVJOcjhvo7pJTlQ1ZLqzte2ecIvfHDKean97uAHEa7I5CRfs9ciOPWn/1bc0omVXR7BJO
GcNPK6lL+vKBHsqr9nAhD+PjEGm0SAM4vTZw6xwcTNh9KXNSrJIuSPbvBviQo2DcHrZ5CeqnQfnv
d6hWowC0se2fMQn93frmrmeTebWPnJX/V8axpJANrf9ADeJedVAoBXRlt1mNytOzwlTOKF5ecQoV
kRDhfug0cWHR7YLN8vE4dchD09nPuS1d9YlaHJw4yZV10kOBUKEuzT48TFxNpOFk0mxqTLDS1E0A
pisw28MmhsEK9lMmKFatM0RlE9LZCTUH+59t4IOl1R+HCCJNVlyvbWQXHy3EZw2hj2YOs3rmfc3U
DDjd/K8wX2oW/soJM6AF/YxVaTSYseWnNZ+qE05zz7nNXgoECnJSQAASd0y0NHyOkyQ2tSnOD59h
a7CxlN/9IEMv1bAt8BCi76pi7ifufl80k+jjIdYd4YmlZdA6Zqbm/3Ut8NEn2oxX0gb/i4+Kq1/t
403jaFmXbyCLHQVjdhv6SQx5xhN9Ae1d1ofqBJ5aUGbxtTEzhd6TV6L4XwU8bj/FNkggxslF9EGq
SmT5qydXNINcdvO2/FEx8gXm+dadgzir/qs8O5aH0oe/j1feh69UtUcxRZPi+V9aGVALk7WNxKHP
nSsPKMYXFPnnV0BjGK5pioVAkWRKdWGI2voTTw+e8o53sFTuhYwgTL2Qg22HUsql+MdKfJ3aSzRf
j8VUQdE8X7jfHIfzT4BbEotol7dbhLAVqmEhv2xrSIrqadsjzqa1M/xgIpSCyGRYj8L2L6Qd1PGV
Kl9t2ZV94iXFIJ9k+83ckPAEer2Ru1bjlQs2YpuwoZjZWwKyDq+mK/kwvL/tJvkp6zJI/24oj/L6
Bsl9jyAZSYFUj9XMRJBwplYAQBp/KtfeD6ZjWXaR3JVrGfxVRbiVWMzM+yrlGYw76SPVPpF+zltg
fXJYo6Mh6/i6AM5AXlpKbdnKKSP3pak58FOcE8BFA3LyzljlrDtwDsS+X3Ljk7yEk7sIEUEmpQ3/
zqr5GTl9TiwqAMqy3jjiSyjP6/1e0alR56p2W+E4I6T0LMJIqk8dHLrgybTWu8XRt7glhZQdSDb2
Oxd3zq1nQ78vE+e5AMX97bClQKH7Jh2zXIW2lgqQFtIzmLc+aNPfEKP2L4uur0A3zIHDaSyI96hm
O2oKd+/64svLD4ul62nONX4dnTFZPTv70qxVeMZcw/XU4rTZU3Nwg4CJa+MnJiJm8pbrHnsQra9Z
m//myi5tX6S7+9+hcmyI8JsiE+m7OiZtIGsUgtg4el3HemlYFluz7A9BCFt8KctrPLpTXxA8vBxx
JSDblr1Qb9o16E0Fl/zl0V1MtivBC/1lJV5n182Zsws0P8IJXWA1QlYvBISvX7UCWyGsyDKLdlWH
5t4znw/e3OAXLBF4wdgaqW5pFEPoAl1KiU8CRvdYxJ6c4fbyNxRGDHtPZ6Jfe5BsT0fhZMaslBCE
KoiLqTlceDz4PFU6SSNzb4SFOfkfoTCNgZR7/A8IXop7aK+I/jmelUfY90NLmhj8LyqbEAPiWcU8
3wB9dgfxtu02OJpLAGYoEnqg/6bii/Wb4mHpnTZrndtnqfXBrP+UX++1GS5OMa5cwZSeufqEpzMt
d0V+7dH4YseqcGIKoK/ooNIgwYlCqvXMm/sn+Fpjcn7wjDLHI0zES90Q/7rXxuA3NT93i/sDaBci
SG+/HGnTPYLLmpY4H5z16RoUbqH6i4X/WtneEiuHeWieKpOIJA5/Bkonz2WpIEkb/zr3BcoeY1j0
haJcsC2QmL0DJq8qjQNuy7ULWL7Asc+PbPJrBW0OV5TU573kASo5W4LMpU/yyiCsYVSO7dxj4Rsj
6zWZDm55v4tU4wlIna6eyLwMNbgwIakCQVOmCpXUlVc+0plS7l66Z6x5uf9/VJ4jpaRh92/QBCUj
Unz2Qc5FshdiVFNV1z6pEhMp35mAYcuPltlKHYlo6cKOTiGXXrJ6Q+Bd2+wujg3f3CExichUmrbj
f21TGBmdrzrx5lnYDwjZC96Llo6/TjsWzALnE9oZCoJjZUgDBSzSm3PuWbWUI/uU2hAEDiZIxXSu
57/DENrla7VbrDoY3Ky1tnvPYPfrDUAdFWUNHljozJ7swyFjRspCJnhxdounSqfIeXo5k9s41l+9
woGOF/vqbFf0YqXxuS5GIQhA2QkE6PXbCFzWSgh/dCtxch1D69APQVowG5VYJkWe+79WW0IOIOJE
ctSfEE5m/H/cl8gooxn9HQn2hF5g/7Q8/YYFN6NmzUGP0MYQI3Yzp2NrWXDjR8m32Ai80aTDtZyc
fLuLNw9Slqh3XK+JWwAYCartiOFYtyN+TTOPMmrHBMIeYcKlPeR4k8wJ6XMRR1Uzno1S+0Rp/Fpz
PkveFVOVggW+QCH1FfWNXkZOXGlKYuU749YgEtE7q7mcSKBuyjJA04K/dCrEDl7ODtP0gDacdk3h
F/GCCTz1V7Q/oZSCresbI6DGxc++HacKMGWU73tvo/enRPFWLLdDzJN2QbqICE4B7lEbfnnXIXAu
fHacSmNDbruGkXGLawCwyK3fqstTEShuZIomlesu/Wh71Gxh/RR2ychKmCiqneFKO/hJwuS2d5kt
cGCq6Tw5MJ6uy4A7rvJbi8bkNbR0JsmvydNdostRTEvJ7D0OB2AAJuxXdbZ7DFtLqM7GHG9MKjym
V9Muv/FWL51+J3pzPxWy9qry8RjpmTsr3+I8X5c1xsXvVnjwiB8JpjTzwaeRZ1L2RlS2NjPmwLbA
a8IHtW23l35qSSKzxrBavvFjHUJNhOFfKL7BMG1jMwPkn92EFNt5yIo2PBJeHWRDAsylYYDA/C0p
Yf/orKU0htROiBycptawJ3AHDAQYKofdUZFPR+Z2tBMwvekp2ashUuSoFaD1K4gFrT4DCg4FSqvU
QGof4aRjrlxEZttoLjEAsxF10BZd0SSc7qgPPpms5IHkm2Ikb2ZOtborMCI506ozUgq2ZM8P9Yvh
dxyiTBJjzdaolUVY+Haowmj9mc9gwPafxdKnq+9fQuJC1ga+UQYSAChJD4MRvPCm2KdeMUcM60qD
861YWOqrRsOdWr5G7D/CoNo+IP8OgueMxkHHx2E1eH8oHZ/QfLFqOo2vGGjeig8LZURpk/pO8j1x
y7l8zzLBWX2LlVewq1QAktr/x55uFtAQE/lPWiJwmsWtG3cuKQyWsyOsMABuGf6k55z304VXabhA
8ohVh1N5JnaSdyiehUMUfnzU3qv9zfqZVdujx0SYdp72J2LGxafBBkeHzJxpwm/GnRR4CoY+V3i4
xgbHjWIfvp4T/eL4qL9I5Wdvp9RCCmDyRVo5oS4EJFozZQGMp9EhVBSDC3uWWDTg5mOg44XtDNE0
URN/x4ScOhbujDf0NWAB1NV4iw1JeEIn7sRlCucIUOAZ3OpONsJYFCXdFZR47HDaimghjQO0Nr35
uSD1R91LuAAsLKpzyejsmftsYqRqg1/WF6rBJAnQsu2/ROcvPRlYGuxMQKWQXjjuh3C1RZiOggsM
X/IIW1BrtI22QvfE0Lz0B7V08LsW6WOf5Q+XOCtddzGwjozAcqZMeK/ILDxmEojdF2tkViDWfMXw
dZ2Cfe6KdNVZedKiDfXpTeNJKBbParEYfPmiIHYgCbyyObfMUXOUD8uPskHcOwMnE1TJHrlC47UU
/zAQip9+/CGNBHJ5e+oRabkUh+88ldCSBIYNrw+qATgVMkRvoS0p63VgKJUZB3gDQ73wktQY5Cqu
hoqplT39ggEKQUWF+Ls7CLOIP2s6n9Goo2sVNzBPj4ueVRoAHAiEkCc2fr52907QX018pzSfY3m2
35gjL4qbgChq+fYP7nuq60QBNvLqDTQps6KzpqAJQmftPALGrZvD3l8C7Z9yUmFF0zb1VNkx/p5e
906ZOSaG7ZLxFIop0e3ZE/h8rtsZ1oo4iuNp5to6ZW1M8GmS0TmG1VCq6PP7cYkr1pyGKRIjhkyl
Dd6Y6/d4KhziI0vmZH4KFAkVoZlJThGtj3dFGS6eQcvxh9OR4f2XfjU7fMtjp5K9EutL9/W7nvdx
WVxK1Wrqj39J/0z6k6F4lLSm7rS1B0Vxg28wVg3r23CdBIgGa1wilsnrBMXPqG0OXM0RVrwI7thn
SrGFMVXcWCgylM6NrVS3Wp8B0gbRdIlSS/P+RYcr8dNX4qgS65OTgOW87wZV1Kyhkjevsw+fuXue
6Q1b1HN07a3hH2iOMLhmPJ/LLf77SOrqF7KOObI7zQqrLwCm/2Ovwf/HB5hD4/tOdbH9cH3zqWfo
GZ7h5IQBxgZorukJaeRi5jxZDUVEH9hxosylWGzMlD1Ah82e1l9hshzgv1NBJDgmibVbcQFcaiko
uGN0PWRd7x6UilmU42hekp+jhBqnwKQkoFggJV1Yg/0DWow3icDXUJnAhYbzX5/+O9UC9x4kyNPT
lW0YIRrGv57stWTeVdwFsBXETg7jbP+E9xQ8eMl9gXt3RjwFJea8772fIDtKnzdg4fwcUvLNBISk
vp3VHtef2dqKX1JZAeGgTdYwp8ipcra+34LdrMx8Cv0PcswEF305DQxtnwSaD0VFFcEv6PgfIFTz
hEKe/VMVEzvCaRg2yNcD+l+Wktp+dr0QwdDe2ZW+MrG28Y5/fik3cMHJZUExmoNqRHPRvLaMyfNz
DzRj8rgffYYscBi2clUSFWJSBhfNg9V+XgAE6UmTd9J/KxHr3sljWMSPm2EX/Xkkf2BGVC4DuAnh
G0wzpPsEUxs+y4lPUe52TKs5gt58Dy/ZsdZl1qP4MeXaVu859cfPni9vHoLuxtTAM+tcXTILCc9q
PoqTNLudoXRxyvllabhzgTlZG3Y41Xhg9nCUFs/kNam8aGvmsAspTgSLfHw3WdNLjwwvIieKoye7
ucyOrHgZelF4zbnEVqRGvB590dL2yDP+7MzsS/q8CByVotzIMZvELUGZoTM8BSAu2bNZJCMsYjQ5
4W9m6RNxC4WmEqjjuPuh/fXwDeR7dqy7dy6Cq/ogqVH5J7MaWn4di7nu2B8ouP7EDYr162xJZCKB
KR1CyNI9xETg97cgrlnI1OFqnOG3vZPYPQ/WLHQ+rRnFJjTUgUE8KqK6OswBQDiRA1hfvKUMVPGt
W7QfLFrGOd85NlmiFM6E9hQ2czexm8B5n1I3okF1JB8oPUlFv32RhKtidc89PlZ66sTZ5S/Kdt3Y
by7LcoRdZfkadE5Jr4XwXv9XoCjterIjxs/E+boB2Sxthnwsf9q/fmpssXvyK+VmhnePAyKPojXH
A8KwuK2QPe1lB+CGHz+7WlD2ncmNX6YDmEogVIUFIQqtFHbuMn47Yz8fWtVbVsFspMG/bcLRe10e
LRvJfHsGXyjisbhNiFSEvlRvtH2oUVMxqaC57CE5knCOAVwIIUODby3ruojiuu79nJNS2eacAxkI
ox5v9yppJr6iidvOubhyj8ScO0B1/vhq94/8YMENlWTZ4QBSlI+8HdhlAxcjRgFJrG264TLjNw02
bcU9Sm3OY1LF/ka2W+JQk+Ax1azOpD0btxQmv0frZGi0+YWiSuEI4smp/1gGR0SInk+2PsBXzfKP
FRO5pDYcZrzMqAbcR17/DP6S9bUyuYvuFYcdppcmkTNyAd2PtzVygDL5FWZLKg6eLYVRXHOwD/DI
MCPOvgV4fx00TpLPBXwkwOkCmRyLMCkBZaT8J6bD55Okunt1OkqNhOZLxG1t1OCKwwSat3MZM1FE
t/XzbeQiNT+6UfGqTihPhHGRw5h4xFbLLdeH+4E243lRLM5r8O01wFhVYWXznXQNA0In40NLVaYg
jni4HiUyUgorwWCH3WjVnYnhaqmkkEN3r0X6cTeqiErgxwbcB9ECSPJ3Sw3FaOXxj+MIyzpoO9fY
hb9GrrVR6lqR2g+LY4Q+HbUdUB2VuAZL6JmFxnCmA1XEkVzA3qVz+fC8Py8Av8Psnv8kMl59XHse
Tb9CMU3Z1XOTJZBcu8IOKjcJZkRVkLuP2d73idFh9DAil//e05eWxuW6XCkUY+WdrBS3HDFatfi8
LHGdklHHDJduNXjgm91e6iQ4G/vSDK/zWX4OVNu5gUmLvdX/7DOlF6VP+WupMZCu+81nmyl5+kNG
AyUi73ADaCHfzVbOAvW/JyINfViCvkst5MIRXEhsW8gMNp5WkDfcSDkq1sWSu+JgNuM6Wl9IK4eL
+2/25hjUgblvrnbgGc4m8ZHw9FYJ3TrA8TMI64uSXGerQaB/9krq2aFNOk90g94ZO9xyfF0xBcbm
v1HjXi06L1lMDHKO+nZkbBTRHerxxGSBgNuD1/oJtAvxivqeuK/bV0g0JuQbTZPDEQ/X1O8+7xzj
ahZ1uruf2l3Mt51kE8PPMkBr9tvCr2NTagms4Lx5wdPoGChW+8LRowYeMEnOIGwbHjik694U+MmI
iBAzFgNMgduIlVrDW/arlI+cKUDFRLsEA3eVwVl9eT92RI8GXJvXRgtXA/ZpeGVXzZC6RIi9jCfU
bV+0PIQPAZ35Ry8W56bn5YNoL6ZReDUY1phc/ad/ByedhPRiD53MO+QrPEtw1AZddS3CTFlsy0uN
ez+d9ecTtgm27fYlQ12l7qjwT1wcLIRfmKbGYO3cxc98CT0I2l7ofwFOGSgg8NjhVienk+aYqrjo
luGlHNnNJH3shhUM2IdLknQHsHP986XtHZpVQ/Rh6ojhZ5DfCqif/p7pVtkJPrtV6miRz8syx0nH
Gu1gX6dQG3gznCSp4tsztZTItl5ZcpY2/8Rp1Meu2nPiIv2t+JfOKJmopqNwSj18NYVrIlt5ulWL
vfPMqaT+fvHrya/NOMPchyLW7Em1HaoZxmnX2bnFbLpKVQo8q/ds9WGXHr8hn46Lf/m01LcgkFKY
r7LymjIf93mGVfo2oXPhtlsgYXrwDJAII+JPs5KiVmnwRdRibXQNtn91yJRLyLixb0w2M8L9OVv5
qP+QN5zeGyRmj/wr2pDiq1W0TKyTEOdF0DdT1X1s5VpqzhSrx47/dyZHXqtKGg8PoSQdtLPZH+Qc
29WKLB3PBonTKoUlbYQOs3mFm6belGUeW/1WV/PHv9S8nMcjr04C6Elkc1kUh71XrNZoW5dK6a4J
FhdPEaOTcAjCqF7FDAccO4qDxo6OGkEUcsWtFZNwF56X6urqbF3O5uSx6wzOHiS8uzQcMptjZuph
IUCCQzzggF2IG1CpAWPRXF9yk87X9HhgpHF65+g9n+LE2EX2CyOjYaBkhXnjxEqeRS2aaaWGiuAd
FWlKlQinUeo6JCB9NtOvPLwK2yYG2IRuv7WiraZnLdPs3MZQpOlz6E4EmXDfQVGapNoHTxPZOzFY
4PqeFAJbUje2GJCA2EMg/DlhUrCRBFePh18Ilxtwcf+CiFzQpfomgH9uzSZ/1L8xwFykdr37h4df
SxNOidLcith9c9+Aj5Z1Th+iZYUr2SIaoh2Si4ygOoK3SseaHyFYYFUS3NujX1WDqL62m7zuaUIM
GMiwMi41cpMiiglesYGuQqJ8wmXx79qFeUBIzpAR9iNJx1yaljBqQxYAvYQRifTCHiG3AYQmylcH
kpyTt59M6kF2v/0vR+yLzvUbLCKFwoRj+coJVxb5yMKbReFWJeiOLkDChTvV3gpkEPjLuNfZww6Q
TjFZAkwdHDT1l44xeROaz5O1WLCggfkJ2Da1N0DCk9yVLmdiSpALEX5dJ+EJBUyfOvU8ceF3l0Cz
1FB+coiAJZlBkduGYom4nkya7jx2q2T3D+XgdrEVK8yV2fjH07xt2PEbFgDXV4QstBFccFRKVlaC
rSGMmq1opUtp3rcDw/T/g1nHmN5ay9uaC7e0CiR0RaYrIlyqacRn/siJlX1RHQlWu1EIB7VHQhOb
RxDQyCM1QTUr1NHq3ljzzeA6B0MqdxXMWR/fia/ThaCGDaW+FmwpbqYvW9Tg6BtVEflzmBrbsY3m
3c1AZPUFX4rQOfoce1w5n1vSWHtPdkoTiMJaWcTa55SqiSfJwA1tKnHNebWL/s2Xg1cJhg8SQf6A
TUzfJAnfxjBF/4y3ioWBp+5G92vjpbNp23VLdKP23JP+iX15jFui7TFeLG3cAnu9OXUvo9Nql9Ux
iTY9jjJz/COXUilRqYLcikgje75fsYvm5xYnAQKpJ6TXXFx5oKpXLMPscyv1V4helIs+Yk18T1mF
ioT6PcwVT/pb07VOScQaxJImQXjKCw0FnOqSD3tgx23jE/JDrDIulYRLVqkFhypMzUJg34LELvfj
0FWqK73V/sw0KLFp4rbMvpFryvn5wKbaEhCI8PXNwNn6Y21EV8cpIE32MQAmsTTF6AK6uPUtwkg7
joki+zsA1rioCYyGqcdWym6gh2he8h+ZpXrPE5B56EPd6D+JS2nG2gU38VuGCuFh99vTpx92gbqZ
AeSh3XuSzX79+YMPmQIt6+LLNDfl5Th1KDTmw0ijLHU40xT22VN8toK6zvxWxglff2EgfJXlT70z
GPRDc8zocEAeEly3HZruPrlCC4md9Pn+kFz08f5CgaAt3txj//fMbDCZyEYRxB8cqJuhNOH7olNu
8zOKVex/iQTzv7qSoBy4lkilZDTfQVf3vFarFZhnxV2eYc7R5nxKXWWVyXiK8KS5Y0heKI7PwskI
RVp942JxpPwrrVSj7dcBPbHCuksy6BUyqi8ZHSEfh459m0m2mhcuXx4gQPAnI6/isxiPiZ04Yspd
XmvPi5/ZZgjUZa9HjjUQQ9diivSJaQ4G0u6hrJAWTywyMe31ajqftfS4J5YNf3l2brl3N/2myYYX
0B8k9Ps8UfyMg6l4Yrhmy4hE4iNvG6ijD96PHLi2u2+aLcBw0syDT+/nOcE3X6ifRAf+5srvZxXI
vwG53bZwI3/q7/m10U5rd2HN8rB0I8MROMGywz+DwEjrWJ5zOo/S+29P3w4WOUNEibTEeLAbiljn
kW1erOpiXBvKNImgM9Hlv0DtT1WM5W4Yp0XrePR6i7aS9bfHK8m4r0LZMQ4gkC84mo4jyiOiBvKQ
+TR5orkZizIUaP0aiE2AzzcMJzBkQ53tUEP/rfGfBPnlRwbuwb7kOR05SYH+X44ODmXsamHb7M8n
HJ/FEr61WC0XrZ36h2QqlVhrEryjlkPosw9dVl6127TemTcVMY7DlV0P/KpPNB7l4qd3sYQ8lg4k
QltZK08fq3Ytof65yDImZaytiY+bM3ADSmwTrUkvPPT+XrAkiB6KXFlNgdGIKfBe2su1ZLOAF0S4
lhmsUKxnpwd8YgL48/gUUg9Q5AuuUEZUCtaGZknwQSmtSW0YUf/+5SwgVBHHB6g14CC3ByH7tpm7
3e9hyp5qMq3uBi3D1ihm8ujC9HdVgFlCf0fSNobiDcn3kpHVmEa+4Gi2lhaxgJkAXbes1KyUiQTn
rU6WAul3lTYtoZjQWSaFk7MwiXTF5LZbNxyzawCvLY7wWSGwM67h6AyGBlVpSKdwOalh4iBZBtYi
qp1uLqifKZH9niNwiKuoHQHnUDYL4IgWdZm2jZE1yLBJsZelKeYUXIv9UfuGeo3kWiqWpXK5ONwc
qa5/6bJSIOZwMwsURkaP/GbfrkPVNXLRoSiLziHnODobIBeo18hY3pNhGcfqs9h6S/X22DXi5aqk
YshHrraAdQmKSrWZGrN/XRr+PNOspW9lQHQ+pM4batDuk/Y/j7JsfNmwfEkDY+Uxr5ZgUPxd8bCn
xNEgHZbXOv+ZxUaoweNkY4eqnxKfas81r9sFjshKpfn8LLgzqwTMNoYDpRi/FYTaTFqLwXj2czcn
GNJaPqdE+A00s3HKaBiEwWkcIpUtIwIQg7p59t8074hxiLWDZHA49mShOZGXNP6irkTta5/C4mRA
kP7AsWz4fr699blrHFQbhM7R7myaiVxlOhmfvTi5aMws7VhPHTKYtpsJoVII3+w8qVC80p8lsa/J
p53pdDKvPK6/cxJtHTC8gT6+63lnGPTnCEqC7JIWk4c2nJE4MWqLxwA/XOIUtKPj2yppwdd9UEec
mutMGqpqvD+YG0XsgpXCwslPGNEMOu+EQnxwQUoznilfMtS75k62reTkcFKa3IDkdmoh30BNY6dc
uDUKnsPSVUKE3H3tyQsV6m3ElNiAImkgAR+O8D89NjFziWCdyfCSTAc94GSVE1v9heFWueT4AP5K
AgbAUdvHx8y+nFCKfO8g5vJKb02AhULsfzN07HoLylx3hG45Ig6KmL3dfKmmnxWbmESFMJQTN8BN
Wtq+oPq48KDbwDNnpovbeltX7pnZjIlYacs6xE9P0QdPeKuVHUm1VfHAxM8o0+t2WsmvQ7q8IMWG
+YEiJOisOv2HsL/h6dOKitnITqLEKUq3INpe0yums462NaPciRN/gZBwfTU08U/EnM/iyQNJk7rg
z2WldYUNBzF9zwKKmJbMyGkPy4nnnN111gbKvwIaiCC4M+sQMxrKggwtthCgua4OXsvORIyiKgN+
a2BYizCxiKzehwFdZ4tKU86dOa/GiUW0xqFtcqAhdcxLxkxOoNLwhv3MY0RF2OVuulHzLpnbtrJe
tCgqHWrx88o6zrd/RiCD4EOQJJla6FK87Zv8UXLlZWKqQePC5ERmULSS87Uy0WUNr3422AKxTLX8
zxvvGbh50W74X8v60IL4wdueK4lngtlssHBW3VCb5MDF3lGqmPNFOlGHXpzFoDJUmhPGBVK5qHzB
k0SrquA73kSkUgcA60pUUHz+9wbbVNkUjh4DaqKnurNkDgkh4X94WNq/nQfGnVMFAv3NeFcurb4i
QbGJtnM7peLIDgYB9a7IMOATHFPVsdSq/fNrEY4eSmtNeNF/dzHJmIFtT9S4czGIxQd5rTwmSPRJ
lzMNKb9GD6RXNz81jnBWOYnsUyGpNXC/msWVPsoukTpCEHSQyQR0xvGABjaEMXdse7IoBGqGmrNk
2tOw+75HUsX9h+U42pteI5H4VF+D4Xohmv/6jQ0V/z9bkfh36NjGoP3FIKVsEj/0KkM99gcOX98+
kr5w5G+pOK1G3rzskosol1750Vis0Ii/9ubwqfJqEyVSYgQsdWPA6TTRTvItmliknFmxmcHgj/cb
wwd5aw3xI2w6da7oGTYeo23x5uXjQvmKOf6Byqm9VxAwHz19VTKlIuTI1oTC7DvYbMFQLbF0LB/s
Q7FhE44/Hqde8/qGGLHCiPl/QxcS+pOJenEfAmsoUs01kci2Payks3VgfCslI1XSKEr0Aoe1m70f
LkSnG6ZZCWQ7zz6dvmtgkbb+3/o+rJqc3c/7NhoAOgJnvUg7qNIQGKgmbrkwzdUuS1gI7dwCVjbz
tesTBr4DZsb0w7wbVNjseF9oJALaw7BiAM9xXEJ8KzY/6a41ElecjQRdsiCjg55AeXjPY7gc4b9g
J9qArYYN+dFd9I2ustmVsOSl8Ke8OIxZWQElHGgsLqum25c05CajcSt4CyGe3m0RlhAM3vF087IJ
5IzQPYIOs4UhmDjlhksDOE3PAjuqkKTfpIymG8TMfMSHicDbWgSytlV8AxefOkrJKbfF2BWJN96f
1wcSk5hOw2K5CzrAgom4FH2KpGrieE7/ayiPTkn54yAlcQIo9E0R511vmkg0HBFcqY8rCVkzcGEA
oI3Sx4XA/brNjWToHDIX5sG9KAIrMvtD93OnUmSVTj6OIr+Zf15UlD01nzjZU69jGdf/iok3EOEi
Kand23yMakzLH6KlriswhetMDBZXCfFRJp9YiE1Xynp499qlFWV+ESpiAWJSXeUlZQzcA+rNKAH8
jWFUKfV/m5rMMrkufsbMp/fBhE/65OiQdGTTNwv28PMN/QqpC3HUMFV43f1Vq9V2nOSJff4Ex2HI
Xr/XaCKXe59qW1aHCY+oLQSnojnnKArzQNSacrXuImKDkmjB/RrQq92YCqa1RAEomMST+opbOm8b
VAzOOAAXL42yG2zF/AP109DkYaboQLIx0kUoleayOQW+MFhTEg6gYYwlk58o3GQ8yZVf0AE9Wubh
5oZ97rYrRbKdhyQksbB8Ni7ntv0Jp4/u/YYm6N4mld/ZbgWuou5U/SkKWdf/AxjiHkIUDGBxJ4Gs
NBjuog1OfhzFgIwGYCASOakFRitY2mTjhPkm4PHVgH+DWnjrgHjot+dSdRbMo/u1t60PiysPzoDM
hoxXyjyRutk9wco8bf0VDl6WyAfxiCgHDO5FfH1bR/o8sdIt3wcC6ZRssrxNja/b9I183eK8DvAT
Ov0e8M24mttTRjOo0DHr4ZIpedm+Tc9Tc6ky7MefkYNlSMhN5z/jidVqUCkGy45m3s1Z7L1fvT0p
+YsmzgYfxKAqkmYUM6vVn7KbLdN7uhroMX4Mvc0rIKMthe9q8k2jF7epgLAg1kjViTF2tuWrWHs2
tgmwj4/3X4Nk5NmO7AgFwU0oDxm856cO7SqvbRz2Y9ENhjqm7jMZADBi092H59k0fr8hdKkAWZ5L
+wf0xYRhKJv2K7VA71s+9cyiFjZEFh4iT4wGq5wsLrSXbS18fo8oU+H9n/AUN6DazP8IqHhE7sDn
tzXzY8qA8uyIMNsf2OmCJsn/WAG7PMjDxTHGtUWr/99nXWIVycXIGz7IFeRW0wRM0S0v35DkMH/d
gI8UUtY/+IBzgvuPa1uxts+ARBhBtofTJuzr59Q7p7DafY43BZO9mQNieNLzppbUJYb5l1tyV4pb
rblAImpRyXtEO+yKY5ZEDVojHFsTIL0ZhpxErk5/QvZ1aSKy6PD12z4FkAWVwhIIsEWmauEPegrh
8oM1NJB+m/og44q7QwuKZJ9mRhwJTXZhkuXVaL7AnCK9qgVK1E+f8XuE1+A6RGEwMGM9Ogh6zTVN
9d5D1wDHmpR6H5lJQUulD68ZuoH7ygP/lfPjQyJcLs4za2bREGTuHMhkZaJ7gyJ2Ju/g/n2tEKDU
rjpWCAeIlu9Su4TsZF3d1Zui0hA46v8kTsglGjOQcyBAtegfhSV7mbW0jHxpjTL8sPwpLZQv5eLA
IQe6j+eS2N/yjoTUrDXvnq5rEsW0p6cd0JqxIksiyPwtB5m+2TlEuLCmqPhC4dC0CA1pLVsDSJgD
Q6qCSvcO/hTJEW/UNxx8RwOPM8l/OJVdA0WGlHY9R5GepOZN5xd9aF75S58suCOKr4xN8JVsocaD
WcAekEhrdu35R71ZBi6VOhCUhzSBoI8QqLivcGoQ4+DgbCXxijPabV5p4dM/fCWT8Si+sk8j/QGX
DTSVinIvKoqPlllZewIU+3pjF/wgywJ8r3FwlMS6CAzLNoQbZbEwu7EcIGTeUBnHwcOsZ/SDVaef
zwtMLzkcN6r6h0FXB5BPs8N71oYliVIpAg/0H2HI0MfVZQ7BWDvfzazEEJsXz/jJKo6AUOmV1p/3
BhQgT0CPjn2h1TCgulNzs6t3NZwY7PmIi76kjWyTNNS6tEcjiHI9CG62+vW0o7A/1GKlmRQHnH4p
riKWFGPo2+QdNj1u7R2Vw+Z6viyMltTo41ExOyZd5teNm7msCc5fppRz9XEzOnmhfSup1TW8pu7e
zCBb9xw/5cwjrmUA+x1oZFVCsKY8pHQgM7iCh5uEHUs99mVrcF6243yDO9O+VGJqUoPSc5Cubfbp
g+xWkTr0fWeP+XjFHhH8N9dE0eYLPusu7VdIsBBGqm//SY+f+TfavoXaYKm32Y+BbCvVJ4OPd+CP
LnS5ZN8jxNn0/fwoVMbmsUMkvtbdacKGCYMDUDZ2fjDFGpqarKCP16luXsJ269lP+/b8UW2EXZcD
xFuIHoJEZX7a+CLBWP5qpMkgVwdh924gi18wGSuywmL7txuLNlzzLAv4ATMeUaRraTTvAeADK2LO
7gfQOztjpXa+KrHKdU5Z/XrEX6M1LKqSf+jKvgrdDN6y1fxNKA8+GObeWjdKu8WwKlKtElrCbjMp
YTggTxi0k5RWkK/TOPC9h0p0M///BYBZHbDF/wjaOmTGM92vtt6A2lhkbKvkbTR2HPPGESd717bV
4/7lN6wFOMswZM5GBN+b1lK3TQ0Epi+mqZGY4iBgNYXgAKR56Wm/uffIa5rZVVhtQJ30/EIFS3nI
/E3AmoMphmhREAsRce4P2bgnB/wIxnEJWCBS+GF9JlMFuvRV73ZtNEuc8oQQHTiuV7o0DLG79/WW
O6LA5fJhfNGd2i28cCJaQg8NpG7PQHlXTvo02WtNmH3wgFMYo92i35KfkUzf2epJgtlPciVKLyyk
vlR73/6c1jxi2Z+uhdF98FSJ25B26aLK344H5MVOK1BrEKBHh0E7DIM8b++bu9asHanSVdyVChUA
XTpbt1gT3r1UT+9XUyGjuvWESktfkfHWzrLjbYBJcYhAnDfxHjqBcYQ63Kt+2wmNEF+3ABjbkgTg
IpXckwW5KUAHhSFhWU8VFnjMwNIepmiPfB9F3qH1na1Ca/vXUKFDsWPyzkBQsDnujE+y+na9e/L4
YGx1KTvvVnGhsRNHnuCxCY1LrIfsfhqez9D9cxVGFscjah3FuQxN5Sl0fzay6JCZFW1EePCbvHNd
cfB1K6V2unUlEr3ZSIYctGIyT869w5+LKe03E7SSzgFLHyd5T17NYodWaepeTvBE3m1IiUf+DycI
1zyuYsRsLuZY+3Dl3Dv8Drdla/heViJ3T+D7ciC34r+wbqIYthsWAYBwngjjGeiwQrVxGifItSHA
2a+oax0CUBbBD6xK0YH6J25+k7uEKFEQAxvchxiwae72PiX0jJLJhnFt2WWBVEsVv1rlRw0w4n4H
az7N4BZ+X8i3Wks1l5+f5oPKuxGWomDheNuVve9wPo2hHnPzKnUrXRRgJ844kzr9+QaZa08kCByc
ofo6AxHnzeNMXMIl7fzdimxbq/0Sa/czutwC8YFCEpAnMAjWDrTjPV9ugl/ccxBFqxaad8ENOyWA
RD605JTNetTi2+crNIjzHtT+9LR0LIu5O1w79VVKUS0MfmuVhvdXTU3BAsz+3SL+Gl4EW0rAotTg
gYXsNTqbTnFe1nY4dI+GPbqUjK/Po7PzA+nqSi5xRxoeDJF7zPyLIb+qb1ZtmWpPFffjMIotjCmr
7A4RiGmk7nA/DK34oxsbg8urlfbbV4YbTNyLe/qZGhbj5oemI1HFpllyYa3R1kDQ8MGXWnXH/Awp
DrjtqdTOXzi6F5fq6tB21ZLGFrrgu0RA7sXph+Y4L2AfEYZZqyEbY/UnS/9uRpZer8Pn7uUbcgqh
0q0W7NOSUFlBHdnSAhenArPtVe5wgtpllPvLAwzElYXQYjCDIgSgDRtAnPpRYrdWlqwyeHP4vIXA
FpcJRT7vWQyEmz1I5Wm8Ag/XBVMHUcFZCuMVE24G3+4h03FtxFl88iCECr8En6g1zOYWZryfQHBk
fKiv5yqNuI475joOvRYiFgBQKxBOoK3LIoC+GLz1SDvf3d2BiFx61wPX2trRjTD/oajuFBwT3+SP
P/7YQcGSHDgG1CHsf4M0hzBZuODl8kxlggNVXaNNR/hgq483N8O7+Jk8ItZEsH9v0U6EcneBNO/H
gqMYgmZL5NAXryCbNqqiR96CBfpfeZVL7qaA8eR+k0Clx+IgmaFmhnvcivFCo/17JrBwG+cEJYdH
vixNDxQtj+0cFlEsAwiQs2zlnda1lb+k/8ZG3ZUe+qcAfHem29Ies+EiPDERsKYKG2mju/rt6qUL
zF718NdaVlpsaQkd1iPN7CsOlysbZdWW5IY+VKuxRUCgAwMkkDYDWT88DqnULsyGmb/ydAI0PdFf
UHtaA74aNC72e0bARyIDCULEfx0TmR03zTggIue+jxhG4bCe5sB//4HOgir+ov3Pkb2+DbdBQ46B
A4VR5Og7E8i94R0si9Qe2fkC/NP/CK1/ckilRXHrawYbBXjKwQFcU/GHxZIDWCY5ufn64kFnYPvV
VPW9TzO3bYRnN7jGL8Jyp/yiHsWdTn1mTEaYbpJwu+WRfRrWXaPHAexAYzEraDFdDI1FXRimGnVg
QBGwXxGIwoX1V43shlox6NaF07lAxyu9RERubjtVh2oWTAzFkDCbAZhlRogfHwNbkHRTYVouRHdA
Z38P0aN/vpdghrADLeUYlOlm0kMwiSl48iNgkT8NYgugMZTUPzv8FWo/xw+NSlgjZRoyq/O9KbRb
o1lzY6l3tki3A7kezjez8cTKbLTCw5IfADUB0xyppG69Jx2o8VzvniMXh3ScBS/M8l5/e4rRFRqu
YTrynQSgEr2inE7DN0E6QzXk1VwdeN6KP07WGTKdEF/hWdMIr8l1YnNCNXUaQMZQhU0M6UkGXFi2
KlUQ7EqYfxjLxFEhXarI5AQCuEssiusJm3hbm811v4rjImfbMG0ETEq3HAiEAmgOPwLtnZIdN2LB
C1ZDUKcRnfExFC7kWXV9nw7Uv5ESiKsA9lVaOpYJt53xDKmZ42KDq7fGd0QLjPSpJN1XtGM8qspL
50ToFnYrRiwRRZzYi701ZP82mxbSBWZ7r7W7D/AWJFBRUtzkfQC6SIx1N/TSwT7B8vIhyhlo5aew
cRJVTJ6fEUXNwAsnLvDCPDPTzSXIbuLf5ibjPJUh63RpuQexfdZOYpdawzt1LJ1btBRcsNgOS4qd
UfgJzpWA8sfeSAZvEbPhndOBPK3PCWv+bJBYZFTINyhAV/ZqYlwx5MaDquEyJy2wG4liPUgDxdIg
AXbyM7T/phPlj5hL3NNuMjHaKsrfb4bH1DdmcSmCZbT2QgArBrEitMeZ3TFzfLe7mKmUgVA/w4oI
TRGLQTOw5XG6FfPok4s6q8kwatd0XxKwE9sSKuqtOLurTAL6bzuJNd1zOznC+QVqTsTKWPenA5Yg
FlR3T4ZuXoRHjPNx8BLBSAQDGqSilNYMncz5u+VoEi+7hEUa31Oo719sOGHJ3MF7dgAr5AcC82ib
/qyFwtNOJxDyuWy3KV1Xx5mDU1sqd1dqmry3oQ/tQi0MAPjwqf+83ZoOxF+OQ/UVq3ATZ/Bef5Rh
igi/JKftr0Mh0PoD4gPXE1bzsnis0TRtcQfRvQRFx9ulKf/bK5rU6e5OfYwLghVdlrpZCSAYhE9i
rmCTPYDKqYwqbGByL4e1ORfgnjGKogeLKCKM2/uU3HWdawrD6xuSya60quZcDbMNe9Cmcnr2mGX5
ozqOeEZIblINytT04iG3DH71w13Rnd0XzTfPCOfYqesifGWEVSM1uSgXXk99Nd3iguRMWtecW9tL
+Q4sM7+2FheENM0TkAsEx0J05drJcLwQeJuJ1BGooBUyQop2aIMRJRpGdV0hOHqOTUrlO5L+KPUM
KhHcJzOn/zKsJTGjVEKWaBJBqWRv/NtQsY8aL5XzA+3dEt/AWJQpaEGkCBlOu11LuxR6Jd0zf2mN
hRKdCn60de0zyc8AHwKtBlPGkMl56rVYP8rSeY1VBBaugwaryLupcr0LsG0Y/uKWpHNW/bQA2Rla
GiRzrBfDdmXxaWlfGbg/UnaPHuQfLGm5ab3fOLe/XVzjYRXnfPpCx1kE1lbz8yM4HulNMTBUPsr4
O07YlUmBaE4ExqgmHvSi/uuoYdbsiNknNrWcX48/g8o+hDmjqhOukLrN1DMGbx2ooAuReaz8WC2r
PGnrWHf4fT5IZVX/AUWYxSQ/Ih+ETgiax7WR76ufPnkaU+GyFFosBcWSVWmQyP31EfcRt3sxBwGj
Poou2bE5eJtYx4m4ay2hOR3mMt1z3k9HT5MPNctrQ+hFFY0rx+I92Ss5P62ZsmYuNN2SPvVOxf7H
rqWtppFXrrQBEaHBUbFhWSRxV15N6N++xHZ7BwVk2uLHFvuLTyjfmaSFxN8d2UcPZt71iIy+cNZq
RyGND+Itq3EkCKw5W1//wUKeoIoRRaiD0ph1yA2+OavzarGw9nSqhOMGxlIAzZIoCZUp7LO58Rwp
XQEO7c1bTZYtOr2+u6og/vG/qW57a8P6ygBr0qA1YHZ2MizlHeNfuZCTppJPY0C1HAYDB6leRYwa
w5U0rImeQcXdZphhVp5eUoT94Mgp7vB+CtQu4zncHJt3Hx6O1GpN7/hT8RdepW8KyUOPL85MeiE3
nkw3DT/8NvcJaIfYrKPd0Xhd8Qi+2S3mdyQRurYUtc+2DS7urAX/3cRqotTwEDMyG6JYOQaakdKc
/WuxM/M4up3R9tORZenmDdCyvMdby9yBWCHNyjG3Bcg+j7ZBsuH89Yqy4lM6xmI5tXhxDpMgBX2u
Kk/ZQBIFWOWIiNWaGYDvlcI2DGlktUiUycrp4rnJIC/Z9emcaZaQwYI7ZwYNSJIsiQr3Snpw8mQ1
iE92Tecwji4q9JJC+cIeAGKUNJvIxEEBX3FxkudqEIaOl1MPtDmJZ8vfDPm1JZ59F18ObuH1jfat
1c4/RRo9cfXwDssjSuR2ZMZKOuYQghn2qMvV83cFxV34xUw4hTQPvWm4P+AdT4YI/GiejlQftQCo
uKaOKOLspprPWi63rctVmz4qVSlR/uPCY3jegrUGP956THmmNj6lZHJS+Y6hZIA2oweBWpgYi4E3
V+REmwwYcAfoHnkVYoImZt97vGFyKKPpnKd07jb4IDJFu0VxlO9BN37vAevQsHatVZz5pt3i1fUZ
iBrUCdAM2N/cfgCXHqoLnWcfjrRP2SYvrsOo2JGVmA72Lnu1SNt0W+IFWo6aptn2/PMFXVHaLqp3
cHmqs3AITRd56O4enET8k1NFhoVeKmyNAZhTmxpMqsYrsTgO2uJx57QsnUSNtoULB+RWe9tGE58G
k2gCaFiTxcCmEyXngoKZcx7IN4A0DwUNIC9w6yXlQMMjII+YtM7SH0yZLS27QnCCyuJcXIVPM0dA
Hhee45Obf4DMPh80noOTGh5c3aaPNu57v6ZwIeSPoWDsOjJLQdPT1V2gZiYJKvZfAcvgPuQ3NOeA
/AhKrly4d8xmGyjWgmn3x6uqD9H0+hkCJKZo8Za+xxy+sri7p3Ownq9UC+p4uIxllUDYec7Md96U
VU/9QIXsiuRT3ByjvLHCpH0RtBnU2jTmWL2Ns0ngsbBRO1aUBAkLBnihDlI9xCD3zBw/tQ7v7lA5
sDgBqcPHE/IzQWarY7J5W4hwfqCW8C+k6mNELa0DoH5LlAmPBPo2w8k7QjryFOVdMwTsbzd/+k+i
Y0QUsYs7D1TXNQlLCLm/2hVZZKoChHftG71JotuBq1o10Si21n1Eh3ZOuwP1ema14kRJMxbIFAGy
npSdTLKP+t9RiMDbe6eAjFbOd0Ph68A2fvqdSHtE4UOSAX3BgcdcHGXLGuuiHkDje7HU03HjQNsn
ez98z0KZiyYfvWScInhH/Ywg8zDX8k/mN0N++BvmyK5oUrfCWg7z5DbGZqA8CZQPUmjcbU6mE9+j
HS644fY2FHjA0uli9ggbbR6JyUCTIbKqZm97hvxYAdD8bXLP5U0KUJONn/UYpwWHyZf1yVCIf4lp
8cwJz1oSyIpSP4ramRZ5DuDjiPCgMTtg0w7YPNYoycJerTjYHI+W2mqQM5Kvw2M2C7xibfIsf1jw
0R/drzrxJBlbkBgv2L32Hvdj9W1MmUXzObWaoFp7ry7rdQQmMbbTrBCDBqW23l85FCT6PBd+CmC6
HxcpJsRa/9lzH+/FBptCb2zcI1606xLsSoHovJcQa4ORKvKd3n2TCKNNwHhH4KphYTgjx9v1dVoC
evNaYv2jZErl+L8LOK4y60GkzAC5mlDvHwlgbJS2BKP/doyJAVJMdxIEGEfdX++AcNks5uSjY57q
gp+19XjnSM85HGPDqfFGvb3csptt+5FFinaWdlGdZV5rZfImBlvywcm8K7r492KYs2NeDa/FN8EO
KKnL8/OsgpXK6o7y3bUFAfhTVsjet55XPl65Fn+oC/gVfrtEYNlt68EnwoqZjsRJ6O61QI+1DzYr
eZWPoQwXmXCzFyWFdmGxVQbAS3gdZnZnNogdCdzzyGKy7mjKnZDMjHGiTcUaP1BV+w5ijoiXXV/q
/1dEo5sOf9+8TVHwNuSCcD4lTkV6WYtay0RD01mrzLcn53+4bMoRLkz2RBNnSsyXVPJt+HqueAQi
haL1hBwFr9dEUbFbwgKExloceQqhIDl97S17KlBNAfFNVftwKDkdeH4XNEobwkXAVojsA4cIXib8
RBq2elKFSDr8gKizfiR5wFFy0rej/HTT/pew8nYZRD5ScgBLaqF1HAH1J1TgXufEcOVRFsdVjoVm
tWuOL2rxevChkPTKH6l6DPEjzUgA1FO7XAOl7w6UMVI8LzlftIJOQLua/IzqBHhPwwozGYldxh+m
Zz92kKX5NJBFVbrgLoII4pcaf/AXBitDa8ljkknQJnPl0aqMJD2h0jSl8CqL2tS2cgJTd7Q6v+6b
CN1UeiFFEkZHNn0ZgH9xhH+slfY4wD8BKSF1/L9qcVlIv/P0A+Sgk6LvuOH4w1Aely7gW+GhZeAb
Kb73ea0nhscmam2Dd2CbBgES0TmjmMHBtLRmsKrtM3ehhA6bfLlk1P8T2Rtu+xOYCyUQ8b3ninho
yridUWApC3Y8xzBnvTCzHuTYsA7p/ohoRfkaN/0RppGVM7bwGIqC3p9GGdZoG+r9a+BMHznRiJoS
Nv8S9+zXmK+ZRmqkZGw8qfWH8H8ZVrt1PTDcDXXPXIJClEPlgoQL3nQLoVxpEee4/weCi3S6S73S
vYaI79274tOfK5RxsMMRDGDdKBSBlhLMQsQnBIOYroQBE14Gn1XwmtUKUmBpzaUqR12Dfr+AEoAd
g/TdlQDGGr4DpTZAYTPgHpsGbF1uL67fjtfiOPVeCjfwlF9EmDClEnxeA0vJ2VFjsmdMZyi9AKn9
VOjTnRD2pHkrAybm40NSjD24ffomxBZd/3hhLDTCs2K76b/4vpfFbH2gnMxdlY517jK4ixN7x2EL
llXlAL7mBVrVUBxB/cIblT8V6PX+7RniAAUivPU3fv20MU+B+UhLrrpYknjTbSv/RBGerhWjZK7I
q6w2YXpNoz5k2opN4AP4spq1qEa6N/bds3Nru88BGnYQGgkjwqZ0ohBzlezoebSfjIA4k6Cx9puU
Vgu3hVWf0N2M2knoA3eDK7F80chgW5ili3oWwiYWGBrJn2IujqpnaF8wL9YyekRzH05mn1vgIUZB
MTVKLZFtl0NASWXpBeeo1SATSbxwt5B2KGQjc2+Vzue/NuYD88+oYYlZj2Bsu8dRCEp8RjelcGHW
jCXhyrse9aekWKKYnXxiIo0Ck9XC+eC4DKtCvhUJ9ruG+9dMZNM5faeMc50Af8ku1epZSJ3RvmvP
frlxMQV/eQ+4TgqIpsQMrmB263P/rbMln8yy8HT9AmtqIZ2ywAY+QE6h09k0g6bIMue9+/mu6Hap
bKLOlC2foVEuFbjfupCnRv+Emelk8LUYZE3Z8pqqeata/0GBjzgKsic8DyJgS3nIwOEKsExVTVaE
U38/W4XGeEsycOQ1djrqpMzFiqCsQHUl5pC6nx1Q2ya2bUtA+0nk3WaD+ZXQcnsFdveeTTnoD01B
denXEGJlkLZnWZiBsAmY7Q5GjLXSGkvK6T3+W+9/PaB74ulaZtTJbH2/MqM8daP/fEaENSE3qGWm
Lldt78evyFVcH9E3mCjyJycjh5l/AvFBJek3qcDMWBB1ZJCdDQkhrR8KD1yr74eKY9Y8fwm7qAqx
eVVy+/VUgHQ77Bp9gIpS2sk33AgkuyUnB+TWrQeFPP+iLf6H9XBBp0+xyuZi/yK0S5cPOXOxIB6+
kr9wcrOZJXP1wuedQ+rMjPcMWezv6BtV3s3yL9Ui+G02TdRiCApykJbz2sowLJKgbMMHnH6/gjMO
WWegrKJ4cXK1MvWFfIAOTruW3dIjK83G/RvyCVH3Xw2vadz3/c/c1gYSZB5S8Igat6vIlvJePtKl
qYfREYCzK7ZstRbs0l88pERzv3QhBMLPHPcwig1khPyF/V7l6K/2Sf4hQvli9Z6Sf+3/FOrhhsdp
I0nBbP4wvUguAHE3A8ASUa0CP2bBhXi6TuSYUtvMxyhp+2vfvO3GBM+SLkI9/4Lot8iOEIeaC2Bh
Fry20tJnROvERX+tTJYSb9mJYEz5FObxyhREIHZJum0ej5qWOvsJHvnIwUSc97mTnQNPxoISvu6I
tQI010f6kcahjKnXV0FaVnm+LPgfjv4KNvPtLigM2toPbmBBWUkrF20R9+M2HxSsoT5Q/MulnidI
tnhFVh4zUdt1gNP6C+8ndaWdA+tR/sIQAk3Csq6DxIU8nUzxx9b2adTUDpZtB3xoflW1GQg96syW
ApzJJJExK6J8aege8Q1dcB0wyeApaO3MQtp15dcX+HNnmXv/UDkMs42+8TqVmpa3JigzIZg+MB9/
LMjc+eMUN/+NS7fCxEXFiZ/GhaD40a2WVGB8+e4U4yuCs9CXxsWdvFHKmGtoV7C2kM6KqPD0v/uP
8WMevvfSoTykDPauvPbgcecbBSi6ErQk2bI8YalVBPl55pCbmoUXrNvYlADGW+DvfKPFmaz0lUf+
qOpVbLLRBFKrHZKmehEw17BAmOnLGBIgqsC+EnO/BFfAZvMGFo+NGh1RK9SiV2HLXTRLdnB8En3T
ilcnwNIDLJ17pv6ey2lhcRHmMH5BdBDN/qx9bEMjWMkWO4WPQy6kCWR59WXXYCOHiDU8ctl5m6mQ
uQ7lmNsHD9nGYC2jKW8BZPDqv4HLXYRb2m4awCRhoi6mV6cXKtVfDfZk1F8Nh+XAfOn5V6rn100Y
dUKHhvwTy7lwQhGPdy+TIb7Yf+02LVCjHZXueHKj/9LDYK7YakxvegDbviJEDCWrDsh7tycqcHPA
MRijaOErj8R1pLg9XwhhV9SBahSppz3XsE0Z8GvGE6pVo6C1U3j9VJejOZKGvGHW7FNCqaIhXcL/
uHC3eoLPrArI+aEYdosm68+BEpqlyx226bnzB0C9+5KPRGGFdAqqUmnZKVHkOgWjukhhE1jnfUHF
EokqRKyXbuVfpVKbrktJpbe7eB29Kqwo6+6wM7WWp7T5woCafoEmf4RYlyRyNW3J0DKFGa9bd76d
LQLjfumidSXkitcyOO/8och5u6CCPRA/BI9JjbkhR6F25xRlojS1z1/eianFtdLQHu95PvlBY05R
WUiu37y9lXtB0bjwNUK6EtuyEls5CdX3o6aTPZIzUznwKpsE51lVzEA635yjocaQZfLiIbBnRUpS
2tDIo+81RgLkZjria5cdpWZvLBzTFwLPimTTEHL62J3T6i98IfPzZ6+E/6+vjLZQ7gtQzDSagx6I
f6W6rue/qRYOvDycaVKD1gAOLjxUcz7jepF7/iIfLQ2mH2N58ut8UosppulwiiTQD1NTbNwyFbnQ
9Rtx4ilmeoQj8WoOuXf8ASRdSRESDmFVF0S3NUsHdEnUUMIqJG4W9FS+hCFycxy6tBa/aTknQ7+x
caU/+44q8mDir6fTqXHfMRdXpdoWEhziOa82x6hh7Qo6daf24IF5m/fb4dRt9fZMnCEhslfuAoEN
RGkA3Qb1O7ncgty03bJbIDFBCFrL00N4GIHqfiMVfmuarmnUSydeDvQ9fLBdg4jVNOx8IHatyxD6
uNG9Z/3/RamRxW1owXEj1mrpxgyH6y7WWnyrEVC0PKKIdWTi9zc0GTNyHrr0Ntn9LxBlpa3QCbEa
k/2gPJtuzs+BZm5+XvMDF8Rt8AG6aFa98nsNIyP26fWuf7hIZbM+eDzeN6ybNBneJgaq7UJIpFp+
FnHYVuoVk1/+x/rbAGg/YusQo7lbTQdRdR+4CjmA3fFhzM7BZ8WBjRYGyhS23dflFAj+N66mKnM1
p+Tw3CD+1x0oSUWKtAD4/FRqh/Umfw5JZ87EOPm5FhTEAtjAwpuo7z00mDYSux69a7xbu0dhcxVp
3HtiXe2f6cqP+eN7IjhVWXlxzFM75tfXCytKlse0GMFR17u03l6SwhZx56GRmJYiwGAuN+uFF3ee
Ff6K3esKZspEPk5IUvsJFscr7KrKJhNOpEG+atOTEXUi9GT/HCOHLZeFBjUF2OKUofpbPEBtqNCi
9dl/nR2xJE3FXoA0k7zt82EUYXc9eQ44WarilRWgcuxKfe5ui0G7f1pbbJyUVCZt8qCV5llWkCmT
5a9wcaUkes07VT3NeN3YzJjr6okYiNxfg+5l2ui8jqZbiyk1FdJCDtUuJt2k4w9f4P+UEe+WvobT
EL/I9D/5tz+kmFjnTm0NyssoTn9zThSdIWc7jz8pBc7a+nfYmzbA0E9MH4MqOD9UXuW6VpifAyz1
BKLkxEnn+HjcgrgeGAAXiiSFPSN/lH1XPajAiilvJyjQBdXLSMhV7aJFtTVYYirx7S57nDXmdTIk
5JtRZG9x1f5kBa6yOfDWEOi+X3u16XnF1RxPW33juMfOOlXwLecKZCA2Po7KAciJZKFPNiOmJIUB
3BfhH3Ab8Kn2qR3JjBCAq/4lclxU1MgJ8DOlPiFjsNbJpOxniQSNvZhUO+Nst1o/crhkMHAm8TgX
Ol7CRoXapJKbKxQ924BJqLmoDfQ=
`protect end_protected
