`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Km2GY+ZxYdb/GRXS5YuxcGoa8WPZL+jkjSPYcbc4pS0r17jjsKrODwAA5X6X8VzfQ8Ezf19MSN7p
Yld6b3u4ww==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZcmjilRc0sHDAXHsNGXqtBscg3WjyPJIawZD+SOyLJW6pbd97JWffW8BNaf7Ngmsr8bPWCocNH0L
jIPlop3GyqO7XyanHN68HeRGp6no2mSgC7brQoXsPWutnqV/0yClvi+3AoB7NYdez7Td3USU6+7h
w89xUAeWvkw9Gp8CUIg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ohcUMzBf0n4wKn1lsaJgu8pMPGDEdABvMey1G5V10BTjTqUeYFimZdvwRGo78L5Pf2o1EWqQxQ/a
mMrm08ZenJLnDM6RW3EnNDb60OJIweAU2w4c0/i4ad5SPqz0KVzf3yDTafL+gYsX2LRiOYArS49t
05hmwFA0l7pKgThqWXiTaRNss20HJq/w32iqEG0SXDDn0tB1NwB3XfxKkQ31pRnD8pTn3M9wRM4C
I8WCNz2uQMN7hj0thJQItU5FE6ZELlzF4ciYmz7Lp75YqANfxHa7gwRAUGRuTN2cTkapsHILsPNb
+q+u9kVrf7FNHkVPsUdTdvQdvI4bL6NW8HuyxA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YGfKdB5kY20CFxCy5nGuM93c2kQLyMwua8YyiMzWcwCm8hJBFvyCqrtIq/Z1lV8ey5tInz3hnXhB
VhpHEo5LYLGeH6ykKdhy2IxyMoMJgPzqZ8tlLkfSzYQJY1BVydqRUMB0CJhUSA47CoAgFyvdtvyB
rxiu8dFcIH4uMJFynQY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Bt3v5fvHVt6RpCYxkUSuQlFLnVBgtiB+rPzl7Is1YlBoSHy6tabwN99dC2leVF7q4pe48HYIKSPj
K3TLXvLloUU45THwxQeMt62kosRzsoApRNSfClOej3DH7tr9OpT+00pqi/Twr3SUuO/mDrgwSMcF
1/l1y8i19+TaFpaH5NofcTFFUsdLQrEKo+hQORN5cL035UjsOEBBOYbb3R5t58DlW+t5yeWe4qiX
HAfRXlzK42DP0hKUtwsWKK9tOvgF+SE1thkRLm50LBJoRcnRtjEDrzgzHNtTb3ia31yYjxbfbWCY
opCeYEMrkIxCdfO/RfhFQ016XWqmNqBP5+1QdA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23344)
`protect data_block
0OkNXOdfAkU+5lQgAML3Ds/ndm2o8EcKEEuGF9GogmwRDy77YXOuiMTmixss7m2CiokIO69e8TW/
9ZTmc6Sopry4SVPGVSJIzBIgb2O6Zc6y+iEaYiNAJ9CZ06kymoQRQmrci1XYzKVZNGX/PH/cscw/
5IM7exkmhlmo0cbcBJ6+xg6KLYKKn3IOS6OVyPrUJ1HSllI1mJIqFLP5C/5BDlO++BN3TOjhhhrv
WGnN1o8Pk6fha9XNI8gjDY6iDGNdpb1GMD98A766sHHv+YFMQb3SjNJoXLktoTt4geLrgm3xTfqN
plVNCAfQBeag9FSaWTpeUO1JlC2dEebb60ZZcHeqfYWPrFazYVZssZ5R607zO0aIM3HLdXjgWDTW
fDdRztlVfIRGHd4RI+zXT2Ai+xq4MJpVRBt0etvkUqeelDpEjkMKrYqZ542aktoemtFbaH7BItbH
/oblS/BJ3Lg/2QOQZE/nevxJsyZmvDXG3jYFFvit/6grAXkGOmNI1FBaWZLL1iSTpJ1hUjUeP+Yx
JRDLQFwmBNzVkIUIwOBms829g8miHEagHS17fPW3W78CW3BGKviyRFFThjKtee5RDvUv0ProwmBU
5yzUB8uIAvQ3ZQ87uCuSUv4bNFNA19MEWdBvvA0Ds4B683a5aWRhza1CgupPSWimq5NEJnJr8IpW
K+FA/OlxGYM+R4od+ruSnZnpC8kpETHVnTW9emVQ9c5Lux4JtsWNopmTs3VUIlmPzY3CBw1e0JTz
bpTIYImsRqpOnXUTKgSbJ2rneRzFSUgzjjzPMuf5N0lU8DZ2H+agqK2Q8D6ZzeVlH1w5BjDS8ujb
XWcTa+YGaiYM/UlQFWUozcEtooI73U6Cb3BoQE4wFPRzI2tCl4XQknn4PcHusIO4x06FQH9Rrs02
q+YgueEtssNnMJWf6gQ5GSbAqHRmF0a90+XWXZqFuuSkylaE02bz4K9N+sD+N3I65OK10fuKHoUH
UBF6P6vTt5RcMqgU4CAGOq4r1/0itzqNmnwhK1Xt1TU7xAIIL+/1ETNUTGO3uKLcp/my0Q6HSnEC
JzO2Ks446NVkVrkJFl+MTMNjnhfL9nco3qvfhtLyQLaeOExYdBkjJpBnBkTXUIKLHnFuR8kxX6i6
Y1ZaQn0XxcEqgtAe/OcXWVQ5kJxkZXh9H9Tp+/bHGk02Y19Eszy+A0vN2/d9IhevW1MMb97XEqnr
qP1ANHoYsttjo3u7ldvS4sHFVCKHGZVsh2UfMY4fADla2rm7mQVexGZ4FA6NeGmEfkwxZb/WFgPt
HkHtzs5SH4QapAWR0enobn03sYbIk4q+gigjvCSPG8CHWWy2n3ls5a0odG5PNZgVVftjVhWOv68x
gkD99owXR0ee+yvsnDakiiwgK5gB+XHYLwO8Ai53nai+yljVbF3vVe5Mp30Gnl+h3l6OkmAl/GjU
vsKqEGwWi3QKraKsAqnlAD6N0IgnKi2ox8YXbwb8sAS99BmkUaVMUTIjAAR52Zhrj0vxC7Pmyfbr
XBcSglPStyOvFglCJ6leEEpS+eiXM/zdEVQz3iaCZfQpsmXFDALhDkMeCeF9Dhuo2Mvjw7dUOQm6
tvJ39qPQFZfIIcPAwk7cSov7PMN40OeqBoDSz+BX/nbojItjJy04C+kcUlR6lTXpIcVEr+uVuUHJ
HX7bDPyemzn385D1hdKt7p2JYcAlRAkbDKxalgXm/xwNSs7Gs3Lr7rltcnFRPOPBQCVdytkDXmU7
A3r2+CHRD427CjQs3JBf+mvvmi8/8xTRf4VpW56hKIlmdTKczMlu9mRIzbuibOzQP10dGcnLh7Zj
X63Z7KUAMxpd9j4YTzSPEtEfVCTfKid1UJPn5+GLbo7Jb81Dqp4kTU/300HdiqxdWhE0K5N8PLZO
oRATtNwXqx0hFqFuSqyg8OuoHT+PycdSUWGQx9WxT1+PTcA+JsBMNBBLpQ1lbMmMGTivA2vPDdTV
mvVs0KTShelhW52w5NbHMdibmE8dnqe1+jagIUGmlzVaaS0bixC5bqwFHVgYF4ZW0TOWt//oVVcu
95P4H22U9h1guM6vAKaf94BstG9mQ4xYhgqVHd0iJ4ysYxoBD+/lIVJh5rbKXEvLRufWFKjt1FaJ
oZCiGbQC6OiGvLD85GONIcE4tsFMvA4oLYJggg1XXj1G2q2kritRE5bVcwivvt4T+L2autsNqYYB
aP/fj+YSgIlN7Vd4rPudkRmURABc8TMDzNCJGDid7jRUxH1ypKHKyq4QSjVGuaGr4nucKPBrgxov
iD1pU1AJv+lByHwGBql/LjZUvxvEp2OPt56ZcvfAMJ1rAUjlfqC7Ri7R4aZ/zRC9xcm5LGnR5pIu
jxxktm2TU/l9jw7DVOYC9aJKKrJ6PssaKkdKukAL3qQfZOnRxI1o7IS1SsPcUIzfeyWlqky6aKtz
umQi/yKL6hM0j4oSM/QZUYAq1XUiokB1M5BfQo0YpjvF9jIJV7YFA2jGUS9zU1sbI5HXdWzH7/pH
Hahk8HJ0jUxKyy7U54Zlmhb+CfJaIEOkIJWEuGFUFnREgWQedZPz6L8tOSM7ODy7GQA5J0jyey2j
9u1GgU1I74aigvXqa1c7LnVFqkKLA4iqMkpkrZgV2IyooBmshNwzX5V/P2Do0CLWl+tyEZxeZdOB
F0BfKKLVAO7c9862DAmsClMdzXaNzcD5yqTmR8zWuLjjcQPAU5tj5uoe0mx+UnNbOBHe7+J8aN5M
J2uSAuvm5idUy5wn9EhWezIcvxWiFN5vYveeAQT9drUKpVYx9eakVSE5/OTgmM+J86B1KAPnVDF+
34vJHdAsAewck3X8igEc4foxdMPbDpv6iVmRvvYxHTPRqkN1GYzEaj/b0//+JI6EePi8QRhm8OPR
x0l/dqRpuPNyxYS0kl5G2qOOpDmjbaRjZIig5LgarprmIjydbA6BFFcR9+MQAQMGiSYtwwoKQAiv
vXVe6u9atFkIEYxsny34StM0jLqZ1gUeiU7TmHyn9zSpX9CB6SqXcwgkt//3UxzoejTFZuU+d9VQ
YqZJQNMJg3gNE99glJJAqGIA2ZMX/IjTVXL/RQoj1znF/cDj4eERmysVyLdtBrsyJX3N57AWdAji
V6/qorT5LOSvn6FulxKMdMHEqBmuZq1PvAwBTwr8MrZLqxcw2a2BqYmLuRBVyui33c6lwW7gHqrM
7k4n7OUNAPj8MBPpsJ5TCMrkK2uy6RiH6nfO+oGACmHhrNiBxVnoejFyjVogyyTJKDgkbT3Cjewb
WL5+hQ7oE/8RvIVu0U1WdNjh7YyTFpj23ao3nFlqcMHxkVNXYvCtneq4UN81cwGjEtj8LCdeHUqd
0CdO8wpnEDTeO+5HQjpw4OrcSTs7tlFb2v9Q12va7RPOCM0t7EHVdW931P/L45GmTi7oy+gADM6p
LbfbVVCLixQ//PeApqF1AyiZ78+WIUoMxn233fgyptpHpKwAVqVvaWeodAu4kCGz3+PQowI0iNE+
JsyUCAi3asjNedJe3M8pCyUhVRpuavoK3+8SQpVf/l0JIl83QEt6LWpC9bGdK7S8m8QPowRbabiV
mWN86t1VwZAe95jdBBn2jpPBNYNo96YBB9hI1XVJnNaUIoAGAQxoTc6hlPt3V5W7ebpk9tTsvM9E
xVBzUl/RINigtiWKaVuz/8E7jnZZsKrXWgPxKCayhOBmNIUxJ+sHdsyv7TgzP7Mi/3hcAkIzMJZL
gH/RXSJAjV5t0aw+bQnBWHWiWuEhd0IzL5b19RphZ/i/6wDrBBk6egNPq5kYz/D6I/VSnGeHNgbl
cjAvobuszs7xSDrrzQdAw1AyqqUNpxEDWpT/kzfNXtMMHpHe9hayoRAAba2CwFGbBaNBAo2G8EtY
/Px+qE2X0l8z1JOeJ9r+rUhUuk7P3IRyGNYXpyjGi82ZxXXhvCyVtyhifJOUTdHfKFgK1/hjDnWe
aEGs0ZIO0QVvUkYuj+wm2A5qrqcYgvCWt2TApfZ3l2Z6DxoIpfofq+25aYGV0mwnbsarwS2cYDZE
OImjtp6rU0M4DJuGDuIc5wyWsPyoItvAMJgtU+ox8+rPtgLIRyoVUPcxCnPutiOzL7pNruAB+b4b
ppfdDIhnwXZqVkXjTanu6weh5IpmCXVmYvINDnLxA3KrgXfvlTGSikX1kIpXX4YdHNLCTA0sXixq
kLYLOlx4BAliBUFxXsuRgqdB4k3fsLb30f7orc6vC+5Tv45EyA8/gpz8f8BPxwVO28yhwtFjUHxF
pJlmMQ3TjrIo0vWYRrSBaFuIh+ki9X8GYKPutW0USS484rNhMgbzi6D7vtLodPkKaAcylwfKyxlE
Pp6DlqhZjhfLOe7rJbSoOVa8/zOkfcpcu/K2dcLKTNa7tWSbYPh3ZgZh063ukYId+AkOkbrtBABp
cw0Awynd3jab/rBKkvFNvQIgUbihVGrZpJfQrCme7r4vRaSmyGGttXjXi6ag0qwnj+L6IZcVVd7x
I45qrIQ87r4VSGmBD4XA9/ZVK+X5CWHVM6Edwg565MWo++6LDhhAxscaxRZuC37R7i3NfytTXRHU
G2RS4vttX3IsFlI97mbU465kz3zqMX3X1+stDIcGx32ZKqEuF2XAXs6WMaTty6jqc4cnCJiTmARk
Czw6YvRHrufqFJP8vB4qev1zNkVI5+d6rpmT+TmrxK5clP50gp8tBgIln+ReJOBZAZc1ML0FQ6Fw
QG9sEL7v02uWhzWZ2y/UfvH05bL7DX+pWNGs7+hfFSRRkXzh/o8weBa0Q1r9ctFGYu1iaX3cD6sv
OTSpufqDYQM2y7XADGbgfMbwYBnN/d3eipLgFGiobccmIf5lCCGE6MBRmF1WvBprcIo/f7nW2uSy
8ORgljDwfOdhUjS0oX3OXutw57IO9DyURkys3qV7d5pB5R+U7vTHYXZDc71ivkr6DoCgMND4BUqt
btJwiLJQQmPQ9LmI1S3gzGAmmdZunOB/6W0OAL3HfKCg0OaGZiSqZLTgQEk6knoPkBX73P6cL47g
OX/9rq6nXODGUqlt4l9ZVtwvVutoVdf+vl/rbNyyve9BtUfMBmPiZawT0J6YI9PfCYBmM9+4XYSf
envlCN2B3cliMXp/y/FSujoRgeb3tJg/5KMiNRGn+Edm213391k6mbyXrZUudFfKM9xkdyRGS2ZA
qVfOd8SPS0qYwB1hkXFueNywID/Ke53L7TNCbxRVOHtVVE1UJ3xkmOt/qJv42ktUVmFbza+5k6eT
LbMsXjyqg9GAfU7ZFbIHrdRR0xYcmCvTN25RL2HOJFOshm0hPcAxl2CHBfZyH66iHJLHDDuvZ/AK
uEA8C+Dbe2iqY3ysZYMEJJ2DyMRo422zaAhek9TLvgNhCvop+RXoN4LJyobkWfZnhTh9BMW707VE
S/u+wYLGuEtwaVxhZXYSHML/L/BINMMiBnTWgk9TR9vQRuXh/Zmg/nJwv6+rEr9s8Sn2Lcndh0T0
UsvC2lrwq5dcwvOnYjb5tuLKw9vUCBEnHIg2IzX6TYr4KDDCRHAko6+nvwdGIRQ8rbA6z+ENlttx
nqEJ1kVVa5R7SASVhLfCbog6cjU3A2hMkqIIAebxMO1AvxlPK5IUi8XuH7PpTGjSbzEPmq4hg6LQ
WO9AwXvIydC8TZZMsChIJzJKjDR//QLcgDcSz/3YRj2XD1qLq2b6zzcMynfUnlwbp0YWJCEVfUxx
FIdeSg7xO3ONkZ8O8S/0CPkgXyXjOUR8vTCl77wlRFAelLgaIJnZf7eZEKI/7C3meFAyjOizhs+p
3VgNRQD1v4PuF9fDPwVc0JK8vtcq0f7Q91LfuQ3d5TjMQLpC5t8zZHVwRGcUlTBGOJnlIc/Rj118
qFYtRM/6P8+Yvdo5BxEOll0UIyJahFb6niKeFn3m5Fv+tpSA05APKLnhFEP42UtvCObLBVq3DtpE
j4L0YwTtutOtDUu+BQD1HYvW28DbzQVQER7+It3vPu+m+gEq2Q7UUvW5pZe01km6RYi1jMkG7J6R
j9dBkjIdJ3h07FvGPO6EoTSuAPek+uYfgkvu0FtLS13pK/Ik5UAJsRW0TztPejkp1ZT6r/Gm4FqN
yzA8rMStccRHWF+YAbUO6b3VFVTc3Az5SrdX+C3wdc5UlHDMfy2F82EQe2GEZX45UqKjwLh6hs+t
Cq+UzjudKWoZf8A3u1tMVNsdmpCHtVq0epn5mAfIqdDh6QlF1GMcUgKkdvBfC+GpYYCeRCvZW2bu
k0Tfk4JXYIXhBEmw0qkZttPweUNkvJF6q7sDCCDTTNF3DZQuYT97RUlwX7HmxfP+CUrQwEm1R+rt
zbudrojHBH0Q1T07HtT6InnarjUlbsyziCbPebbvsQNDJcDAVuiA8cSa6/wWGr+PnL6koY/cUmG3
LA/YHGEvENg6h4cRtIUtt9K3ozh4QKHQQ5KrJP7qIfTpuzunJdm9lYo4c9lS8ODaOZEwWRswsguh
j8Gf6uvUz+ht8rXIjVSqVVw/cbKHUI5VZN/ike9Y3LVrFlu5MECY0hyJzvehyNsxUjj59FHCo8VY
XzFe8B6yKqSmIqoIJmJF9iMcwVtpwho3BxWQVhhPexHD+R56UbKLba3VqFrmeTJHfTpkunT7ZzEL
2Alcj4KT2JRGmyV1C7WgOK/Ouj4YRZgBNkNxUy3hWQVYMdo6O4PnDP2OdvkuLzMin/pMPcvQGi9l
06aZzPQnWte6/Puj/r3JfLp05Fbvg51Q6JWtizK5Ji2QLh9RK8PSGZNXrskZ8fd/tycHcfyclDZl
QXE9RgEXNm4Y13nBTT2H1I1KBFoPhQnez2+Iu/oxzsKHhau8hQ3FYXNF9VMMa3JrRv4r06tEWhbr
HemxX1SOSsNizj6s310deUbpEThg1sunBfR5NAkfOC1wrXCXDCugqvFL0xKYksIyST1rkC03AKG8
yEMs46+PL0Jx7UBIqIlqXFNkeOjNVn88PN5Sf1bq4UzKiN3arHIIjzKbQGaQ/zcFM73ISuGtNf06
5rW4RJiD/x4xNPvfCld+pohJt3HsQemr56+F3e5PvJlA2Yff4fEX3hqml+XZF/OQ3pe1KI2VapsH
ImH2S1iEwne3M4sp2IZwwU2RHl3sYwxpahGUp78H9808cYgn+GaeZ2hbfBm7eOaFD/LPTO88G7F6
KdW/Dz8dwgrMvTBjURsDXWpiYBz4cUl0igrsZxYweitqg/WDAMbxBJAp4nx7q72whei0+UwU775v
nCIYngpTRBojpagc1nRgjYmFWVC3lzhFSTgya3nI0Y2RgktURAY2vKIA1Qt1p6CsdNsQvJb7QQ9E
5RMR6NIHbI6yR4+I1NOVkRky/f9uaOe9Ts87UMFK9tzjcoHPUh/nBlmRNyJnFAQOojq7xduEnU4C
hfYAJyRDn5jdUtvxGe3blQXRwsBx9aouQmhuiG5K0QfMp9xEC5beglBD2Q5jIbNN8g1J+jrGRCBL
Rk4OCFAUvtSUSR4FPw9Qe9CfBgJoGMbJeV0QXwQaC+k6SY4CtoHvUKIJHUhaecBK/9xCwSQuTcZH
1K0q5W5gORnZWkk4A1O8l3bAhjlDWXVxOoicfYOASnwqzsuHjlz8cK93o/wseQl7hEBgixwM75cK
lw8TKSX68jid8EX3gLMk4igoISwa5rdm+UsQq/bhxHWdaYOEGQjP9dh1J8LSFlw0+qBMu2xiu8Z6
8qy+la0+p4GKWawFhtkRDWKY8uuwnI+mir3JF/JhjHgQnvQTiiudX1AoIJBjlJIX+/rVm6b+zMxA
9oTDPOt0LH/TVnXOvBnT2aZyAibqsA5RKlGF0GMXWJhoDnMph6cznLwZZ6LOyOnMnlxuj/2JjjJ3
2PkbV56C1hg5Z8dg+4vkHZt0CeBptrTqJMzCZEezvsFtrEtuv/gYW5v7Q1B0Rtlm33YeMF4FK6zS
1vfQ+WctnEDInxArNAwkIqTLrDWRpA255rSMsrvVU64Yi3POVXsdPvkCBZrIlH3gwOp/AoryzB7R
58QHg6pnRSxxAe74ElAqbiLanP97lEXw/XWRfbpD0takYqUR+aLBRfCClCn8/z3yyYYW5AxCr2gw
pwjLZTu4bdLHCPL7H1xLRpWRwQtw1n+VbxorwAFhKRhFeCOcDtjwwLXqQ5FBN8qBMlcTWf7oXvPe
qy9MtUfIBs5Lke0c9m0/hUIm3a/+lfiQrNMeQdZ4f/Ir8+EQpXSopjI38UHleoFClLzkIf8eD6bM
Uoga1j0+N46xy8vh+7xUdXmS+96cHIU8ab+ZXEkUZqaSx9bz57W9HFe0IBR9AtypcNFrn+vn7QLN
3v8uwK9vZVDK+sBsYqNdZ9c25CC2WW5CpQ4AXQfIsA8QvwERMA4pn4J2lZ2MJmCZJ1DCE7oF/aUb
igfc+qMp2PoJc29omfnSs920ygK1mw5QHqBfMu2NOoYWY56Mkyi1eaJVgjgfDmazVSC9KNvbYN3Y
kB3sMfepbOE/9JFC07R9jzOjxFtWC/Iusg3zvIDJpQxRiwjEd7UH4rdZqzoehnMhi55i9OnqNK2q
XQ9k5hr5vV8ToVXeUtiKf8WMaNqxkZRBbt5/6QqICKRMolQfQokPJyiM57TAcUI9SzkeTYM2O5fS
A8Kod3EaNpU20MwBFo9jfOITEs8PgWFzilHdSHP+kjeYHNYOQheqwM2LSrJJDOVCtLICGvF1eCq0
JKXOFfTDOE+qoBjXEKUr3uVFmcAXUprAzDPzsYdiREljmpBc8LNXNC2RKcSdpj4bBucya9+cBcXG
gTB9YHABKOlaEvCzdtuogiPu6ZI+ftYZVjItIq3RGgh3hD+V42PRbQ1LtsErCkqanwxjcehn0vQO
Qbjifqkty/51iuBIiWjcJgJm0Kdm/qVfDWNDrLzcK61JwAxXaCfEPs2iKnwmMwCTcTEqC7LUhjtU
7yorfKskrFORk0zZOTvyOoh//ooIZVrcsfKGGWPqMOKTABg8G7bOHyeYbVFfl6NDy+HvsLAskyia
EtHpF0rgbMWb593ipId1M/rm++3ME3GnYEpd3BEPN5g/XVy3alxyU1+Qf5uEuPoiF9EueDFJhSdK
SnjeIyQ+uy58kYCB4Tmuy0sd4rgx3XSvLV5AR25g2kJvGvEg7Uu1hjrwOtZvDbNTA8YZ2/JhTtkW
AWaj2N4bXb9kk0fRgnc4HHDukGqGHJm+cw2O2yjbQlFxKVABH4NIA2AueCyKrofz1UI3e3dYBzod
d2rRJmvA46Kxk2XyWS/i1aYVCKC86zMNgQohtS79d0v0oiFEZIzsBUzpBcXcSd2Ss8pyu5pJrtar
t6hqGDcYlGxLUa2obLFmvg6q2wbjdLOgH+yqW2BzpWzuhaQWooaaIZjKwjn0CQt4asmRnmKumgLE
rSPVybg603qw7Jb4lvXx1FPPHcSDeRi2leRS0f0mWcobvVksJ917RzL6ri//82q3OD6e2KZwoDcS
WctPeJJ4t33WDRviXxiYsE++9Lr//1Djh/f+D7iTAPpNUSDoxGtmJivNqpO1ht7mnfN8xT08pkc9
eSrsE85rmLoSqXGldeCmPA81P0X1XYEwzoTvSLIDTG88kXhVOby6hjjuAks6w6+IyODd9qX5+NYm
vER58zaOpFfmSUTcjxmTcYF2//MJ8VvW+z6M2KDLLT7XRBkSPKiMYHFzGOcmVIABx97aeSaftuRR
3waT2PH0rZCQI9UXKSFUhjgbvIXdFUY45TDHNn+md2yNBeJ2Rghp8Il4h7qqFQ1+5TXTF0OY15o6
w/1uoygkGiJF7TfkjdTLkqx8Y5PtMp9Ysl/87x1ER+PkkQFjs/rfOnO7SJUVOb3ojL8bKIAPnUvb
sAt4ldxkDt2UN8GSz5/G5H8qnPQTerTllNGerVPX8TLM8xCdMZ8AQ4lZu54YZhWSFKLc8JpwtSwM
dJ7gk7pHhVyp06/t2eCXRoapGMYsoEd3Nqri7Jvq2o2NgJjNYoNSM6ezcpyyhNUK02upYDLl4Per
ZGViaq2rfy+c2IJzwK33VCDe8Nk6q9thu50bC+yNk6QW/1umma1/fbCna8cy0Ur/ez/GAHckqgiR
3+bGjCjJj6AE+iTiFc9dC+bGJCgwVv5qqrVor4DNh/Mrc32GLyX9DJqygAu2jLhrAQJh2LoMnV97
hJaGLtfZr15WGHz9cAgdpDTj1X8mePVFwCPXvZymCirMb7PgAc9pNDyknQQ+LCMex0nEkI936ug1
/+HWPX92/MySPhARKS90ciV7I4MH4mxHJ9b3+y6PZnbJFKtY17NN1v/R3aYYQOtbr7dcg2nMvKbV
eE2RnuqpSokP48CldZH69hrU1S79yfc2M139Bz/Dqq2EiXLpJvHYBGDd7EHORzOos1SHkaHm86qB
khNKY7z9/S1ZP1mg9cGG/ONqTyPYHzE6gqqR1wLM2g8IMZZD5VdaYyTS+fKXgoNTGu2VJthKTq22
OKPINRCVzYUooTlgzAcduZsPUeUkun3vQPSngQFVWWSSqPuaHiwacssuLkYO1XvHuRt4ay1XvLPd
pgEcafcTLNcGELURqCIvBjvlmUbOlOyY9/bIl7wFM6HYAZJigcWXs/gkdUzhYcjD8iEhANlytD1I
iRm4AndctTmY9e831dccSfVGCcqD4F7mavIZ/eSYpIhjTlXEJeby6OAtLfUOhlec/dk0RP/zgMTn
RYqztXyYxvCHUQLWBBoG1ok/Bxz8vLnA6dFtcz35Be5FtnDLV6CE2GwZ0Q40p16ULVBF2PgDVedD
6DehsfKb4KioJrwezO9gD5eCgiFt1WTvFsYB8IvTzZgNC21iQoEOFmvUQgls2Ljgl1ppkDRtlsUy
CUidpE5hWrz01zhQ0beLLNXpei8Dzb0K0oM7ak+5s4ftxD0Y4Ehq0ZTJOGCg6tgL0PE7R1a6Ft52
qVAJjYmQd39GglvYVa0m8BTLppwnyRUujch7aTFyky/IK6XkSZihwNlsG4c5I2mqLZj9b/h5of0n
S7Uu69HGeOaYljys7Su0ZMPeUCXDaVKOxTWUrb55CzWjV/zNzXFga8AhL+nF4om6GPjNB+Rl30Aw
cVwXy/ghkuUG75vYVt8cdIZmNBJoO65Ft4PZhz9lHZLBD6LPViPNgC8vr4zRbvVSOteLOcgKOuZF
ehLEG95/mZ4pZUgIPUSFb9yvxc2fYCdJEmZdT8u4S0BSN2hWpXVGUGqU9fcin1MY9nEaA/UYsgNL
M2oJxaYGdEDZfp+mcmKScR7psGOElhvFq6QIvzaeAByzY3/Z4rsmJR+LHZgY+Fk+e8oLgrp7CJD7
FiCrSusZlOH5ZlBC5w2RKD/DUsvzbOvAq+Y537sfZ3uYpGTR4y7Hp4SDrsywkDdXPzUdxE8WgpN6
m4pHRgOGcZuz1/4Tc5V9h083amQmartS07XSmFnM9s9bKiWGar8uEqDoR++Brw7lE7u/gACtTEmP
8U3VggST9jglvdcSjg17YvQ6GbETFkcEu+KMVE24dxU2kPCO4G8vw3MMyQna+NvboleVa/yQ/754
JfyBlQFsjr3qWUtQ08XxInFOjVP3lfxyobFBVbXW9R6oTwWXkdTKpiU3YOQaTlxEN4KfF872zn54
OcxN8dFc5cSEQjaFzPdQJL29iPznQWoFdnWRa7AyE51tcwAHMKatP7ne/+D7ehcif+qNSPJilFMQ
IdOkJ/+Pg2bD7Au3ybD8pDN20uz8JlozkbHAKU2Sz91zuFIlU2jJgB8pOrxX/u9POs3ea3ZfWcIA
mz5zlJ8iZV8aAlhay3x4+Jat4aLpLAzhnioIFfnXezF7wQQZRSJNeld4MO8CeXfe1Fk9UhncUht3
idjoJ56mk31HH7EpGLUOA+aZ3VnY5YtmyYXNrieZj68vG5Afvd7ucij/I4iXEtNIKg0/kelo7bDA
gGZXOKCHkgfKSOVtLuTox/aTYV1z0ZNXpGODRtBsMI97eI42sBLlswDeGD05BfS4MJV27a4vG5lp
JXhNePIuqFe44kkamqHsaRlNP2uvtRlnH0Cl46yOQ9G9HaVNx6BNxCSaWmEzbqxy842OB811Y3f6
777BWNhhdWDTa5Dv/Qje4I9mBhfW1TBajqKyrYgwLHiJFvyMG1qTP/RGCKEkZfRGARxFqmea+Phw
Z+telDieRxjT0qjoAxOEmq+++uFzEwC0U14FI1PlIRl0zVgQR26mrHpGkbCV3FNjcjaSD3RGy1Vs
Jyig8cAiBiifVehq6CNzOQuP+Huno4ecmDYC7S7X3rFMVglwF1gi8hSf+PzTaN2w2wmrhZjH7pQa
z1amxqgXW83dcdJoDRV+V/QwgCuCL5tBsmZEP78fa7ABaN0O4/TqiLLzPU1DXnkqUnyRYcze0yD/
MQu2oXSgDDKHp2QKz+w9RjwJbSIPHyv4INdbUDFDOJZ2BxmMbP+RMIU5TQbf13mfam//I6vdp8Gb
g25YZhOP4+68dlv/zGlr64Zn3kfM6h9YtZwgLUyhK26k55f9Mx4m59uwOtQ+kW13u0jv8WMcV6y+
zwILCAyKbsI0okNi21+5zEqlEMCU8KTKaAT3nr4uOAqrRpjJ0RXbW7/Mr5Z/SM+VQR45DzDvPj30
4KQdV1MPCZmnmV3Sb4jUZp5nii/+3hJMLeHIeId5VMrB4GvRRX59DY0vNJBSQ5VgZfOkXT8N8blb
kLcaFZV90tWo4GxdjgalR97BgArMhQXobUlgecXCNP++ZJ60ow40QKa4Lc8k7JO3/6snyr/qMjzA
RCdVDyeYNxnkOwGoyMlD65oxKLRg2Cw0Y+qtPI/vF+zJY37U3VV1q3gPgU8CstULeoUmLBJH1pBf
/rbaShK6DKtw4Anq4+/QmqH7Z6BAbJdYIjiFKhvnSbegzO+JqbSM96biu1Sdp25N6THYEFRKkhcf
rGOOxkbepLhQx95oDTOtwGbkFKHLmUoDG/gyccXvg0TYQeU3g46iy1KhVyOivCtgemEYesZ0rZip
HEtHJVK6h/O2kHR6+75MKltXAtLSqV0+jozieSJuNk1QrnWMTKwyySXBPXH95ASwic2ISVI5QKBG
8o9eNarxwKNPli16XZfNyvrHLuY4tGcd8q1Java5kVEt0UvmdfM/gBrRXyEf7XCEQfUuK/GBY/WT
8wO4b7XcPhRzCjTd9zWa2ysk1elJxFu6/ceAgUvYvOmL8Z9v9D7UUWy3tAC8Xnt36208FcoAivh6
TmLEWkRT5QJUAlYkTMcISKP3ngiVu7Ls0CiKBiDhPHxk9EsoJnGjtPySXiTUpW13oiptz6O2eij2
iwnHAB7OOdjm0l9KQZ5iziZaOjzIKzKU4pk/yU2AStYnxPKieZ2wdQZce/tBFtpgdzDoWUmg4yE6
hxoKG3n7B2NJlLiX9oMRNpfWUMtc7/y/PJV9lGpI7wvo6ab37IwNJ5n8Q9s8LX39HYMyYptZhFAG
QWMaxf7f9yrLXTH2/xRATvhBeN6NjPx17CZqwXlMkuEC6TnEMWosi8vByFnyKzJ9G435pXmMhtHq
LwWty8nWrhAdIHFE9mrizIBvdLC1LUycTEdyjwzAK1KSwXAJ/dPy3sye7WtiI3Fd95qqVh82Egsr
DPIqcTbhbhPoy5f9E1KYjpBpBEEX8upKipyQ4CTFs7QLVLBOgVC6QzTkQWoGk0fs7rhMofMTNluI
ePBzpay6FeReVfPLPqQIDBgMfa0NveLN6e9rX7jl7IKd1VRDUETtvAA1tyXE5T/YVIsJom+MJ4QR
LnrKyv5p7pR7Wkl7tj5CSVro7FWxrrpPdrtukXM7+dl82YSzOnJq3UvsxA0l/yYuvqtZFK5veVI8
Q5A1siJYqbUWSSXqLg+t3mLqMwgdUq3jbkG7IL6K5eFbZVk8hujH4Qefm2kNUr9dLZZvWBsh8mfK
9LS0QvP1236XlpxkqPLMZfJ8Ou7xK1n7WPV/HBbRE2ikGjm7XG+8JNjyQNyPkb2ULnYfvdsbBMi4
pN0dZqFKrcDeVoh8pg2PB7ggkWgM/mVu4+kXLB2TFPuVRqW6Ux7qFRpb5IIkZxAdqGuUq/Eiq6X0
N4A7s3biX+J4OcQNqoUFlhzmsN/wyXd9O9J/o/ItUJ2C88z4KTBeBy5WCZCMgKNMyohlFrXiJu9e
ywciywDhTLldGZ00zRXf62kSnEnLujMnq7Iw8Nn05DgAEQNYMOnnSEdZN9velctGVutIEbrk3fSv
fGPDrp9qNQod2Ed9gbW1zlpkMDskZlKgqsmh+q7oIF+Y+8LycvhDzOO6biD5cAmDllRJQ69nIEhX
mfE/KLj1rqhlgZwcHlDXb1dOBbjmZ1v6E5w6Sdar4RrJgs/5X6BK4hq9TIcLIKK5ECyMLB20zEVE
IMhb+46IShXH35LI2aUMzW8i6BY5Kc8DCwk7wv3PJoq68gNUfwT6Duamh2Mqr49TYxFUXS2q0mTb
N1AzXIVjoRNZFIEx6OcL1XffWf7S9JOAp93xc/rUyODsCOlxTLUOu9WvQ9Wu015ahAbm95Wb/wen
HCsrTgRAlAUApN6xEXcN8cROAteKbsFMDEUQBhV0+SA19E7yqpkluVqRvwcKlzUa68GFVP49N3vx
U54M0u+6GoSBFLmlCUu+mEo6l7sYGp9I5vxK4F0iahBJ+laiZxMJlRb75X+hcgJjPUUehD5Cx8F0
3Ot+XpGi9AfyWgwtB9yR7rcsHjqyhGMJB5OU6vAgIZxp0RihyziE/poZltJ/q6WU0PApmIDjQdVo
yKjSaqWH8QMXLEldH1PACkpL8ppxZ25xUzp1fsg2V3ZRkKIN7Tb/GUYPAB9b091NpiCb83ZWdS5z
n2b0YaC/14X0w5fx+mBP0Y87W8UzqBvOoEczFmG2aPgFGGfpNp2wvi4sUAXbQcVJuXb9DenmLB/x
66+7M9MTgbT6pjPqCzLQtwD1F6szaFqYIFlWoOFfeeoUL/GTvt4zRZKBtDwzLqOL0jwt0BHr8hE4
s+zVsJGfk50cMF2+EU362w/cseV8zcAQz13gNtfv53GogjrVREwN9X584KAYC2bZ8ETC6ApDcC01
4AQeQBLkmDUbbZOzxEwW8WCe4Hw57IJpepaiMn3Qnstr187XP01WqGgSjecNzTHoo3HZP3/ioVt8
x73f/DJ9BgIeutsIwa5yO5ErSqJIMIW3vKsaR+vZCRCZjD0E6ulwqbAyhpFQFYxXQJeIUqTamdiO
vj12L8DclCA6kRz4CsZbRVD0psCKqwc1G8QuE9aaPwEkWzdzyR93i3OHRVpompuXZDito5hhf6kj
5GKJMWyFRQhQYqRZRYUdJL3PX/FQw2w2ZBf1nkjVgSegvhaKSGL+3DVh8cych7sp3l4RVoxSPseS
UTVEcGuNFeoTkz0VmJ8eNV0nKvCRkYnbXIaJTj4FeO7vBaOvQ5MP5uDIYCyp0xLtsfH1ph2QQL0p
t2bq6S/ZqyziQZvbBevK+u4WASD/BjyauAOrmKLrt4MRFvZ5a/8es72w5PA8JCCymLkYqrFQIZ8g
uxltBc+89NJCBzb1zOmb88y2CASr4VmfrneRDrab+5o9ITiHYmQePPJ7Sx20xQETMWn2dawKPI7M
3WiQX66WO6pajTC884RS8YrlH2fnWzTDFAHFgPpQMTqShI3e0qGgHhcFWZznQX1MVmStz7EWaTZU
vV7/hR7s7V24YlB23/4tsRJgMSgKKMn8gsf0ayOjprN1D+NPHiJf2W6Q0XPMnOfTrzkdIf5oAfY2
8L6o/XgiVrdYcYbH4sTx3t+ntg2F1V8nFfD4oIklZ1aMmGsFnhfcK8wLPv6BIgbbWla2+naZPDz7
sRRw0CusebjidG4Vw7dDi6cvdtKUFWsfSSWnOYmHV3NRNiRDCO+dz/FuDyWdpRHZBUi93KD1cces
MhMsE4jWKIFUrk+ac1JnF0mjPPu7eBTy2qo7EQz4Ca7Sm62HC0HjJQGhkioPEd42C/u18lcMYP7Z
tlWpZm930r0Daoz2emBQFE2wqPMRUmElUwZekfMvZH32v1KrmohUdP58bp4ZFwYMkv6Movz+j8Gt
F6p9iKNenUX1n283nvVxXrgN0ZdepiVle24c4E522Sn14ciS+fjZT9RYqB8P9LHf0wjPTN4HY1Kz
22s7rPk+FFsZID/UqiSB9h21XAZOf/IZr+IXfH94WVY/Uts53zMVqtcatVd8bhTJM7R3dnvNhviy
bkXlPdzDSveZ8tBeQBWxai7+4+tLroamq0G9EC/oXi+jnpw0LhFqVxHOaj+isMnn9LCLmIigX6Xs
hfZ89nAo9F9c2Z/NdpWwHB0G/TeAuUVyCjnEYnDd1nNMhREvCD5AINGfjdnSyy/RYEDkdU/k5egS
vP/E8bVf45xHVZANpMCHpqBAuGft05FDxkZxUO1a0E/U7hFHSdxMW6o2+F9SOknS1s1+v0ojcttb
nqZzbZisVD8Ch+PobJCW7fX58pyWaT4HjaQCN9PZU3G4DA+z9nBr9FQqC9ROZ1rikoCPdWc37y33
OqWqCgWruxaFucYVZlGOs2Sn1tzDdY85GjLQ1m4n9h58mLkq+wxKOEHDZITGmvsRO0Ovw0VK2Ar8
WWn2++owrNKOONypXiHv2acVe7DGyBX6BcOsn+vsj1QQyOdfVZx7ULA6nKl+RJenD5ms3dVoRMYR
xNlIpAWoewG2g9NoNQQCyNRJiPmKR9myP2ZRpKyU1ZC/aAuYaUcCHtOvq/wJGrKFkgKF5ByyJoo2
INLtV+8Z20oRig0ftjcexyVshKvI72t0OGy4bBkhuS46TVBxy2bV4gwWpcWpv9KrenEJ8iObrZEp
QMPPDz0i3Ji9NdQZmrWfvdWqu2eEjBgH+NiPVllO60Tj26SgPpQQVC0dwv7EPqpbgXmsPIvd3LY4
iB6zPABQK9fzKCjuVUnPmm9ZcnXDa/eoLoai+mTIZNPkm9F2bbdoMtq0fJT15os9wKTwrXw8kNIJ
bI1HcCU5fHnR+LnFSotih+ZHd+qUjvlqjTpnMjHCuYN6ejz+KNOgrtEiHXZghB/yhyBh3CsiEH+n
pfKt8mCYXuXqubNhHQYmYc1TTOCR7Fr9OSXBcHKTNwqC8ZCmPG1gO+wb5I8oTO9lJkPNAvCyo6xO
gr4m+PCWCitMiRvLDVLAWNCZleuBDD7wuNh+KrhIIyEzBZKFHt7K2ZXqUPleIJZFvd6JA/W73zZR
Czm/D40YdVfO+b4ay4V5dhPopEbL94SuMAfLrHwh6eD58QtTbreRjOo/ZbtuW1IoG4Cn8oUiKBf0
Pbk9dGXgLQf67mqUB7631/lvwbiwHhtGjDqqTCWdGOTVEsM9zwLbpdfOOSfmfuwMQcyI5b8oksIp
d7q42wqnrJiLTm9maghBlddGY4tW/wwF+LVNwo8H2N41W5LUb9bjON9GtiSxeZU6LS3N0lhTaEuU
QrxMW7na6uUzPB+LJryBpVAqKqmBSSyM9qykK8Qq88KqOwJ2a11iCgFdNi/autby+mZagsaZls7t
NwtFQ+oZmql4b95O/p7Mcj+1Ky21Fh71ZV4CZUdfvzlHpXDTroPlqDQlQFw4xu7PjGi0LsVTaL0W
XunDYEiwI5A7UytTokDEQbWgZyXEVbM+R/8deYvHf1RsoMAhgpRljah9T2dRXSc07oH8jTYRN15e
z8juvjq7u6BLjv+lX7GBaDI5+peQCGxTFdPyo+mE6NrqcamiFy+JXNAvz0ky9vLxGX6cETHlrRdm
YJoyBN4gwWarJQttBQCZuj0Ag78JvijAvdQgL+uY6sYQal8z5oCYdTwkzKmE+4Dq11weB34jPHiX
uzY0kmQ4M2AY49BCxDvioHStLEtcPjNgzlVB25RSNSwpZ9vouOZNW6StqJTzhVhoG2ioCqR51z9J
QGac1Uj96ikohnd+rka8UCMZlcrwOQ1f8g/+jKxXDtJK/HkV3AnKidVenECa26IJcxlq6NJacQxd
G8znojhL8Lm2/ZUyIqWVALsWVAamcXvB8Gatgiw6f52m3+LL3oe61wIE1ZDhsDRIeJmmNfDIji/S
Z370SEcJIQBu7XtTnXccpETJ0ZWbyvlq3zkFzdM2afb8vuE9p8QFS+A6gPnJXpJr+JCujTFB80Mx
3B9g9P57dkq5qsTBV9smDPoiv5/jc8y8hdv6YX1DT17r+5B/FxgMdoGbiq4uQuex3jx8p5NSI4nm
Ga/vnQd58v8ppKrQ0mVbifndULuhvBEUla1ivQfObp8xDoiibaXSBA0GgIAjwbV+QGI9G3DDP4lP
q1M2AhAXxzmer2lwIw0TikD8VC49gzI0t7yA7Ex43KB3mMCDtmpbEEtsZ2fIK+E5pOp/cPJrnrkj
062Mpq9v+TCAih5BSyITRyPE+lC6hMtQp+hzDBueVa4zvFRdQocWDbtXVFBm6jp1OdBHbQks+AWw
xaAxP4EQx5Js6iAh7jzUcBlwQgKBMZNHIYZAYi9dClrRBTh96ZfXUokPkVE9XGrpsrylhPMPDO2R
KyC3xvexw9Rv0m5gpwmHJvdmbleqWb7tGC7dwq8npVQNNU/s5W+d8j55/c39yjd3xlP5p/IEO5+m
9PX8jFu6VX0W9x+zx/SjIZizAvnSNd62qcMiEQppqtrI43Mg3cDDPdaUx2qxgF5wz8ti7vmoHDYx
rcxR4IFp1Hnm0je3MUQTDpHW8eV0zXWcHq/1cBTp7EaVqgqg8aWm8u8XMf9rgj3McQwzVMoHlsYj
Ysa+KNhStsOePqiuiYPfNPozG9RWBOwKS4LJP0B93ZnWfeJCkRaxrNQqkceuDeH35XSk/Yek4mvP
k6PNwxXZ3rb2aPqrzfV3qOR9HZNSJWCI6P2ThENMXtfCANq1kC3TqyJxhx7+Dao25WJhJgYnveuG
npXiw2KVmpY34eFU0ftvr4xFl+MJjVYkOyxnVE6R2hjHTGf4jnAtl+qIKWXTCzbJqjskTyKWBD+V
XsDYGl9dqBt1Yq/nIj7GQAHXczFyRzlZjduNgAGItuJQwvrpfSRMgoOdTjTPIZUh4taeDJjajMeD
18lMzvrXmozxGCH6OYpHRSe3iHncGofv3q/vXUE3Bxk36TlU5CjRVyTLH/JeqzeMpjDgmHLMTQaa
Ma8j8rtRzAPjNvNxzdrx00XCklSQnmAPy1TYXnTm0hFy5rLwcd6veZTh4uSv+kaSKvkfsPYrbkMO
kVX40/QJB1q38pao2B2ANgnCmlR7AltPiZwtAnCazd2VOv7EeH62XpM9Nac+FJHfNFTcfa4TK8xF
04/WY1PtIiGLc20qsLKrdgw7VNnNkmgCHlDf1KsHBh7iZzuOSiatHfn5TP+kqwkI8frizpNeDfnE
e2JxAW6bv+pf/3OnGrGaMsG6EXCMek/CRLzkz7jkgY3++PTH23yrMUCcMQMBAIzlTAts1xGon3Hi
snU9Sr9qyQSX7CaZdyYFG3+LgVVVC7K7v5X1dUcJKS5ylSiXxCXLi7cXwA0vBQNtB4kVCFSZFEvy
Y5fLkPmVOwPmjOAe1P3Va48MfOsYbw+lClNPxyQf4pkzFiJYmiWPOajOG5BdBlWU8wmlzSIBBZEt
7kCa8BLPDque78NHyZiwZ5T4MtZNo0IsZrBAuYkpmZZrS1fmxRcd2GxveJkntRXaDgh8avLqOcW4
XYCLkKF3nl2YTFxmso1kuEsZkPjobO7FUUL5ZfY1IuREdyfqTLEexWxaLCCuYcM151h+mUC802ih
SUidiJXDnOHw9Y5mRuHXajuxvTrxG5Cabtcxd++Bof0GAYqLyliqXcm3BSoxqvfFsriwNmoQiN9O
fZrn4MNsp3CiebOH7kkgUwQtAYSvlt+g3iTgdlLJAMlAcbH73c1rI1SinnrqA+XP3R8zUAfe4dA6
Bz9TISiL7+p9H7n+gTxaUeZJKWvRvujt09ixQ6aBfmv9hkmg99TuVqzlZ5VenV3bC0YzJ2qqzQxm
eUv4EtNetCNCJpwzvAHJOKl84fVCd0ZVLI2DRqnx+qj5C+TFomZrnvfFkCB+HaRnSmD9OZYBXOcl
wpZhFDB4e5lZMvPAW+/EtDv1BqIL0jfR3HyXou2LeVlimZXskMBr23r/2dQ36+vrpH9pW9YibppJ
/sybnaXwzu4gFLq1lFBCE4dqs5nc+mk8xB1xWmzKKqXe9Hj/fBKodPnR6+aKTCdD9aWUZOvCcaJS
aMBp596FuUc90TfhIchutSDW9OiOdg7fooq4V4NIfKFVdpN84fgSbUFops57CeIa/zkGytKj2t05
cmccqeyzxkiEjSsAYFgoWdbnLkCzGkiMj7bQVhitzFt/outbfdKIChlNrXIRTR4snE5k3psLYYrV
oRFMiJ/1ZhfL5hd2ntNBR+4qot+ek1iLWsWPICaGzRNdDh/cwFKwaylKv0NLvuijGDHbL+Y2PSvx
g48XQ02aBD0UZJYRqj6aac5MJaeDLMMeLELqLHD2a1b6dnVAxfucEqGxdcXDocJpH23QKS7Wik6o
KuzsD+E6Y9sN25fLzUJaokbrbqA4YzIZWTRAAQ1tdOEwkPmP8ypSjQIstC8N38ff+zIGE0YBxDZg
08jz7jg56YuXZSmXDLI3/HOLBHGu1XYdkYAPxwaLRW6BG1v6i4FsRiim/Y9Ye6aa5keH8nvrNxqI
O3sUwBEhbHGY0NI5bJpyKyr1g04Bkv7Vvw/DyBXtf2u8+7sWLNoR6lOIQl1fEnAhlMzCyr2BLIYO
BD41I/lfo6yyRb+bg/ys6hQC83SgVtZhDuJmimh5fCV0Yk1KUdnrbJKdFCwtCugohZECngTAk5wR
aP2o9flNrMQx705GF8VQ3dU4WKVLpJV3twOK6L20H/fL5zpyqkd12pZxX+1MsZmtapS54dnRl9tI
+HOOzFwNtqCP1HfE/sid3Aa7+QyNMltSGI51ZMm/QP3x4eAjYx9EPBhANg5uBvfrBItjBMjE8221
mbYN85fDDsvFL5ythsN/S1mvdQwnrHoJZbuq5mYj5PXs8HO/MB84TxikSJeSrtnX5maONCovxAUX
NSNMknre9aX4FYjjZeXHTieAxxFG5Ot0NI3W8fa2pVNQ4E6/SgY4mAWFopIYWimPlmXPwa+6JTn6
QLmy6+svUIE2606zI/ufwHJJeso3CF8Jbl0kuNx/E2NVbUMNIeBDyB0yfsHiEXTw993OK4+bTSKl
PEst02h4widQPJOL7ECvGg+ORvWIg/W+weDFSUSGDYeCH4/OhWppxirfiBuN4dtQe7/8eNMBGgkl
HXSO3QEkdMkmNy1uqgGCqXGfC3Z5sc3YUKdnG12pDMeiBeBFoIEZfk5p4mo6YBNumhxl6uOAp3lf
BiepkLuKb3/xfH7EPv6RB7i/ebHqnNbpX0AjFGAAdfm99SUm3SjMulFFK+SxCKj1IDjs+ViM+X45
PL5opFDPaoceFAcx5FBvJY8kl8IVfe/xi+TbxaVQn0CyGyvt4xUpI5cALyxtEq76X2cjTli9+YBT
aXvJvjatTelpAFKbcupDxk/zLTZyMgvV/h/XuB7ywRlG+ghNQudk7qvoXQSS3i0TBDPG1lU0Tkt6
XycdDknxCqjhcnTvOk736cr6vYrN6t7vvI/hP+5NxaUzmOOtvrahtu/+7UKKwyF2HGSodD+HgqV6
Nwuov0IJ5QDGC321mTLkrCdI4vEg/0vRel8jWT6tLYfdSyKn3Y4rcYn5eVSnZ7cW2sgFxqIIWZQ0
M1bI6gcQqY9yljnbDuLa7QqJTHENXRAXsrtBEmNnHII4tb4j6vw8kABqfqHlEZoraJvLI2ZxmaGE
FC49exiZ6DtUGLQ4ttarhkFXeuDH1ILELr2SpaMyFiYLIY8oD3vHZvKfCUnUh4FOmFY2txMGnV8G
42XaImT/DIRpXXCmJ7ChDZ1rW2qbvWASQGDJE4C8sMenmSuu0aHdAm+cv0Mgsj8D/TD/ovgLf93F
aFOExqSw023BhPOVhuv35jST1RE3XtUTDMWlks1WjDF4TIYxhOzEFb0TPKMQEoSHGnQzLYnH/iof
uMFAI6FK/dFqV9znOu/Eh6hbDzEHBnQaZ2GN4Mjju1EcboFFd3S90XgKSTEFktLnCVqNRb8HWP/I
gv0e0Eq7SomReV4xBn8staGrOuLvAlyFASY7Rq2pqH6/A79uMlM3GI0UO6Ht0Rbt5Y9MdZF6yEIc
VmrIj/CQ0UOtVvAmdD0pR5Iq9lcv0t3ihQlutuoxur7KQXsUkAGlE/s2eO/wFrLhwzYItUt/0s+x
Z/UiOzwrN9LT+w7XT9/v1cjcjsSTm3H6p83XZndrn36UWD1zBwjbBwHjNzCSkXWpM3qmPQlshh3Q
1RXgswHpdEnGkePxUIsNSSYtJAlOOEDi2DBLCn6G2kkuAhAiU7MJCSZ8WWI+sQuvdK1WPqgAZhOS
6mcPMZjyUEOsN7p2gOix0W004w8Vo1oxRTp2A+jK2MUod48fsgF5W1ejnMo9PHHS7uiuvTl7D4Qz
MSDQwYtWWMzkxA37XdjIpsQU9MhrU41xIFs6SXJEs6Zk3ExnwH7VKA+QafNYZ9jQ6va+GEUqoHhD
8sk0VFzrTpSqP4qdkcJ4x6PMHUZmygyAmBU3k+wGOzJ7yTMhKEi9uhOC7HW+CmL6nru2VthQ8mn/
lNlsYNKz+lCy01E4ggTfyqwp495CkHfKordLFjvRaimBFO/uogG500F/n6pmdmD6xCKLHXR2XZM6
yTKp3tvzxhUda2QkuamHs5IeRV+BB2vLNVNjl96DoOnRwxoNekH/7CyiMPnSqu9Z7mydQid+ADhl
R0/QbHGhApQMaSdZWaZG/eD8IsRxWCRGHed9ra2OICCHY0KAJtlVRCczQ02u4havuDvxnF+kRJmx
lY57Z29bUHUTDDjoLWVs+6CKpelVyKKcY+CtcuDB/uYI+cOOihgP4kj1UtOxcNsEVdaaXNAYzEFM
sF6m3HOEY+7ip0DHTm6YBy90BCyl6J/kTpyqEMRLu7I1vbZZFJVelN/xovMIHrZ/CtxMMdb6QEw/
V9XS2I+E9H9fqTDKdWzQowzA46XtvBBbQFYPwh/3jMRJaEeBjiMRLWkNBu8AnSu3KffS0D4JXVnJ
xSQo7dEr0Zd2M9M2C9k9Q3yexAFqxH5Lt6jC7FUkywLApMaibMiHuv21bhHUuIsPKiYFief2cvKC
uzrVoznEwG/N9iEE5euECneaGVNbmb3s0WCgzy+B1r6qRR6GWSyfrvbx03tiMqVFz5c6pvCwarYq
SMuEQ/U08d6ytWjtD7Lhv4YrbRwHiYLJsrW4LTnYRYtLa9rE4qeRuYisw4/7TjiOCO2XyjNNGH8J
0T+dcDPvn68O9dq+61oIZYD5QaiGjTNdHDHZyYIcRczmc5j7nHsGE0x/U9fMXUnHSRL5aB5r1Hx6
VuxKyKhNlTCElm0rrvg+lobf40ak6sl/f+X9HnIB049eWp+VjVWGUXHMxrktDPm4RjWrck5L7EB3
vjc/+JC4YkXbJTG/GinndeZ4F/mt3GrEG6Ntq3OQyLxo7QbVKe43wEwpgSIORT7p2WhTP7aem59z
sVqYIckwRFq5t3koNSWMls7omndMCGVXBsbgToZ8wKdVGkqC90s51JUi8vwL4BQckdB4kPUwS8fU
j9qTaFDNnH7Acb+deiId3FJkmBcfPKY2O431E32InkTIyw/aQIv1S2FWif4I1SBbht1xJ/cUdmYs
q/i8A2mmlEENHPtlvdFVjyK5EOK6+P9QlOfb2vAgU0wewCjxmdLAynLYnzWJiVyJEjw0OEfH6pqR
syH9v1xlB16qdFDeJgKqg3ogI60pVmwGXUJqJ0YtVugOGgVPjEbQfVhcck+Y2Sn93defSg+26vBL
PwbaVnHmWSDD9dLLnvubtm1TS715OtQCtF8ClFIcCmuAII8mLSAJWE9dBqf+bm4z4KSz0LFU3JAo
dYBzBxX7KRJ9loG5UMu3+eLUD7jfSy6u1srtaUr8ZkSplrgmfulRyvK8EbJbgJlILBJd/vwFKvka
3VwlUqL2BWx6fG9D/3pLbSeF4waU08BX6C+nYUVn6XKH8FYdiwu0kCZ4fYEH6LTw7L8dg/6q4NWe
ifwBCdw1C40BZ7YgxV5UfZfJsJbCbNVMMUaPDzVGvnnmZmLvUPdK9EFUo//faOYIpyGJWDFJ/M4R
hzrRbqAErP0tqirEQeFjzEtvUb9qj9x2VqQTuWWrXegyLcfBkjoacakvfz5iY0ATJPwwh7eMdB6G
6t8DzcwNJuXMgJTZ/zk6nKE8cJ9tCmjkA+Za6sKyyF08TLevSylnDgYY8eAtG7egC0xWMEdz9x8k
RNo8zUOboQ6pOCwNdveB69pJtUjL3YAb0yzoBJTUbjkdGTKo9qmVE6NbxRutrRzb/Wnd9QkmZ0aY
jcFbyDaYh6Ichh3gNMKH2R6a/zGN1SYIIb0PuO0gylfpIakrv1x9bwblhq+NgBWAtdF5pYEjF4mN
tfzvTer01szTA3GDauXkKhQ1fXRF5Spy7ppzpBybXoqjjLTyLWb5RVx3KJ21a+j9ZiENleNfGqoH
+rTo4C6SZqkWPAE3ktwaxrP3isM3bI6f5s0Tv2DYKBkIw26Puk8iLIuLiN8ac7p0u0X1Mq/EDB9N
koHUMAGd5jtyDC9FIfJ+hhUbHeJ+Nld3WUblMrF8pUON4oZv4Ckvx94Ze1mojLZ6F62lI04a76TD
g8zduAWcFmP5euu/2CuvxBm1+gVQzMGb/i4gXtTjzHB4wJrInkEVY82wsw/G5HHomuieKUxu4Tfs
7aorC4R3wJxsFtJaXkaI53n6l3mO/SwRoIjURGY4/93drOqZGCk/jM8PKfAoH79Yp/iBwL6MqoG7
GckqfpHqUfYrZBGjWJKuGZP/1J05P5HGqgdHPmaR0uzxKUF87jawdBHNMzQYoH6elpQ+a+ubxPgb
Wi+xRh0vqxDd7RHIxvjSUlXCvFcyhwVqwbIUoqL4GhLLr41Z7e8NBUhMx1GdbrBGe6FMK4pTVmhe
I8g/XgsUH0Q/33hCtVxQLCbwmIEgLh5qGLFgUW1oJZxkPWQ/HPXhFZNvqy7PiWZW3JHMN8SAiF16
kDq2/7OjnY2Ipph+L5ot6QLshXQ/Yk3brxSWKtG/8AzB1YbbIQeV5Z0ByuVPo2gsZHfrn+Fd3K2V
3DQHBwnzgEqvdaebcJEtUNK+INXYXc/N5x7XpvWlfFOFuUFMNh4HnHX7+4ItTCIv4BaL0sWijdUa
cUhMWLPN6v4XACWA8ZS33oF/nZ4zq+BuJr/pVnyv/43wHsm8s9InWzl2ejgQeE6I54OEhm0lRjMr
C7Hpjn7AZtyHDZF+uBAmnwRLccy5dfs2cp6ZviEltWvC1zjNVl20UU4VQQ4q37Aqw3wCWY4qX9P6
VYeOc4SCFBqp2OpOXTC+hxn8guSRlxOke5Weyu/L9sVeWiuG746eBsxvpB25cMmpNAqm4NqqfC1g
0p2zCZbYawn+lNQ+IEmB/TdnqPwc/oQaBIZjxfAZ3/bMD4H0RE9HVTNmuEn45Lxzh7L8Ud1YqRa2
x6kmnrbSaODrYPZgx6vgWSCa5ifWW6mElAfkRxc4uVUSCmdha3aw23LUg5negosi3PN2SVuEFwRn
r9crFmT+B5G7XGaIGrWv8KtvsfO1KpU4xbxmGEbLajJaGyesFGhN7kXOsAQWPwm2UP2EroCczYvU
gjm3qoXlaKZQt3/PnH2UDgcNXS+YBKglXgkTsUSifz6dCF/CGNDZ/rnPKhVv22cHLoIhenED9NkL
ymp0SVqx2yYIJwcziyZGdntyWuqCq0xH8/6XfhFuJzOMz1RkXGOn3xhTjFdp6oGAcL7PXVBynGPG
0VDTbE9PHrZUf0vMZ8V1ha73F+H3XLdMOsfxFqk9xT7x6uQY6WfQ/D3kPQMZv7PU4ABhQUb1yxkf
HDWxw3uq80GAVsyi7wqTlKvfY2BXjmfsvxqe8ftZj8hskonj60tbnQGFNyv8FviOhioRyDxMFAby
T8Jwvn84tloBKJCzbEw8zZz7U/KwX7qnzqx5IbLqF1xlwYyKKbZfH+URl5Ksj1hvWIss845xzRFy
/tQKXUBVeb0/dviysAPUq04vYlgP2rsku/W83SXHGHbgF8LrubOrzhXFn/HG9cH7dG5BrHP9nhS2
H2XenlYzk57Ty/CQrCrAi6ipgJTCGw2nMvfP1xqUg7inajmY+R1v7t7B2EHEissRFiWT/9qpVeE4
1GnXNVi88rxHWtJ3nK3YyocwrIxhdEAjNZGXPrzS/oaXNpyEz3K+V4ntzuK9TZVHLzWi54DBVml8
21aqCaIFXhfFF5pe5kGPRHxuz8CYp77ntFhOKQmz04Q4mwsJUPLQPa0g7km7WrMFdbL8J00xIXYS
RghjQOnYJwE5lYfqt+EOjaZXq4cRATOzWlSg1PKz8hHEmy6uzPPPXObiujGmbXfYAG8iSGSD56X+
KaGZNNS8XptWVAT7iQcdXeVmYmkCe3fRit50W4yt/Tku+djCtW6sr+YbLM7pRR/Uc0W+rOCmNbuT
YGPg1s0kORTLXeuS0d/hhfLquH5Ui8Z0ZAeaqMdCx7HFhl2sdfbphQSZ02gyq9dQWEVByNwj20Fl
P2Y7fvqfJmbYcC3OFB721MvaKuqrV0W6HbHJBvHskq2gvpud2Hau1tp2T/6MxiwoO8uyBrA2T3h6
1YzLD5QeKq6g3WZPkBnERATLFHDCJEW27FOuZyX64sQAazROQXlyvVzm9JROc+zwVU+tBWsmSrp0
GhQUrx24rRay4mKtqHaugPV7mqiI5OMpG241A+vserJU//nWi3M9ZlpdSB6+w9HVp88zLcXVkyeS
WoZ/mv7IDoLLuTI7eB5Q9hdazWh/1Oarb6KckUgITRnFGtj+n/pgaGgyVO0lU1zqYm+mPfl74kJt
Rybbw4eQS1IaVOnvu4UGNl94b1PORUTkqqm+/4FxLuHJdTD8NvJT+QPWChj+L5kYjr1kAlZyotFq
2A9KPeDe9Y0WvIIyVE3sBzmAmoO/l0ZigbF/fC9KgPAe+QqQ4ReEtJgxK6ibWSMbqQwR4mNOr4zp
66rI6o6ArK5r+Fop5K4ErdIEonP/VFjKGtG7iq9FAWOXQ5tMgoHvFwaxRjFeLC13e+/ktaPAAcum
H5H+YfnJYK1i2IJnFz23HWvfpxeUmmIhIc9wimnDkeyfjwFLVLrWrRTuBhj3hc5pf2ZwtVwNc10q
CQRV8E6frQlK2dXabuDcQzQ+0ffGQEUa4bVTREIVmC5CqtPX6T/gboJjEScMoi3CjntnTrBKSD8o
gdulfyWEbIEKwUU6GSG2Z7gN+Y7Fc1VN+vAxQcTugU84NK4sQlvTzrHa5y8zwrmzvyWTk4+1KmSI
aGt+raLsrCEzLo59AP34ak6LtoVkksIHHDA89QJ0EHEcqY6Hd42eqYopm7Dg+85SjE6PTitNKFIp
IA4MpH3KqFGu+LrJ2KeWoYXqpROrvVq/D8N9wGknv08Ip85EA9QUPE1PoK6lLi/FK4DlRvH0RrnW
mXyg9KkZt7a07wFyjxTftaIl0IU6HFs0PV3h+poTvr6/0N4HqMI4BoZJl6ARAhaklyxAe7ir7ktX
2VanIMXHfFgSKKyiwG+5BXqR48Bi8hCDD/lgcSMKtI8lfRfe4mRWYfwPmFYh5mGoe3zuAH+OEysj
Yl1t4f2W2zjGUVYdMBk1RBMi6+szF7ZLO8WEMELFXwThUvacWqmpkcbZhy2Em3sjSpOWNbmyuEbB
Ag4gA6kXpWujjrh/ruQ/GFESHGOVv+TazGp18rE05HEKhSVjPB3iFIeDWptzBmt0AIHf/FLNefrT
TwUAYz/3fcSTcQs7iLDL6WbpUJb6BCRTQEbEyHGTBVS1TRBZgupJNAA9+6CcvQ6Zc6USvpwdVVtq
IuXGnk9ES4ZlEpy7xhAhpERynYKJlIZWs6avtbxczgVHtuJMPtYK+QCuf61vfDNOKIGlKtOEcMhj
md0zE56mpf5phpDlUsJD0VzUCYUCvhKSJt8TNn9t2In9YpqEyF3IefEI/6lPp7A6uJixZrW1MkAK
rr5zzlN3xlYHlUk9DIWNhPA1uGINwDbS+cn1SRGJ7dCH7oVRSBx6r1ju7Bq2EczNUcEQt/bGVvPB
CbmkoDG+vqGyoO9imf8gIHTr8f/xRhH54izjz13jslhD6Xio2RzCiSlIPbCMUNOnlgO7mLU4nviI
/Pqtyu4ugL0aJSeYD6JMvr6ccp7eEOSIbdyY9xlUA3JMV+m/CIPNdrEM5AxMSCWVczL6+T7+IeQC
894ZXXS/Nd5rU4uDAkSmqXsR650yzXZ1i18DGbtiucEyf4yIBFskp1UELrm9x06JdcweALCsbil3
pQOAnoe+yfrst+a+a7D7XkOoRQFgBE7kqZCyw37U+m3u9uqPwiIbn3pM+ul4Yn8OgZ86xI1rlTIH
fodMtsDas6LZZU4DHhLfhSpatl3S6i3SxArC4o75Dze2WHFerqC5jy3EZSBNpmDQyprgrcVXEyrC
yrum8tpgeKWU6yftcyad4NGHzIeXqIVBdSjL3mU+7Y82Oap+Z3HftTwWLELOxTYK0yELZ4HyGwl1
myZzaCh4Ed/wThRODdkKt7hJtCDK6dKT+XfSWs7qL0zmUmOEm87ELb9h6M2XV8RrvrXoQIE3OteY
wlvdJhTuuer4jIMrJCM2ya5ojeHsNV876qebho3xIlwQ6hw+M9gxl4TMmkeZX+64CbiT7A3AnAmV
W3HWJtTTSVs5NtEKguZMgRRsZppLU8T8cHPao8ygXqg4b23bvtB+qRXMOGrwNBRr1/qva7oLOD6Z
ZaLMpwL2/tm46WqHanM3JK1UHGqaN0D8OCgcBzLcqGms0++2zaTyMJsS5d3b3rVDdU1VdiJTYUi4
Kk0mLaw+kjYoDsNqN0mQ4yAZ2RuYF7x0zoncGDRE1jecF5ZFF/wGRJqVEVHSXYcFNNm4nVJl2qdy
FHn9gajXIn972KGDJgd0hfrGt5w9PQcsH69axzilmclRp9yWV5vixv8u5gPSdvwWVXC+y1B7dzoT
hMTDaFlRE9fageY1zd2r9Im+CCc/hQn8e/2U/cG3nvLPKH2cCyM065hG7+ifWBUNoepGOkqVFkoO
oCKwKwd54S6I0+E3dH5AdbxeYSyof+dnBDyBeHg+C56VUwstlWHl4kL+l5yTeYfVFV6HrWJg31g4
NVsOQhi8wrDyADarvlaFSiy6VrxVw74+5SY89cJVEnbkvxeNwNqJ5mytUDlHTsLWCafqqYhD21+O
V3FXB3UzPbqVKFfQ8GYIqwVkgPyT01l2VC6eMAqirkRg0qCljsvEoP1kmX8n39fwySBX9GzG3iOI
eQf8RNzjzFF99FvZCT5MEwmzAVaQ3EclBOBqUv9MV6yMryN5NCGrdni18QEPvRvYRK4Me/vdyus5
iDGcq5p2p2RbcYilSg8kObwtq3MMqPGNLGyVf6JLoik8WLXJPAWhgL3mDFlIp3nCXBuTCw3akSar
CTgDmsRxNFhcctzW9Myn8ux5UXbpGTaEWbvZDuxzVl82EkRYwR/i3MsxaOgfZ3S+souFFPfi52Gt
GUT0fNUQE+how63gtmYcUp48knUzDsQhzz52UANoy+zWWVlGivFg56RfVfkw2UXlwD5hZ3zuCsn4
izainRf5+mSwnQPCfwRuMqPLf4g11Fx3Mf3QVX6pXGmi2bt8LHdjY0N3B5gA1QAsrUHZSNZqNvaH
EUkmLQyUiUHxfcIafpMemxOXUtrf/d+1t2qQAC9i/2vHDe0TYwL0PTDb3yGwHvNXyadNxiE67Inp
zcHlSk4JKV+lLyt5+qeopmNZU5tyet+zeoloYNckAqsBRAd4u/G+dPxKUS0U2cQPsUj5YUd/UEDy
s/I380ut6pGF5cmUYP+0tnPllGWOR3ddV+JAjLfMaRrzXYnx/d3jev7lVrNyNhkU1ddSx6fiW6j1
K4fOSniu5/zTQ/Iio98B7ID3g+CM63APWZVH7W+IYGbd0JUzBF7+20DaqHc6a0FVBDSMIdejW8e9
4txLHsQ5m5fu8cvA6pgOvlKeiq8C6R4eFOalyuVaRaQRdz3Gqk9NtwUu1mS5Mzfzxj3rjQkNrrtO
DFn5X45Dc1rbpzV3koG7uAI5T+GrhiRcvx62eKXX4Dvmkj28bDHpSYAZwVVw68JU1eh4pVMqxiMr
e2gueNjTEzB7BA/s+JtPOOrkZgaWfGUFo3fKsXIdDpRPC0VI4pWkFdBXUbSOF2I1onoMm5viMv+X
9NwaZ8r0jiB7RsozGWOi70Z4raS/DLeajxbbHM0uG/TLJYbbbiit4G7YGxIsZYtBjHe4YfgPQDjG
DW4o/ZgPwtW1ykULERfifMNYs01B9OfEvWU5yYD4IRAhVHpcYDuzElaVIegwig0rnHc+/Yt/foCm
RWNiNyrPnbWfvb/tYEENl5wHQfRrIyLsJFyIE0df2ioi0IRumyZfKstn4MjGnknXGsJiG9yuDiIc
mBr1nh1+KFy9Noy5sG9O3COkc3OSRKbmq2dkpCA/cuwCF3Lg0OaA+u6QULGXZMyGVR0FHm5AZhrh
dh/yKDN66tef+pJv/sPR+rFMin9wQ2MVeJPOb5m5/feiVp6DHtIjc/TiBCE7JN+l+5fA9EFYN34x
0VBKLVRI/oCazRYDYjA81vQVDuk0H7tt4Mf2mBD3nKACNKT/0BeAx0Z+XP9Fy0zDtrAa4PL13uYw
hYHlTc3WgMaxptPZLGOibo5gLmlWqMuI9EW2X7psidmXs1colQZdFdMh4s96Fan1XJ41wF/GxjFm
fu0uc4fRMNh7T1/PdaMtxG8L5t682KsX8srx2W6nagnUzBUgEESQuF57rwsI8+KJE2SluPaycDM5
MLxHmAyR8v+KXsgO98yh1G3LF3CjFZqh6DPyAT3/VDiMzlG/t7F8jP1Y+rEpsH+kV9uHEo6MExHr
brCXYkBWVK2EuyX7Qen4nGey+WjQ8AyeHnDNv26A60eJIObL/JSGwOjDCxMrIX111+AikrEn5j6+
rxDe82qfg/LQmbqu5AZgxm8ya/TeeCQWHso0K9MJTCCgjZCxcIqCGuLWNXleYmtvxOnk+F8ODNHN
7MKw+tZ1JHserANlb6iTrWmPKZBJVyXHJHTLMeRTnHOeMnDKCygu+gKrSNN6LC16nMYkJ7xjOq4Z
EVIVPM0H0qPF6MSA6y5fWbnEPs28C8rw74RbyGw0Jx4PK0eW+bbecHTV6WQ0YLaakHO0KH+TWMhm
7ecoZ07AIq+yblOYHcobq8gNe6G1bLMGhEWuSFkg7A==
`protect end_protected
