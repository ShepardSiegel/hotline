`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JyL1uJTLeQenORltKoxVI6J87l6xaQ/OmqACMHXb7wrTTDOMQ4evIbkrErci+EwREJm1QLQPKNMC
zw2aBAK69g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pjsUZL0ijjfXG95IdmAKBqzJ0jfN8lhUU73Lb1bZPVHVTHR2kJUhsNb6vBAzglN5za2KXl2NtLAI
Xiuxi/HKM961xpjPpqaLS+pKAxxAwm1ByiOexTb55OS7iNpNyylWzuzH6WfPSLOvk08odk3Hks9g
093YVpybYeKd4H1cDZU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TI+2I4wB3b1rQxUvQoeKRQd60x0uw2a/zLpYWfww+/9oDhaIQ9RBmWFnSzEUNoX/doAUhuI3MAMD
CkLrDmTrqkiNJGFx8ncTP8CqJdojcKx4a5JPp+/EF8zG++GC957JIaQYmFD1qS6E6miGrVFoxuks
Prz8uDRpH2s63R/IHKsph4pSuaKtLNTkWTY8O284w4Tge91XCqkSkBe/nCieGi4jxbh/tnUQuF6z
F/lE67Lg58qArBG3l9v40pjUkT2vOrgn2ECqN/eP7HJGXCz72MDUJOjl04t5Hz2idseL7Md6cR2m
Js1QE0k1NQS2z5zUJqYalR/NDFBA3EqaBEDjhQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4r39se5hvppSF3zaex2FflAUfJ00DHUZZXqygOiAxLm0gfDlnG9FzTa6tgGqbNNJ6asYGXVqn+3S
RDVffGn8cZcJiW5ddeXmIdORzghtbuUfPG/RuenbcfCmNOwQiGw082rrfjyk58yPHkfER8UvWaPq
/RcKiQW7SRs9//yVksg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IGu3saax/51kgktjicaWAT7rQK6KGNX3rNaJ3MyGZT6ere0cV0KsRuIxO+5+hwliSADcVmkYrcq1
oZQaAs47s7lMGMgtTLSjiqx3W9PeSzAGHFsO7r8b/EW9Y6JvnrQZ/MhRGhGIxSSVhn7sZdpHR0uy
rVeBQ0hK3drlhad0hb2uVP/t4E4UOF+rPBtp/k3gUaZ+ID2ccoTFdrymH5vX2LowdXs0jUN3BRiN
Fdn1bN8m6BHLzVQ0ltJFrdDb2oZXSWCa/WJ2XBtY+lbGrh4A1vTAMgh39ccHT5DrlbKQQmUXkNEe
TA0X7MwiYjfe83vUhnNFZFtYMyJt3fXtU2lO6w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 28320)
`protect data_block
n0bizoK3hNkX2JLAu2JoWeMcMoQMxJ0QjCPwGO36VCDhpSCGv/Eg3n3gnM4fM5OU8LsFEuXvzsTk
r7BZS2ay4nuKg/FAojmDgM1S/50mfNGyXbNb7isPMUcGIIbUez5atF4BL8wr+zepWD9t9w/gCNhd
vCawIT3v8981y9JE3qpbX3LWu3yNqMCuXVmWg+VumT+zR/VaAWAm3xH1Bh3VS2l5z5/evtwZZ/4W
COzht6zk+Q8pq4kvav4I4f8b/7Xd98ODTfPSy1h1G7iniUbt/eSmKGD1Q/n8yLHXqLFd+fMzo7yE
YKJaeHnwJidrTjj0XKTRRxL7uZWpqQcWZHxKX5KtvFqs4t0r7dr/VIJekBss03VmNcHSiYYDzzR0
7Sj4SF6LOHxLvPYQO9tB2qiEqPIv5I0md/rTIsA9IbeU2SgW98tATRd/Por/8zevA4N/67jT3X2W
jhqM/EVOLF5zT1zInO5dVTRJMKg+bi4nw71FZxtlufwMjFEYyzvPSBSUBlsbAMRaYrw673mCbkPc
MEQZULMGSaiwW6OLG/v+7DXSl7nbcF2Di9S10b6Xc1CLCSgBd4VTBpU8EDEtJ8yJUwUNwFamJ5wH
YNJ+fCM9R4L1uoofWDhlgEAEQDFpQB45zmu2a/wOw/J/ndN0MrljINvwPgDG3sVBKqMqxymKM7m3
aa8GtKcFecXhLKslKCh54bdmNOh54kh7jD+em28UfIx7CmtfYTm2oVtGgf4VP8QXaE2ZSze4PbSJ
IKM6ftJ1cXAUCNfaWnu1qK3n+TtYRowRcqwmrVXIaTdsBoNl78gOOOqDXOzJPHsyMPzEQkhsiUii
aAZF/iacaBvYcPKw82WWUgnERTX2Z/+Ha50aC24xDO49wIAfW5h3fd8dlF3lUckP1DlTqsiQ4fzs
jABw9UP4GUY0BrSdiYfETF0OJHTmECzjCU3MR/iOu2M7nIx3n51bjNoYY0l2e7/qVeYSjqkDGzvS
os5Rx80ZPaQPoDi5Ex09UNQVF65TKfJ4wqxAJ/r7vRg4xPQU6Y5tq6iuLu156JM8TEzLhU3fqy7Q
0pP4cWf4ydtOnaC0FLjfQHPzQ7MoPkSq/134+4iAt+JpKRZFUea8NKgDNICha062Li3bDQUW6UnY
eCrX8y0Fq4iP2fdMvek8UueV4ifZuatNmgVJHGDtfoCd6GJLS+zzi/AvZy8bBDIfZcAp7j/jiTRl
URBrivFT6fAhMps0nWRNJYRrR+oJ9/wCi1CPsYEE0ZOKh9fmg2U1gGnjf5mfAUX3jHfjgBt58SKW
oheWfxIS1/GOBTxHHvlxk+ibiwAzs6JzWtd7LdiMruuRfOmsXpJxCFzlNnhfrivj7KDP8owzsrf0
wWeEJoEk8pywvlUIEXbGpAEIbN6CyRhln+KsI6WipXPQlZmWxHkYHZjG6pXLYk3NL89LxkVfv17o
WSTmDtMOO6u1RYnfW8kpY7R61jEbTSnHETIacmo5Dcd047WaLfEfPAAGZgxng9AmSmNuotVx1ing
tcd2tVwHg1b/2djLDtM8OvlxvsI24y/mu0LEe8y+6zp+Q3tu7Cl0EnHmQVGtaK9WKdgoqsTtmYry
/YLWuEeqyOIe++p1N9phdUryKZtYCaWGjcOQJbp8ll+jyEm4HYVhO4XWMUYZUcy5BEZHywOsIz8b
7gFLW/9vHJgrvd0oSU+tWGAvFEX5CrVBB8HRExDrSYMjdurahWnqVOM2KEDb2NyDymb8YSwAT8/F
qrDbT6QYHM6WUIsiNnTeiT5g3XO01twAGIEvWDPrtMoTmNXwH9H8ga4SGwCYtzsPI7R3OLBR9rtl
Fyv0rmKDlytGnpQTS8PONun1JAFvTAL0TuXYl3ZstVfh4frcxS+DWzgHPvt8ppQPSdFyJhQOdUwR
xK56Q3XfdPxvstqzhhd/qbslUSP6YodZpLtrtaI3LbzhBi51vg11/8Hbrao5s1Ehfyfjf4v9hyX4
ZLvd1h4xf90OnreQCkAGxonW9fuVp7o2rfQzfKlkBNwQrBIN5mtCaeDj8Jp20ljCIq/CKcyM4oab
uXcvMw36IZR1AlyqniKHED5eCUgCQkMY7iX0YajxQBtp+BCb3o08XqmcJix16uaV+xT2EglNquD9
JJwC21U79v/GMyp0Tsl0SxaV4d9aZ0qX0xV9S/BOtj/JeHqEkchv7HLTbLrcV43pjYiZkwNKxo5l
FSgmnuSI3bTa96vVAnZb40qK7WyQUwdPbY8tcpWI3Im6wKeNLXmVUM17FwY6S5WExkelEiAQQpXH
f8XNp+rOCg+w1AsIQTQ1qBaZYEZngZMw9ROyEzipNutek911ZSe8RGHkUwqLQ9du6W6jv/Sh5WCs
zkEBLBhV9QT5EOkmqKVLqu/2UqTbC/5C3oUYKi/OkbllmsGTQT+rXtd8aZO/ctX0JXWw8ghR79l3
KrnqwY177+Vl0lN1ElwdMGLWe7yFz/me4dQ6Z+hvySyjVimc2wpkD+X8z5PovwZS93x9D66o7oYC
D/8W5VsdnaEC7wwmDH4jpkbNQqAZ5c53CEDlTJ1ytY1oyRIb+b6WrBn9/PoczVbUoB3a9XDkAOnA
0seOSIEEkrO2uJMrFl9LPUt5cgVRLDJg+3FfsYx8nYPtlnaLGzjlDE8d3Hny3JXnjth2NXR4qvhk
jri2YMKgUryXuE4iroW+u/h9GR5IEoqix7Qr5b63WMEQmZxjqOoUe/HdAAOCqc7yv0eSs6pCPPTT
2k3jfQkVzfqZqIn+paZt6Ryo6aorwTLfEyzV3mAzSuXEyhXiifRpNaHx74aWxjWucnnslYx6o0jw
Y9U7CZt731Qatqd0cMmQinahvkACStPm1zYbKJtFipAIb76qm1ptEmLyJ6O4YdZ8x4myD4llxpWN
Urmz253INbpBaLAemKp9c9hTUB98+ghEn6vXbZoHVZHe2OncwRSVix7r+krgeJdCtNO+VNxn39rn
YbXeUa9LMXE1uVpmPixqK8HIpfhL9xL9sG22dEW3keo1JKITmetxqWy8VXD3V4lKBxohWkHewI/Q
QH8Ui5aoR4LbqVklJfLWDbBCXtV3/DaqzgL9i03tD4bM/scdaIUus1VnHC5fBy2IVlpWe2KvdZ4C
zXu9TKzvOmo8L7/f7erv1nsnWf3bi1ZwPUZNNfsTkAuOLbxTirhrtNRrSxeOOzxn3bfniqpSqAkh
XSUx0i6+R9Yl3pASs89NyS5rIWuakcdHu3E9/wtF9FOsDwkH+LyCuDHrm0hJfWNQtVof/sAW2W3J
Nc5cIjgLQT1FcRnDlDDRFp0yUfL5kyXiTZFDJFcZy4mKMo8AaOFK94ONBnIbHJrMdFuSeY/sIK3f
xfiT20zcIZAzs5Bns3mrr7uZVx+fME+UgMYk6cc6AdmdUFv22lXZx+38558zKvt7Gd4n6oT9ZJE3
8bmj1a87cR9f1EUHBlGSVQuRXHgC2+xM4/FtNTmN0nwYLuijALpFyLA7TwoGgFBN6JrbXqx/FQiV
rAa/Mroa4Jy6oca6kcXsvzIP90R1+ISnUlrZtnE464a1dgACICYuntHTPVoKYJoAH2jvNkcQjvlm
oA8FFZofynUleuR8HMKoooI5lOIJ/c/Q+PCC2SdUk4RKG6K/0ZmoAe1ZLr4JgpQgvHz69+PWKp9N
19rCSMC150DDMUvySM2c6p5RXhfZ1SF9l8L5orxkmu01omrFzx95nxKH4PeAP3BoB+57UGqihPXK
u+/Bug0k8iCJhXuqdXwuZoMgL6Qmd2xGVLFwobEND5wzd8zoqkswO754iYhNUDNvOSnG3XtnhJ5G
p6JfNxHuA74h0D9Zp+XF+lIlfL5wTc5C3HESbGf/jS+wAZQgDogDQzpctEWBCPniT3jo5JkFEuwx
B6NUmhB7H9e8EUj7xCWjV4kuWKWmJ0AzUYJ/Pfu7KeKzIUmkBXIL3HRskiw3cRBVJgpFh3LucbkN
u3V+tXN955djwkf44ni912CXjTX6mjTcRdewvjbtyGtzHHgnUbK9ZI0bo1to/7o11CwhEoaxpw0G
9bnNzCFLSlLqimwgtKjkdinYaQRZ+2Srh4tINWQenRd0qQFqLRGgZRArY3wdyqgWwaWcNLUIh+em
cOo6vwptQYiX+jNo5Ag3qFEKfL1hYytacAiqt9/VhsDLEFEqPlzNnSChfsucg5hZPcHMtiREldC2
kkVsC+cV54Q1UAnJaPURTGEQIUKD/3BU2gDAneV1NYNliQHifnQRC0vb5S+1pno5Y1xLhRlhff44
RQ8EotCs4V7Kl9gJ5cttc823LcKZDqtYnEsbmqlHozDNb/qSJpPQKadcMJ69RfYcCXo8hmyPQ5lw
5fytUpGpySnIjKQ6gGuviyFFHyhaCkTzZChrz5KOIEuK5xfwrrRYhag4hLNESers2oZIpxMtkNUs
2qi633bsngiJ+g6sJMcSbXFRYnS39fjb7/u2rwqHK4bnxhJ+qLq/0uWWuzot9SF6qW4MNlcpXrPD
kTIE9JHTdEzbuyxF4Sj2bj/lZp5YLLmQeU03YeLYave9pbAEEC3hwFQwG3davfA2/1FvXeSQlC3/
FetrAlBK2jOwP2apIXyFLLawq8S18QE1cNapy7DeJDzO8nDI6jEie95W8Y8wtdXp+l8LunTsJlul
kO7rv9KyPctH83eLkrQXeFcLyovhNn5ATUABSZgF2TQVKBVLAF3OrDEcOaJljbfv/vZImXQ+fyfD
oMqivarg3EPC9cJauzhIkefMv+19vcCC4GE7/Tpv0KFkIudoN5/5WM79XHzCtT11V/DgxY8WQOfu
E2vcps2u1c8fYW5fCIc0UdBaVv0rNXqwjx1JxIIwXu+ZVNGQxIkuMVz+W/gZ/JgYn2hPpS3ziTSM
oaldRLBAMQd0daI0olcfEV+TbsgGm1db7CvZ74zYddIl5EKD3EuhK1q/lWYvX8XQcv99svoXM3QQ
w0xmpzQTQPbT2tII2eU4oP3OwIXSaELQwW2S0JyPHtbfqbCSmUfnZPiNj/Sydi7euK6JaMmF4FxT
PlcmzT4r1BmhsHQSEGBvskXFcT7FZOlQjC9Bm6hv6LUuahMDZwAqQ3DLwMTVdKH8E7+y9P7QR3qN
JtYIvVxR4yqJ4WlQ+gi/yfpx7T60Xla4gS3pHVj4ezoxkX6qdaX0JsVyuF5wiwdWANK4bJj2wgBC
VU5Xonf0Sq0XFMOdgLsI7bKHqwjVBh0FHvEdLwOy3ZYyqixNHANCnWWoA1FBryt3yxfVV2KMaZhV
GiSwKuQVW02PVmxoamvXk9O3Xfrbwc6PjKQ/m28dleR1JBJRrmoUH9yRUlIOvcMzXkisk1CLYND2
SBA/4mkWB005AbOzg+q4ivnmqSN6BAwxdFsanXnyjY/uVH7lDQUb8PKqPLhd6peqbI1rpprOsYvL
JkD+PaypD7gvfk7BViVB5gGQKXL47cy5R3HoWrOcBxJ6/Lol7Zgr8TemQCbB9TKeyHQ9nUOj61Oe
bgkBdI8AkzLl1yA9WOJ7PX5CR46zyEO1k8pGZmCnuy/ldA6i6xoPy/cm2PzKQewpBq76kZ4u3Xj4
5znJl97i016CNVQOdM+og0SCrlfz0Qx15HuzK8QZiAHe4LiH9F+cvgBQjPfFlOiVBlx+jTOV3ZPA
ALvolSZuKrJ64ye2z4s5UfQzFkpzuabVV68MJM9J7DZ3zhOP9f6mTq8q80c+Y1+ru0KsHO5nTein
XmoDkTsylxkuRWTdiwi4j+L5OJqnCsYxdH7wIwIeyYS4Usr017IZW1Dyi2EggOPh8phQJu6LMfZi
1dFzBWGuoQ47FXp9c3/xhofOJ5wd4jd/nJFOxrNLwrDhH6/LqDc7SQs99zS+SDHF/3dDorp+K9OF
QKd9TFFbwWQSfDKQqXqDZukXTJP+u879/q2BhzjBBh2BvhVLyR3XUzZUsW6cF6Z6H9qblGoeZv+m
g+9k2jyXZTV7guCnJ67uqVboXMrPACx2AzGE2MjNA3FEvssmD9mhQ0/Wrlcv7SA1NEzB4qGQrxWX
xDJx3B+vA8W//7d9G94toVoBL9olCoK8H0lWdEdf6DhvakgtnUKIGEA5qcan1JyAGa/O1FKL3RMS
/fB8wcOsvVkdCDOoeLDF/5Ql610v01bUcxBgG4CbQ0qQbsQpPjZOnsEHyPaFoAxgq4Rp3GHITKxg
oZHd4tUUcGn2Wx+suI2X4ovVQZK7Ad0MBAsMEu9ZwXF2p1S/0VefFB7R+wsLMVEcgX9jn81ww6U0
5ntkOPKy2PyJSg2dfP0ee+ASOhGwC69qQ4+Jfl4vL2PtkgulEPLhdayHIirDuc4mIEaHg1swtW3U
M8J0tqcfQL0xiyZ9D8FWDDGj24tctmHyAhXdJjEZYEGCTCBOBlTJSnwMiHzA0ksj5/eG0ogS3teV
Q2fQ2eexC7xtbPsDmhVIN8DiXyfGtY8mKKbhYdfW+sT8fYWiZoG/mX/2GXhsFums5DY+McMaBgAL
ONvT1mZPW8PQzbJFtvea+ovRGB1gFhnH38gbpMNe0dlfWsa3vWPrW1TlAwH/rwLk21lH1v31zq2w
mPY6AVeV/MIVn24UHMx7XLuaa69sg6V+7I60sTEwb07iE6EKKxDI7Ib1b8XbifKBwvYwQTtWEslY
W1wLBHAZChoeTulBcoKpBEj6qv4wK5/Bff+pCFi3MevuHVupzyXWynIDBa5kRuyuJwAiRDbn1eKO
T1ISG2RPdQzinFLwDRUq7Duut6lHH+HHi9230NrmnMGoM3S75T/Fvl2lrh4Zqfagp9Y5ojrr79xZ
ZS0cLTvh9VOEBCIXeQ3WH9ZfwvNvy4R1lJAv9cjxVDCFkCk4SaBq/tF+Ndnz2f7lmOyGENIdlq4u
NVpyFKNqAfViukeqrm52eObJE0x1kh2yP+xJzXi+qNaCSxtl98Zpx8cfS8+WGA9AIWC4av0IBwbl
kD2d1lqGxb9bOdzqYHiZw/tV3Hiu7piZMNoKW/ZdOf8M46yOgek2SFyny3pX4ghvEiXXFdETP3Ju
BbH41hHYvTtmvNkD96Vo/Gk0SP0gxg+6EzfYh3ZzHVOehKx3j1MvGdWWynoQFaCS+cTg9+tzbaq8
1QhhMsbXGD9LipmUS/3YFeBtwx/TeXNfjor4DF4soINW8kK5xoBzFVBtRZX8SJpCZRmuULFQsTMX
+bjl30ETO7m7Le/B1pvD0fzgD+pmomrDzf9bN09ZRLGk5/GLSdoUXc5fWX8IOWsn0qIB66oaiomI
H+Ls2cXgtfdpwyUsj4UUp7FW4B8m9nI/KrTYylTs2QJ6L6hLxlWasyNoYdAq4ZxBDotcKHm2n6IY
dZJBu3idcOIfqfh+7v67SVsaWalSc1aS/cMe502LnuMPfwPCQ4v4nhgrkwoOJYdX4eU4VEV8N3wn
qyVLrHJnIJyoejqHVWwA68Sl9r+9aPP+BnsHENWFg68x7PUYQdfqicA+Foxm3hftizyNRL2mB1iF
94bmvBxtiaO2hQ5N1ZqQNKpA3SddWUtzJ3Ju1kmtLttfCB/hjR92chz0lNmvi21qO91p0+bKdn/x
im8zCcs/v43jy4VYCgq/oBcSDgL/LzUeHcJvCLDwU9kIa32vWD7qQFU9hMxMRmSXG0BIgSGVEZVS
9j0Gq2oPJ6NQrxhdROCGlO8Vg8QUnj+iM23GIK6HDOf5fE5IjIDtGl7Sotw0ELqXlUZYD5uWPvs4
BvO/ZZLEWMUbX81MeHsKalG1uQbXFI79YyFUzJOZXElZYura/PTX+Yf5K9Vy+EDUPF1PQiGn1i10
JdbO7v5rttZ1IPg4xswfYLH7IJchTs6WOO2qd118FlJNsWsUVdcWWNDC/GTBepFdTp96Dl1VWcS6
m4bA9hwYESIUodlcScYQSYm44cUtxvbBE18SkI1bxwESOfQDykRxUZWM+07Whwm+YGR9H1B2hsIp
k/OPO5ibtJusA0WH4rhm+9i04k1YhVqgtv7/kMlsHzUq9TiQ8GfRY9ig7vcCdrykvvEmIpusAjY4
A9Isg1TI5zQv4vdD4HdImOkwAKruta/bpc1g91RlfnNJ17R9KDvHrKuNCF37ubdyyMh9E+ER7y87
w3S8jpf9Cp53hl+AcSnMXhjVVS8OhQ0BXirf3bT66usQpNoHkmiahdBdq4zOh+84gW4iI5kCGqFO
t7ZxWEPzQ9A2KRHohyRLvZZfsyiG5mz3F68bacbpZyxgSZszVutD5FT5vahpuA0ESJpUyVcKT+BB
uhHjAU6iiDkYjjiMjW983Vf7Tfa50SydxoeN8T1/TF8T/zR5K/lpDtPCHFJ7+RfXzxYR5gYnUqat
tJcq/ge0ql1cnMTxIQs/llUHfG7/7csm7G8u2Vh550mDfbp5UBvLmZEXIjM3I/LBFlDCcmHC2jJQ
8Kr8IsitdwxBVnrv61VEdJYJ1AS1LAtKENtdDURBATbBZz9co86bGtSE7WPSY9cvTcYOc8DAD6TO
uN5joVixCqNhO7SJ8IpSfSR2PRCsjMFupAJJaiezNq4yC+/UU4ZAcNoqOKV+cn2um/MYDk7tEb8Q
bVaFIxhFWZ9dmhUD2rmxUrBeIoviMyvMGwdfyTH/tEo+vdYgy8SIFd6vdXJJD8jDGPOLMrkQc0jI
lKmkh2yAeRKy9M7zqsiGVgorZpSpPGv8KxLRkeRimdkZEAqBRpZiz9jYhp7yXdVl2FOsH80BBU6C
Z99tKazAsASxx7sRuZTJULGKdDA9C/fqm/0On2wg/hw2QSx0zKLwITQVjQSe+7b5c+LZfxB+RkCe
dMxC89qYCXw0w9xrzvA3SvmBZl6My4aLadJd9KsdrLbQhIOfosga3e6AbMgK8N/ru8et7ag8AucX
BgRDcN/7bdegcZ9mgG2pk5PvpJCLxgF0Xk8HRJ6f4Ag+k0sT1EXn9xZzBIQE5tc134PFQkNs3DKg
KcdYFns8J7ZZ6qcVcTxQT5GRQUuZc+pYUwAsdCTH9m8g/9dUPntgQfa2snmh/21gKKbj9KkxGZfR
5UkOirfE/NWK7PUs2nb/1X9sOQ5mKW6BJHxFiILmppcoOKdY4psldcY4GckEHIX5nl5dAKHH8p21
3lJ3vuBAYFRQBbYepDBgJaHt5kHX+k+lse+CdoQZfSNjtPPKgFJ9meRD4yDetHhAQ7pqj2l2B318
p1IKj/CRl354pObeN5JVzyFq17yCcdcNay+yq7NKUNoa70qawDkZ4I8yp9FTMbwsvECeFvgm6WXj
HcMCjShefR33Kg7sTLHpv+gLv0ENxEMiSDk3ab/7AyICqaZNg6psK10v6/yMgdZnjTv/29TxxQ3z
bbLuPj7KwhfNKd0AaLaY+f/IeCfkdCT5bsog/X4Fmii9Y2o8fNfEC6lXztY6RMKvzp4LiLGriSmG
SKoGtKXDQkP3H8yXdwhdN9IfDKRCxqBHNBQ61eerzmmnW2NOKlGTQxkX7J84XlurK3viRwxZCJy2
ip2KVQiZtAnjLJ/18pqgmy4M8nrSZ5TdTe9Flk8adU1LEughRJGqwZM0rvR5qEmvxy4Ocw8sAF+6
WZ59KEHltuNSGW0I20dVIsVvdLScmvTeI31uAdp9NPROYQgbUX60GbZewBrBLJBOBYTl2ruvDhvO
zUAjAjxsUmCa9A6jej01C3u+JD7hbTkEjLKFsFG3bDtOQO2mUZXVMPCBg7qUUAImNImzlmGP04tn
BUuaokAFwaf+L5rIxO5XZO/gjweT6UKvlLUgBXHeVH8b/Kb/QN28jvVuWVofnmXb5/Xchp/RDUm4
X92kelTpI85sRxJD+D57+c2AiCdt3+UxxrNk8rniek3YX9iWeX+np06yArZFP3K272gBLP3s4syk
U8GWXAyakDIzdB5h1vEaO5y29nOzT0K+RcciyAAJENR+VNqJjWmCyxyfBouvn1LA3JoGfB0Y4SCP
YUOHXGXMIsG7ZV3LtX3Hpe/ybT7gXGmnOs6Tu9DpFuoUCQ9hLqsj0IQTnjxChtTaU/uftPKZNMfg
OlcADpBDiLdq5brnZ1c8Oyfdx/hx9jHDLyi0CeT9ZjOH3/EoorMB1LnXu2opQpLEnuODTNC4nJCT
9FEwRNRkRRDupeiow01LDn/bscPUV/M6Qh7rv5GBOv8o6IbfC6gHvjBbF9pEZx7XPHqK81XYA83y
aNYAEQy1X/XIn9RvTnweSm264so+kxE4dxzFrihEGhzq2bYMa22eBhsGqvx49d4r2pLfKqEiGNoI
8GEqaxpYlhzwxRIisMWMFc4Ypyi4PIPP88LYUjBEFi+a3UWWlmRUmaLgp42K3YsU8JAnqMhXvtqz
pS+q2Ub+hPHKrl84MAD69dX/ViZYCeoNndQ9O2oNeZrft/Gl7U8OyoMwj5pEftwdeVJq/OB/BkVM
NxQjNYs5Lt4C+iTA/eyy/0qCnlsp+y/27wHKf7t7ixinxfj0eM7ZvtQZ8mgNKygvEJTtovqE4/p3
MVyTeRbPvuWuviKiVHyjHF/CgzxuqxJPVM/11D3i8MNNVLjkzYtTqYp8kwiwr6MUYu4ZY/AMMGit
lZWTUzlJhExSiitNQ383ZUSfeyq42bF2HzcBpRcgYKMgQLTcGpVG+yK7rm07PdztWX6+7r+rewsa
8xso7vHhVM+Y9RJl58m/u/XRgBYeQ39T2bkgGRlI//yI89CwgbrzGo1orVW7MY8p6v7wzrFKI4Ax
R3UoVeBv0w5gUfMsyTCDEzgW21/yz5XvD+PyR7iqolAicy1q4Dxtr6RcNO8IkuVvIPSxhgsMhxqt
rqSlydKVtt3l/Nik23fdAnPOrazDazC+5D5/NP6hTcLzZuO4FRsX7k9Qy3fJ/89XfrPjisNWbM6g
vC0XZpKBWSXFrXwjAPvIUzvUIkBeDaFgTPC9PiHeCVZPXnsSf7tL4fPDbpQM1dE7lP6Vs3+df3Up
Y5Ax9zvt0pHIPxIKLFUSeJKNrQZ4KaAmPLZGzoAnmR6qKxtg2pRT+C6DXQPSJOm7KjmWHF94N3VK
Bwcuk6qSy59IcUWO8rafU7w0VUMkEayRXfwi42jsp67lH8O3pO1jE8ajXia46ZUWmDFcln2uHgCM
04bqaNUMyHwr3sw9pMY+orIeI5EnqQ195O0S2OcPahM98XVuEBnyoD7NOybSPUR+rrVtMgkrgwMZ
1m/ZaXTpsXvuahrWMslRo/tQQtxT5UHUdEiPsIY4sbd0lZSsqqMYdRTflKXEoWP67rWha7CfAtYU
XfHkKGzhB9sLGSAqkPeZJ2qct54udfPsHaSbbyJqNRKUZT1ElgOfHfBgIWTXTZH0ugtEIg3VHlJc
dx96t8IJ38hOLWXAmuiDLacH3xuDpRKpZ0qvQi2bPyK3Wqygc9AFXRmQSUodDGXySqR1yve3SXAu
wOvKLYU9mCqJbP91Kb/74BT7t2MK6tCOzYGUEW1h0YJBTaa/oU+ROw2SuRBbcYHxtmWERBKWcBPj
2TDhNl73R+GgKlFqMAIIjOF2ZA0GtDKTjek+nEJGgz63Ag+Ac6XqSnDzazyOZPx4mWrZvwo+w6HS
hWdMHLXmqsCrqqysc6F4gYksDYIvK5yMuSeIU6WW9GjcqlgJv03TrCAia9b99k268zlEiEzKwIAx
sbdMPoLfDYospiLr5ELvfYVZmug3Sf35DDZPwJ+7k1BqYE1P6K4Oe0JPclc264PigTCAuZRX7nAt
sDshbsktKfaowDJSKR/6KQVfiQsbyod82V92fIszkLcmygvmn2HoLLEsscNW/M3W9WsNOv1VjDcj
ETVOA7/xbgSKp92lHplrYqtSJsKb9f/gmaXM5GYcdH1uGbylmlFq3bOcG3i6qgVMMdiaML1B4TiE
eg9hT7Kt1i7/x2+ao/bGArX51EZZjcSsNYmC4cPOQfS8orZcZjPT88DXjYestE0G0U3QCEheRW1S
Ob6Y84y+ZnyJeEiKRO8W9BlLVY8gQGFw2Sn6OuZtD4kkZUvK8FUQkYKG4wBXa+toWLSyoDtmhDdA
5o3yFCqXKVesdK66k2Sy9mUGrc1dNCUCLP59uY6L3kEtp0515tO8Ir4VDedPCrtNnSDpp94ywNOX
9QytcDyQ4o71B0mWwbnwOxo4oz9Aef/MrkzUcPdZ/hAmg+UGwPqJYazAhi2Z7h044c1ZvnjHpMBp
YIT80EGlZr2Iol2BM/Bamwpw9NDtKu1QHXs/MMIcY1iC3kftYofCrvPI4oYUyAjS4KsT37I4663u
udXNxJkPu3kgXLxfldA97TOBHLrsU4zotsrUGR8pX4ZPZQdUHGfts5AF8uKznNOwplunwt4SVzD9
LGa5it03V1I7ycs0JI1TadKOA9uWWxje2iwu8Ycs5Rl6AwfZxIB2XPbGPTkwNAQ1HU9NMzk/C4tg
riwvoGDfPq96RoXqWevzAjsjrpwhxP47ixmOI+LX82vfs2YIV8JHvubzp9YX2S2zzgPWeV3lwPhB
dh2LOzCBIHqI+vd0DPUmYN9+lr4+vXxtXrB2bV1+0pz8b2fPbdeOK3vOI03xpj67v5KtTgSjzRpB
9+Pu/2QKpzJAyJOS1bBnKORFu+hJaBfZTqpZ4CCG8cTnPy6jOAl5FQ49kFQpzIIIWh/gmx3uz5d5
SkeU/d8XUFoU0NLzJbgCCt0s5v/xsowYhvCmeJn/Z4EAh1Yi29wRAWjIOr7nFR9FTwP+0peOsyO7
vLpriOtWh1odi9f4nFChXPyITw79uQtrYo1c1lx+yiIynLE95eiLieYOwLrUeqaOfxZRfYSV14b6
uqUp5kPBT9DbrXo1/2yXL7yWc4SLV2l4Z9KcGtBHi5g4RMv+5EXgs9C0v7/BgqnV3E1aqF7S1J+j
WKsQHn1MtXyNGy9WAfl2RwwvcnHsChCUNDv9ItD7u2z4KQyYQsWtmYbLAYw2X7+da/pLruvOI2ho
w0CZW4EuLvc23prZQTT5mtgLvcZFNsy9Yp6mxWvwTc3bB8m6ciojpOVc1B04Mtd0pCGeYCOQUDes
GvFVzIw+eKyUTacZpR6177NIBex41uO4NWxTtNZywRFUJM5ajYpE2/PSlUx9FoAaQ910WUmZCOzN
1y5U3bf2XN9bkjfXTWYGLkDP2S5SIZ/R8YZRfVCsGan0q3wkOERQFPwRWthB3GFech2dIiMy0Fmi
U7UjHFumdLuxQk7Xp89dLyvt1lAyCer62ZoZquobQ9tKAEPaPxYNgbtjBvzplkXs575ponkmSm2e
JsFdLMcE9ymUQ4ebvwbGyqzxM/Xpdiord9oOPnZJOTTUXCz4AVwc5Y3DpYuswo78LSzSXwA/PlSt
IpCiq8LMV2ucagSYo/q/UnlrmdehIPat/SyHQqynGdjmVutNGihf9UHMzvtNtRVVg+BY3xH9xikd
raSs3llZuRFWBtqklwXXhCP75ftcT8MeFSa9/12I0BwgIVGTmowyi6oxND34aClxDsqlw+tUbxa9
QR0Gs3Ua76ZB+Zttj0a4qBzSE/zni/di+L1pt8X5CcbS7VWhT6/jCc9td9OJbytnKPa1awibe1uh
kzju8aYRZXvi5F9yZdxX+hHLrS7+3dAGYk5TbbE++PxniAup/f8vWDIFStpYRG2uBAGOIemgX4G/
sO2r8xO4rOgo4PuD9Djo3aCNy0GX97iM3NxRUAiUrGdEL/by7jxd7JdQbCkca3gLa+P0q1VTvYwH
zocRAl3HwgP4v0t1zDu3Y+FR0SGE7RDxRLiROcN1NL/s3+4QVhDJxvZTSG6ovpHpqUGUpCcl1Ull
U5WhN2S7M6a+WjpVZxEge2FELrhrvBFbdFeBcgxFJ/CFQdIvfG1pA9CqCpmTBrdqkiD5q8NTVWld
yvzVENPT6fBKjXn7mi3BR7wmSFTMEQ8g/11EFe1uGQgjxIoXxhHSRaDfQAWanSvyxW/uJj/2TDzz
hP7515coiSreJCeQEq+LNME1p6kGcJZ6bLRTTO2na6kImUoBd/LXCztAfGCIG46eQwQ4//0C7CIa
/14x55MIwxkzBv5BR/G23YycczB8lfY1goAPaPiUffC6a4uiFfRt1Y1NLq7GNFZgoU3ByK4m6v+t
g5pQkStWvcNc83wQJAXWgE2iQ+NfGxoCCqi+ZVrij8W8+pk95PJz05uRUBRbhktBjDuE+DBF3jsP
AG8O2QuD7+FziobFrjYsoLJRd07WDuiKKW4BdYDLI08JQMG3qM6pVJf5BsgTLo7cynt3MJnGb+xi
dOcpIsBGO/uBe/xHhgcoSaIF0b9a9Igpjewh6j24i22BUNsC4tPHbnQVZvLSIKut6vePXyGyM0GJ
tPQx2WzxKvEBlFgTnAgU8rtzH5jym+WlzyKTAKfuIW1/q0hSmUV12fyOlvkiJROSLxQJGF6Swgf4
eKxCJxQojnPKHDH2GDr0ZirmlCp2AF7TU28IWNw5/R7lxsub4OSF/gOzXQIhl0/qYnYwdZU5xDg5
9Ll1CRUYNdV2wGmDmDeKqYNbu+/RSHuqturXR2O2nS0/0Eh9JAXslKiLDqLkVeorcc+5EtHohhK9
6JtBo8LxnXf+KO/QL/5QQSHPBcSng5DWiYXk5+zVUylPMgrFqayyglMGhKJTz3QjhRIGQU3H8Ga9
ydXnWtG2CULnaKlXXqyHyxn91Myt52uWkJ1H+j+/iD4YPRwOZVlVSrHOAjNm/W5eSePkqSyECJfp
cXeln9GdRSRfxuvF3qV7+R3GqPqwa85N/NGPr+ePI7bOxffPyMxd/yN/SfKTTOgbjiB7gALmlpHL
099W5Vo4Fr45dk+GCAC8Pa/WvA0pVoazk/1vqIUNCESFFHVt5x01RufVaukW4T6OTHTM/kHo/RQt
1ESnB6d2JltQFymE8s1BqQfe7Y4rvjAOks4gwPtPi+mW49Zkos3EprE5UonfNnBWpoYB+3IJW6K2
oq5etdwUVyEwQISoTflURx69z68HE71bCLoRot7BjtMqJKq0L/JzA3doXS2QUpasx1CmulglssfL
vbmw/I/DnIQbVgH94g03XRsDUWhm9ZBBDiwe+dxvPN4P3OQMxoV9CmLJGymkW9xoSzbRhb3vloT/
sBmvlVut992huOWMUkL6VqJ5Nfqbp4YTZiCgr4Kl+miQoMyYuawErzTuFJmhukWwbC656Lxcg93C
wUklo+ETqdMFfFPsWBoXXapqz+gmJQ9ojaBUrQRQLFOm49dRJXllkX2Ot6zjeroVVyGVoqAMleVX
mzb1z+T/EBGIcQWehXTSaG6zJId7hh2kZiIa2XJRhyphar2LV3Dq5w9RP9D83sVA4+hXoWrU6vXt
I0vv/uLZtGMCM2gw2QXqOC93DUNFBe3TRkfG74VUm8IuRgTHejZ1soaoBg1xWPoJ2lQkKZc3Lpwz
I3OUnXUC4IyOqOP8lvsUuYN7/mhAPinQFwTuy7K/Nior0KSLJ2NSB8FBTmRV9DDpwlKvREaJto5o
SJAUllfS021o7K9iWxQgzndN1JW3ao67N49O74AWpGHg2+66YBCHPurY7FRd35khdAr2P51er3Z8
0wrhbq+BX3hYRVsIDQ5Ha9uJvMtQDopjJq0L4qMtf54CRp6TVLcuDPwRHhVji7XcclyRRkWXeGgi
MmRS4vrSzC4rTJ1J7G+PlcWE+zf4hp+bPALEfrCHiCp5yFFoiP/gjA7TOoPpPXCo3vnIJ0N6kW79
YsE8XxtY7sdCANgLlj4WUCc4UGBXfDZe4XuBc1BoTwZwsJ6Vs2jYcQtPYcz7XPNnQMbE9okGJuK0
Dfr3kwSdzJQHqYE8OG7rO9M6a88+f/IWZEW3DCUprF0igdpmkNFIVe+IhtvthlzUPjMsRVd2icN7
J1/sYkitCqDlUWs3FbqN1EDnPWJ14t8eBR/toO7+UFVM//y/Bx7vu0q0fjlcECSV+YQnTK+jGDgS
4jfDBelVO+I6CXAiOmttB7GqLHUlq/hAVRw7dWheGAf0tOsKqzyuUszTLeh77bLIstZYNiKZduXt
UgDpoBvIaNUH1f+0uOQR9TSqjtnZEqrAGTVFgDDg0rYdydc2xA08BY2bl8Ramd2Rtgz9d7AcBMRH
QD5WOCpoVYf7N8FdbKg5aDtCMSdN/17SGLscXLHK1oR3yVbtzkGWjkiFuCGf/Gih1XjJZTJXBNMz
svbw2zeieDKXEA7UtUSDCUVcMyQwUVH1Zfje+SNE2clM/Wze9NoKpDH8W1EIGtCWbvrCf/y8Cefg
/QAzuZPg+OadHjT5UPFaltFc3XB2i91dCR05gJNHn9mR9GKtdlZvGj//PtmoVYeVlRo/P7/c0AE9
PDdhExmFpjSzblKk+dE82jsEPNVX0SI1/0EEeiLpp7yQvcT2Bh8e9DEG174v71PN6iLY+yb7MK7p
hQ8bACUCvwEloKh9ay3oz2edvX9zvJIiHtr1qG3Yhs3Xb3APb5MAraJJ0XRKQmpgcopVsxGg+qCz
rX/vlGzLBRbDiw4vKXIPe/V2MMQyGUDviinAGmEaWLekw69St1jPqRFEtt0SQUPpBP5xZEpgVxSt
DNZ9YUbQGzCqri4Ki7iCeqEs9VbvnHgnbHrmLL5STPesJNSuid/Lg0RnRB+M+/Mk9vE4qeruJtdR
53Vn7EyEiekKGjgUR46ZYkv4UzfpshwGNhSvD/t1EX1WCpgtlsf4Jj+D0VKI4MQ4hsKdxRDCIf4H
grKq9wA+RcCyWUpps6d3Sx7Hdnwt6C7zUr7iWWc2+EpQvpq8zd5AiazatNqF/RMhMSB9/EoxJig/
dc34PGFkDbG57o4esS4ZNVWRWvykCWhBaiywz+UGPAEmYsECoSObkfMGTPWa6tbRNZRDEA77Ti3P
gFPZ3I6LGT46I0ye3ttyDTuX9So211erbjvccVnS7sRIhh707yETZHu3Op8+fHX1DUEFXu0o2Zfk
8Va4aKHhE21Zv4BTWQmtwvgaDybCBH5z2l31O4VwjNi8F2u2u29oBRgnJ+VzDOLDLSgI+jttrOGn
QoDYyBMIONzi/Nq1V+WlkDl4lrlu5jOpxsDhjXSot1vO7ZWq+K/utViNe4BjI7Ik7gIwLL5NWV7/
0LN7KJouDCJAi9BQGX7QAOvNXZdBYLbgvW2t6hcC7lt8eKv0AaSTg+CrCFejd/tLLeQ88hMlBz6g
/xcfD8Oo5O3jAEMG2CdMP4qTOaOxlqHN7cGkV0FsAnnafTF/boBkDtQDftrYU0/5yxpIA8+PbfWE
+kVYTkQInx9frJKTUgoaBic5El2TYu5qV3JC6/N78yUsV9xGtC8Cffszm7iS4tTqtgmn41egpCu1
vv7+7dr6Al7rp4KrFsH+hIrhUd0+7yAxovp546OWhcP9Cav83Lj3GqsdsEacAWK7JnlYzLtXuxl5
3GWkTnjf6yCZ1P7et5ypm540tuNEtvZANbSVU0YRkrMuQn5zg2Ss4g+KIkKdWocaY0bJZRLMKHmW
C9ck5g66N68CBoE3FJ7+jGj4NJcK2RM6s7FiGQoZ9AYo0w9V1iwmVmcx7DCxnDdU+YnUa9clyDAV
hnvAhqQuIyVdYTRhbjW8+RxiJq+bg5oJrXMuOByDO4b6s4RG1844MMzm6HAa7dM6DYNuIzew+RzT
B6/SN2w/0xPcrWcLyk2VrV2GshhqwrW13MK1Ji807AGQ4e63QZgvc1es/lGSftwALkguInk0rp3Q
+AlZj72NP3Xno0h6DOTlse4za4/us2K3Z3SRCBtlryF9EZgYAJinE2Son9OGsD7JmRI2dNAMxn0l
iG79fp98VHWcPg0M81571TXOs8fpwKAiUcB+c0SntlF/xHnJIDvsf/PKniew8gqP2iK54XkQNZT6
nj92HacOJ2ZrQbdsRFmyH2A+tIF8N+aZdOZr0U9t7zDvPNO2uPS11AyYne6+K4NbJpmw2Oj+822k
sWxxGoHeVptitvlpAvVuyjdvBDkAKUgeCb728SqGRWoZ2Ah54eDNQnMV+xHNgaAGXRhOIXLVr7yO
ttcCUmaBG46PyvIZFDUQ5LLx4TLRMRQPhx0s2ZnmnR2SpNlGTRD6jv0hcvkommrTv7FOEunQLd3p
UQmw24PSqtPqtzNGHr5Cgm9q9xGvNUU1O7I5Qq49TIz7XUqMizJ77qhcaIFXFcfgqAnLdG7fCf/1
XCDJ+5y9ibPCpkgrs4vmo/i47PB7s8LxNjumILWcmE799V+B0Yii8eFEcr62YeurvzHvYdJaVvOm
2c+U9eZJBcfXaCb3SrS0qOJb/D6Qch/C8fXAXf3ZvdpCreVWNCw1J1b30ain2kYPoPiRy5YmnLyP
+SyCRHPqiEtgFCXbtRVEFeW4ZuGakqtETx1ayK49I76ckOIspiisxkrrXDq+Qrv8DhPY7b356Oir
HXOQZ06W74KQmaRaa6KCyxJfvinyb9GMyfN2tMI+nhqWiyM4rwpwuaSIHe2uQ4mD0MYMyKWQE1Z9
XxpkSnp82/wWoSEf1SmBHTi6BFVJ0VM4qK6S8swYlsXPSKsf7ruTs4ZPagy47cllR4/lahtvGKUd
5T4a/rqMHz58RvvI3hP5J6lxLf9UKNBwva/xOCnQnF/8FTWenUbxQL2AYkIexMmINfC2dIvuijLE
5K1u+2fJEBop3o8wdPJlPrSSRB8dyrotCls6XmFZHMWloqMIQtndKfsq0Ck0bvnAkwZwfLd1ZfZt
UOdkTqPkb1ziW4BrzlGpLYPlDyI/4Ruk/ECWZjYE29KSyW6dPZRJ+eXjuIUaXyfkmjG4yCgQ9AtI
TekUhZhpzUinM61y7m+9X2j4KD64JwKfC8BhYG+h0H/oAIecHyMmR6XkaORo8WwFpqeaPfDVfUgd
T6KPLgCJNRz2vzIA7UOfH9aZCJ2N8xsh0UbgwW+FYMX2GEsKXTbK6y1yisVeC2GOfEivBMHu+O0j
opz2MtxK/AYZ5cD1IvDJEzanNRFyGJa62BF+DjYeCYRJ6D05BFIzmZXz56V2MH9AIJfHCm2YmhF1
4ijHrf1kU5yYHK/oi00gN20eGcI4hG4ljLlXcsCyX/Gyp3Ig13W0Vid2cSPHSz7Nxb42mBqZUuZu
ZDITGdjhj7/E1M4w/Cx6D9F/o8urWH+lsUqs2pcdXy7lfQ6F1S5/+QlSKoXoDpA2rDctfLPrJnyG
tDCySEGkucdGwr937hPVH17tr/hi8SQET4HJ8ZG7eCzCiLv2qheYlVBMypBZLuwPq64wmn0/8gM8
I2B6TWZfq+V0876+++vsMFN82DzOdQilOJY5KdYuiwuQXJLFDxQN31GqeiLkq+/g9/bXHW/afzNC
HLqwBMZCm8gmR0dsd4J76H9pLlqoA8NYv9OGmO6D58mZ8NqzXsn7Pizhzm3cIjyZIND6eOM5YfBa
Ir31zGlg12r7kUGMrhJTBalGE3XwtgL/XzGQjBJKW/dNXTOa5+Woye/78k8gaFfhBfFYX3iptK7G
Ju9xacPBK4HnEtPQokjRx1FAgaDPT0l1ym4InKXLzI+KwwGQY3XZTNOCMVQxGOW/akcoOsu5F82c
4U5RqbM1GQ6YpFaXp/2xQw7+iLDDgZ1V0Mi4/3QKLLpVDNu2sR8ExONvlSELR5i5orefIzprmtFJ
PyGgINSMuZcwjinBV6nK3ZD/9uw/gEW/2DJLnUkBVvi5eEOM5oqXOVwTR8uM6FKFGaD485qpo5mY
iCLKoxLOhaWTLzC5Q0dpuhjBlU9jq+9uVvhhxF4MmPVskew26vlAiKQBE7nAyUjDozpm8jsnYlNG
uJDcjzOED1fSSADyMvK9NTAWP0vux0QBjIMw5qyWsxuaefzdP87pudX3fyOthr+GnPRZYpGIxGD9
Rn2R6w5HSjARjLZBOgLiQrTVb3dw3kFQZhyZjEFNYANynluN4lzwnlZDc486Z9c3ISJioNeCtXRU
G6i/HuCBoYgWl6PSDTq0XefPuzspPPRA1jFoibAJXGNCvRwhA/eFOzBteNUqp8RVN1J497f/gw6E
nDtD+3NemYH6RWSnL0p/zOgvizkFkMfwLJh0JLkJews1TMLvTtZrJty0FcytoEeFpBncIC62PP0f
OuwTiRsqJbHGeNAVktDhYii+yFv661P2Fw6qSka8LDBz9Vp8kARS2r3cNQmjcLOFvtwsgNkWitX9
pephDZva+Vu1JTZbK59LCBQjOUUx8SCM4i7jbO69Z9N0hmjLuLHehGZ1lykl1NzVXtdI+sblOtSN
2sIpiv0fxIbCSamIHLPPxxX77ZHP3tZe933h7tTuqYeIfwfYUhR/G27jRwRxoTKt5d6Nz3G3ZkP6
sd4lLz5wmg7Tx/y3U7HZq9Yi4QP72OCDJhEaHpJ7pBR+DCpcdPT/jqya+npz26+mIawcKpO8XnrN
YKTz49Xxl86a+rwJCbSPJJYQUJ1mYHyytP7o9CZ+k0rZkhtqmuVYD+Im4/sCWRovopsL4SDQgJGU
1Zeu8tsYJFbuV5yfmlCSOcNk+SlsU3+AAmbH71No512Kd8SspAy4MwLBN/I9GZJpVIS0myHpt/Br
USmskXlmpRrqgs6wRfsbYNbLSMGITf0Ta9Wa6bC4HwHxnrKSrQARgcvoYvHBRC1SIFu1f7Z8xRU0
1HyDHBqV4Rda3dP319nGg55tbaTXKHCg39Q9492MfDcAcx3xx9BMrOeBpNeRy5vAfIrhFgSmfy9V
1I0alnTG2TUPvg0nq/R8rqySoaQF+mkVt+7S6Rq5FLgD2VBoUVr05HJX1yVjZGCxDW09NeFIkL1w
CfFbWXN1IOwOIVz9zKBPsw3VkfB/pmiHusI+Icu1WQmje+EuR+dv/hmaDsAXgkdM5neD/e6zezK+
ybqAs1ntibsdhDWeNpu3ha9kdrrwlFP6Df21hoRxQWc1r/Fi/5QAH5oif0sgKLvTot9Z9QCakG+I
DsB+t9fIcpN2yzFhQb1OEd2WUDcnBL1KmWgkrUIwdCwfAP+JRA3n/f85he6QsQN41rkqJuL8zbwN
V/KPdq8+wIm6fPwCQzamzCJF5OvzAdyV0fIVD5IVnJvHAlrc7VHFuYD3qumVEeXZ4UsHtuv+inSi
oZJmZPxDTBkMBMVdNrHbm5hopKXXVT/rG6OPxjQHXoefgJwNjwgMl+avQSNadd/VVTqsxA2kIzWQ
bAV978fpZ9E9O1SyBKakM9erVB9zSiFFuKXR30WnLy1gKjAoSWqv1AivesmJFa2pxLaHBPRbBEby
ThZRffWvM0Zn1ZsdsO70DTVu9zSUnOAqOBDMmQpiVJ7XfEUA8SoPqMm3nOy/a2eEfFxadTXueXJ/
Srks0XD4GdBndJcsiELZ0Ft/Hn+xTKtpP2JzYIB5mk30pDkKNWYc3AHM57ZhRydlwfmHm0hK0DKF
OLwQMwJhLWjQIq0kPXvKAtXyKi5XOcFtgRIY67AomRXLEFAzU5b5ERPM6VEkEXD224P8LUa/16Ed
aAkfaswOq1rLDOB3iiKYWroTUnW1i836RCob8QLXayDIWRqDayDek/O4HdAecTdzzE6OciNXou3z
pTMOZFZpzRzTZ3c3p58OZVV0ECKJy5tR7OZ8+CuuiBgkutNrXgMpC/J+D9Yw1eiNLuUzQLjhMRPr
nFhXo+PxRHhimBWRKcwVs0Aj2mpiqnYe4Md+YRCho6/WkMS8ZHO7aSqjs/9jsHZZ1jMo8ic4M2Gm
DzzQx80XaLbiFsre/bRHHBk4JkFE7OgbdYrc5Wza7B7iO7JEkKlnmDeKZlm4ltXPUKT7LmH3+gE/
vM2zPEPIiXkrWLFA47FGWpuHjTSX3ez0kZVt6mYqroOipEvBWJm/pNELr35a0kA+LNfQH6VZQVv9
R/5QYVwRX5J/2y2XQYZhcq86orErRFgVGzsqNwrbjmsrMOmnJBLyrVLU88tCNG3WzLihsGnVpAEm
SN7mxXoaMY62h+7GQYvapIGlSUhUgvMHKi04iqDbCtk11xJfBbyJnUySqfdv0hlTvotyFAWf4540
Dl+MsksdfNGUCzEKdOpk1F7Dgs9jTCxWkQ4qOHxKuFt5Z1PZMH9o/Zv/IfnRpX9hJX8Oy+hikEZt
hUkHBLQCU/WazPcHIUFpdbtNgRApfHv9hNpACr3sZRPY4+OmyTewQAtlSuFyJXqdLxlH22PvuJaW
bGp+3H9M7gKMZBFHPsRKHoIhbK6ainwDBs73nd6Q39LH6YZhNQkD18QX194O6+ax5/B1Z7YAkUdH
lPNSEf8JYgPsCAiTHlwCQ3pkpYPGzURweFCYPovkE4/tl9JSfXVY3oTe7qQVuykZCuxtswEzpDhS
RniIf0n1Zp6xLVV/1pUMNxpT2LFppAnYxdmoagzRGJI6Giozd1WOqgJaj9PEltXr7QD/IXUqGaTb
CGn4oTVWp+MPhfJu+Bmt5laZKc5E/kXViIdk9zvQhfakluWWigxjEhSFuaE7TTkpxnd2zRZ5DdY9
0xkC/qj2DCsBS9u+Q9MD35KSb6DGpXJZvltrtK1bQSDWZw0TPwFX0Htyptg/E/4ZOrrPKt9ya3f0
WopXSMo7WEEyvqqvt2ZOtBl2Mba9cQHQrMQL+i8NmFVReSHO3j4xUP/bWXeA6/Gf8bf90IbCsUPd
A+4+qLgVVoEER6/mUN9/8Dz0nTF27LwUzfWtXVpLYFZHYMnoMbTcWF4cpdSOdwILhJZdfZ4uh+lk
mhzwvkpJ27L6FhqUVnIuxGhg2brhMw2kiKQpjcfskmgRMN97152ldKs/D7olwgbSzgZuxOEsvivH
dF9ZnQrP+9t1dF5gVoixOtVptda3Zb36n9q23O244CwCMjDM9RGnOooKMteab6/UtO2IDLf5B7Vv
H6yZ0i/97ZVqd4o4gHrXYiNVen35Knfzj4AU33XWnSzvE8Al5fRATqb/oIMF+D6JDRZAcAb3AiDm
WYA30n3plqixtqnxL8WstTP5ixRwxVryelxtlUJ5Qg79Iqr7j6oSSIbsk4Ocq3qjGocEA8pZel7u
IObMh6dvUok0XC2jJelUs5X4/L0vkQWWPSZteHNn1YYq/cS7NrZ3nrZq+BP0EYEG1FEY6f8O6up6
ZtC6WTfoWMyhpjr8fqGpVCSdLyBw+mKvqs6f5kV4Vw4evuSF5t5DnBUQEV/MNSAGEXSqz+U7Osph
HfIFLq4hIAkbiJD9USuOkar0+viiNWAbDHnq+c3XIVzsTBLd/AAlVLk0Wh62LgM+/J1gXG/NTxcN
YWWvBI+SvbTWw9/3csTrbXodhtrir26vSO4A+P66ATqONQslYj5Ks0xYmX0nijj4bZGdN5vx/AQ0
Z8Nf49j7sCYWQzT9cP5WKbPFnpprTAq9V7Afb3NHcSqniDrVzPf8LYm8NQp000w34Ctrw6rKSSvr
WxaVo1+E9yGwXw59PafXQ+ICLs1QkbitPZH79+OnyZ3AsvHoqOjcEpj1y8qqH0YSdsQxDk4Pw0rt
bf7adHWRbPqiVfwjR1FOt7t2paHV1zIQHWdJD5dQ0S80Ae4UuDA9aXUYDxPd9gGnSXTn3QrTthuz
4IX9xuwuB/LE2NF5gu8Drqx810AE5b6ApMxlhxasrf4v+glIKwmHeNHKNijZmcrsHZiqjjcrNfhw
hzAT9QmLs+9zk1oLtOIt/Y7NFKw1ejRiAw4xJS13lBfcuAhopBGwPZnBR8/4z2EEyWtTCuk9WTGd
bv/PYGmo+/rqBdDYnP9WMWk3ytZ1cmez8dYZ5HxmQEAPZQYPpb1JE7zvqMLBIMda7V4R2pU36Krt
giU+aRVJsgun91s4NY/5V2KDw0exdUWVkTHkV6TGyoHhPodiOxwWdV3POyovsxgBAdp8ArfSNhsM
PBLx2VAcIPreTqqWWE/lRfh3L219TsQQDZh95Ei8icTbgsaFpgGY4KBFgmGAUiteniy/Kl7biueI
1zKqn9C3XnPhe8TpHuBY5+wYjniwn4S/CECje5PyViD9qQrmT1RSi2wLehddbZv1ZzWUY+uPT2fZ
6nM6n1dgze0OJl6uMzOZf2Y5qfcvxPwZAr6Kms7wqywJje9XK1wMxZ5IW+xacmf5QkxVoirjtgfe
c3NYL81efGqviHxLsdFpLA1InvIhLZfvjrTmpewn1lqPQw9+0/Flz5wolY3bIMHdwVg3TgUxXy6K
FUR8ty/+E+XFKA2zEyXmoJ5J9XmZtb/6ZnkO0NcxkVtfF9CEOmv3RpvLgVNKq5YHci7sT+yGhlB8
PHTnzpQDocdaWfBpji4e+8wNzsMBL5VaRV603kF5vkR3uQBbzRxlTKg0egYfxgM0jdyJfST3ro1p
zyJJFbS4yLtCGk0/+wRSkAqgZAkl0vz/aMDD+O8RRbHozG3PvfpgiUujwKOYALbRrsevyc86yUTK
vgpfN7RT1ukhc8V/fzDX7KZl0CyPXLsTWgEGFwIPEyzE4rJGjkvIrP03kOunWBn4owRM89YXba48
G4UpCvPuUIybph4N0knisDZs928YKHTqzTtcbL7mz6RYIEzPq8zo/F78kzWUohQD2jAQHdaPSL8y
aB6kAsp+0mKRz7omsdbZ18+cz5Keomzi7jK0qBWSLvf5lEmebhQNzn2vinSvjEllu8+Wx5b9D+CY
8FD31ocwCT0qvzBP4+4crtxYrGSJMoCmlPOsyeBcY20p7mxMN2jwUSqK2Zf0RGH+pFP/X+X7dpzD
uw1SOcv2JfK+9iAStZBYQFY8BlFqYxHobd4Q14xPJeuWOkLFY5zi8FxC0qc3LswfOdYpnlUXTt1Y
tOHvD43q2ExxKUfXMFsMzUXD5Z/BdNMynS5Vo+QZysB0OJJACEWb3/N2cKgQFfspAbpAeZQ7tMBO
D32omd0fHtNuKdhBTEckXH9Od4X+8NllqctFrRre7yTMPpDDeORi/cMB/wJsAmPOma86rULsOyQz
S1UpyrddaKTM8hRtI0XFImV7EB1NZOEUWw6ecpyC4mJKvB1gORfGtIvyEHXRMBnkZvZTlZV3VqE7
DnvHQ8GRQZb5m20XZNie8ai7nX4W1H2keNeVkI1vcOm8r3MvEkm2rVID542lHj2TkL21hZWkfAKR
houzI+jF1OYhVICwfqt2H9hscQ7INVroR4MZlMjRrEbGZoZDvLdpEX3S/RArNSbdJegRgzMr0mAQ
6TkvVSjPQ5LpaewnXYQYJ2I9fom4czhECK8jtgr/XIPbhQM+54xsHwYQBpgT/bDunWQ0Sa7RwKBm
bYELvy4mnB4bu+CGmthxNlCMFH7CQM3sQPktlN2Pfug8i0OHcFxpO0AufSaAgNxtNjRKoy1S8Ksj
eNLzVQKPzZw85VzjBKNuYj5C7nCsc3GW20VX8QiuE3dKZRV22HP2kNCLrI+kfoPUtyxSu2L+aS+F
grNSbi+Lvu0wGwZSYSyvn0jcEwwwPgUk2AB4F5WU/6sJgOuWWry71uMJWd20thA5HusaO9EDdHPb
qznH4Mvkdm5++NIsE5QD5qBoeS8DOB4iNTxC1fb2bpBHnqd8dHhJVnsGFmKDnt3uqTR8tZTu3LwB
qkZVbYVARxsJFYlBit8tNVU46B/G0DNtunnPDHUtjF6h2qqguH013S6x4x4CNI3nH6qcpoAA1E4/
GKTNV6iy8tsJ3MdzK58edWnhCcA43mui++FBdXbrgLCrcroIgHxYzZ9/H8LLOYLlXnAXi/XypqkY
Sfoav17EMRLR/bc9QvoWueAWiRofJh23kOyZ7ZnHpMiiItf01S7JW1+/sC7tk6XFp8BK4PUEa1XQ
6412JiAx6fwP+f/5UK4JPglj74VPGKW6ZTplOtEzcG+1obPT25XPgX/Ht/UEXz5cr6Yfjdk5ZUfE
xjRaM1qUgeer+49cs3vyVnGQE12CnrARRj6vk7al2MiEtaffmOsvo60TRBUUDe67MjydEiAIM6b9
Swko8klSBy3Tz1kHBVfA9cRFdzDvs7H4wlbTPDC+q1bMfMW4KqPvGWSbrYi8cBRiayIK1s152/kL
0fgXePGSZhBQJIT+85Rtu+AcN47yX1cy4LZz12utgn0CM/xrteFPy8O92QcSu+A2OVUV6Iw0/Hbh
v0KHDKk/PcV8xO8Zb2qMEh7FGDL1o02J3u2nUwkIqVZfs4+5YfXONW+flrTduV2v17UOwZoD/E+Q
F5oDrf2KprCIoErpm8sWtAxoAHyXOiEemlaAplVKVexae5Jnzvvviv2cNIp2O6ptVv+TBO9Yyy0z
Y8MwobSeOgGSpasqsnSMQWbyteTvc06iFhrFolsm7WRdffKUNZGLS1+8FWD8KShoTtl62avghSjx
2kJxAi/gKYzct5od+pSeKmf0xphaAlE3WV4sRdApWCozZwM+woD28THg+YVVju3L/Rcat5O7SzNQ
nX2zBcwEuJ0UY/D8VXosLzDkAUuf21TQJM6eMK11zxJWWgTsU7uoAnov2wwQ3r7+oCv0vk/AhAOQ
mNzIJB/wQIaVURPbUIylx3LReyyPQSL3qBizAMErQpeVOYVvpqFqJgN+0Nvc2bgmqvRXSV0qD5hg
ECuyHyl3MNp0iitg2AHDpMxGZwJDspefrss1QWaoSnk7CpPuieV+yCKprmL5rsGANmhNgLH6h6/m
KT+ReeOtdRzPVHGxWAkjlChBI3tO8LKo6MSy/KwZZ8t5/wFAK1yIlzgbiL9eRIUvOBXZuMqpCC3F
CI7czjPKTgj6Z68n9Vwrh9Mau/cbGESlAmb1q4Ql+izuAzpZtFkU3/Z+C+xNiO8RTyB7+Bmbu00K
aEOvRyk6wRP1sV+0FSKTVpoCQMLE0mZ0QVY7rvixes2BDOkzcv9qdmMhmX1acOuIe8AsRdEcUv62
dmtHrD3RPfqO4BrCvd504L2QHwnBn/Yy2cGtLfUa7W996cTiOQSr0oMPNSnDkLbsEBeKioTtWiF6
y9Ir5o0PXR1LQ/p2lIzkxz+tBmpfoRr1RbBiMr51xARC9LFdR95rneUy0lSyp8AJzeWLm5+0vDSc
gy7v8/qLT5fqe+eGMQ8cVLLOVOKqdamo5Sdd8ZOXn2NkzJGQVOwL9L4nbZ60IJtQXJ2vJvLNEK/A
oif2TKerTI4wpNyK4IWaGC+lBt56rYHGMlvegAvYBhzNXSxb8MGY3kFN0s9VnLdixQIGoPQFYNlt
l2z+lstaDzwrvSQrUqGG0AeIL8kcZlg4Cfitr3tEk5h4ViP/3NbfiCO8JtPAe9QrrZMiEn8rgaPf
WE2k91U9E8C5h+VSgDeu6JUETW4zoXMrbhnEOFYAbW8dlOXyuuGrFN9UlDc4GHAnu44bCBxqwh8k
Ie3w58BFAu74dVA2T5FXveBILLQbFE689Vk1OBQpQ/yFyXiCXiSm8ZbT7y4fV05MbTQ18jcX9AoQ
/eaMgMmotrCAkd/6kvT5z9q50+NX5QPUBDGXW9GRGsM2m/r6osQGoSdIpTQqktJPrMa7WNQ0LoV5
XwirCD7nLi4y5VolVurdvE4/29nhATN1PHNZ6lttE+s08sPlFIndkfBKvF++yKkUI2LgRyhU/gOY
/S9eW2OTxYLtPxrI/CrQMfJ7dYZNJsnyFO9+kR7/04+/NxaTq5juCHN+0Esw8zX7pc4AVORz/dDe
jT3IrH+KFWpqKQeVOvTfoDyDVxAPE+AbJRyVQLwYUwbnloXdw1JiFFME3UM+ACH8eHAW/cz75SgL
R3w/yHCA0pGU26Y6qZvoyikyZg/XDZa5KH6NhrlJUVbwfcE0y0gsPBcax9W8rxmKNcPYUwYqiN+K
Y6U/3yrdnuQluZ7ogwMacsfRWhg6SchpTiAv4RwdICItJQaiyzLJm/Q+7nLXaUffX1HlXAHP58/0
9TGwfgrppSkHasVde0+LZVf2oIJvv0pBqKDCR0CBsDWfOBIiaENcLjz9kNFo2LnTON/7Oh0AghXP
iJANY1F7yDBrqq6Xzf+rl1tzOy5auoXYc1gfu7H06DLHO4WNiMOf6tyHaqHTJ8uZFM4/ICfdA+wX
1516n46d8dywLRACIPw4NH0GuiKdbDYdyMqQORu1CbvOTX0QHTn10uljqsReuRGGB99Eo/q/7A8h
vP2SZaKkj4LK4H1eMbSj1egyS1mJ0hsN49qQBZDygF9BTxFNWiWZDnzbcWGpak+SW8zFmbrtyVBf
SYVOW7vADKWT+vo920W7eM4BXivuOe9q2JR7F+wDS99keQLAbQtDnX+vRoiLvxyhGXflrHfDlOSQ
9FqQlGUxU0/7dLagecoDdAhbKZpzmjSrh0v+y38uHMCl81dCK2yDyTpM40PzHE2Bl7wDeAd+TDi9
7+7L2o/v3M1LSAKraXAc+iedEclCy1mJ+P9N86Aw2KKAqhW1laZa8iLFT8zrHf6tcSUZICBS27bP
cXoL+SY6TTfoBssMfM2oRabPp881bB97DUKBOIeNiXlJpZ7tMhRpJU2AiF4Vq2FaHs86gey+JUN4
rhQUMFF7K08b+UcEIrwEWKM80DL08n6RDEps83Ok6EOdq5qECqylvibjUvwXsFKz645duMqQnPVM
uTTX7NrEbfvDV3f4jMJb6/R3fUllInsOzu/girsyigKk/k2K7zW5L7130RYLFJB+crBv6xmMFQAE
t3cuidYBZCyjlnPS/ggBHu4b2muOneYod4lOp7YzIXl2vdxXROujSGkNYDIf0fvoqF/l8uebQKhJ
MW3aZ+mhsElwtkB0DbKUC12su0S7tKjetoVylwXfRIV3U9SW4LwdzN732KQY7BtT430legAupPiZ
b2ztg0Cm7TPovvPQyEHLbnNPrZXvFIdj3Xd1vlw2xd53GRnX8GDqFpMDC2a4nxlSAoUVVpertzvW
x53drgfseHcptOAdSZ08Cz5SL7bjGCPfpsiIWFCLkzI9NJF24SwKjiDtyBX2m0vlCIrm1tvz8qN6
DpJeELNm2YXIDZtq/z861YqcQM/efIq9UemY95SD0BevUPMEh+ms3FxHRmxS8awI+aYkOpEhtThN
hJz+MqwivFsqZOq8fkVva/JnUifdqG/ow7+Kpaqi+YNANnr6UOpdQZYO2WjQSB1oa+UMIegxTpi/
tmbzQIkUHRf9BXlmFElnRtr0xZFH44JyKBossWLtxtW1TFUC3ygJCvfxOZz4Ig2O2Hxuf5DWtcqh
5ycnew+NZhbJNMl3MbXB46dBK16VcizwWU0K+fswkoHwUmboplILSTb7LdiBWsmSDH/xIpy3kJ/V
/moKIVFgMJ81JlJRp9TbjNfhweD1mRTNToFgIwDkqc61k/G8ayR7uL5Svr/JZ6W4zBHIZ0P6PYph
eZdcWs448TstvWWdIcrCs78DCH34vQL1uJWCvxYItxazNdz7hDfyyvU+In3GS2riRsK7tMXyoVT6
EiuO+FZ2mccMb7lRVxqx1qgy0qnKV6vCGxLn10qDcdLAu+RlAo5a486GUJ0+4yOvXf8q1PydRqMK
0nd6/De2QfRxn9DZGO5oQHue5hYM1+GmPCM9oEQfTRugzEEyVhFgS6LOmzrlDsppC86tuEEYH3wY
ruhYQWVJfFXMDbdAJQuS13Ej/6WRCGBwVbcdEH2TYPvmZGlEUvcRQI8yf0fx6htyrG92fnBLUxTf
rFsjfK8DjSzfYLRUcCPi8gGU5WAdgSb2QyGWobwfThbQmZJgu+/5UKKffzE6UUYCCQSu2S67w0jB
yegQpxneI5SQYdUjIBc+35YEyD0A62Dvj/HHjLsbKbLXfqv3RevpUvdiAOjfRPsf5vpv1yp8iwUe
EwtfNK24sy1oK151DT/3N7NzRkYnD98Lte7n8XQtdHswplY4GLoq4/timnyQ7Osj1dLInV12u5it
8SMVp3O9SOiwAPSRpFqtP2sGLAQ00wpYc6YVCN4O1/I1SEOoZlAHdGu9kJ2KJetx8B0HBFHBz/iJ
UZdXRiSMaidvKGMa61oHBETB4AyPqWR4V6074ipIbUKDPU98PYCXefR5QVRMaXI+TThfqq2hUQve
4JFbQx6GLtj9JQqbhBMqWrXqVY5ehIM8V987niJ/VBwtvOQze6/fdN6mylbkAvj0g2tLcUE6hV9C
pESIvpxedLH2Y3xu+ho3OPKhx/cBJn31MbdnYIOZZY11cjYrMZc+7KryBypxZv+oxVQNfyYBeB/q
Fgg45sraHamVZ308gsUEgToBFZfjO6hJEEcg64QhzyCy5+bG6Le037vzHGhru75lgzdIgmBrl7jv
FdQJAaJRdLj4hletLodvDXwhqszDM6qvtkQX+nHnJ8XfPflNrckG7nVcuEAlf2zAL0j6r6+/yiR+
y50tSJ7A8BdZXgQZMG/TKPbdQZukRVqiA3Ko8AFaJxw2Ma9i3auPJiqwnR5YqfFrTKadQUnINY6F
eAt6Lwo1PxXUCXlg3MoChVyfM+eANSDrQd5PHjrN7WzNswZn6u4BwYSEWh5DNe53SyEZwMY+BYPJ
RuEoVh3Mcj2UG7k5Q/bGDU5MEPNYBzcy2hOIWOdPjnV21H0JrFbLew0oUaldOkvXGeb6N7geKmw3
EQTR5p/Wrx9SFKnndWM35CwenZBgsL1t3z+DHJ/TXQhucbsOswOyGiixg7UfQODBiPjnUBQLBl+G
XSkAYcVjhoKE2kuWS/CLklfTyohVicvM3aijHNSdnkTWId6o8Iv1buKOF9ROWkaS/8hs5ukntVHd
BGfrfWBuef8DfHNkEebWzwPPoFrWI538ykUJRXZ88leX9eEuujf9mg5qjW+xzEP1Ve8qdlL9rgBE
Ozow456yDLA1xPDXRYTQn8/PnH6hO5ZNagkBmnUOYJcKktcFeAwfpRTiNjz/lnIn/B5RKHV5aHAK
Lq28OpGMpubxjoB6j1w/OU1PO+6DV2LWQ1rD31hX58+5IGWoLd1uqYnSCP42c0HfL+wuXSaE16Sy
hHVCLrI64MgvlFrzO70nVUXnI59i9iqM02mPcL8JXYvM2qtHDFxiXgym2ruiiAhCScwvOm88MbX/
dkdjWch8HET8px+ERUPMUrCz060NcCVZceRcrVJ3chjrHySfIuwil2FqeUB2WFDF1Si0AJltKGTX
G9H+Qg5p9uiZABQMxvAXw1gtTeTzaCjl6ovtptbdlsMq76uS1ASWomOxE++Fu7r/6aJedrtUG/as
p9eE+z9GCj8PkwoXb+V1hJQhqZ//HP5PvEwKZ1befxy5J5Suf9nma7Gdg2txzanVGTXm2qbrZuik
XEQuUsXrPBlCKVj+bpDy1ldOC/rtyEKeNL7lGZy995MN7n0ZeLzZGdb7DvI2S6IlzvdFNJeRqgxX
0Zvjk21ZQX9hvrjftTXk2nazF1FzOhSRoJog6HkuYN7Q3yPSsS06/TYS5KMSeD/JAMVzEc8J79pD
JzIuZDpCHh82isol44T2V316L0Q3TTxtPLpxuUZBV01N5yJ2NerGVyw5Rf6/jIACKURX6ao6QNAP
m29MW3M8YaN5rDHs/frV/9S475c+ppGgOyHWHDcUMoSLcOwM3q2hI72m23539LNYoxZGh4f+iAL1
gZ/mNwMaeN/P8ilhUhi1k6YQ/yztR3PqTtBIhRAJ8wDqGwr6AxVjBD/t6oKbyaBlEnz2Lr930uUZ
eUdNCJa822c4qLE530QxNKYKn4gd/tujcVt5AK5NSPPIQD3WKlx6wVfMALVtlRlZg42fyGqruo+s
D/+43i1v8wWqZOlQYOSLJxUvGbib8CrufKwzSXvR+x61pV00G7gKEFOMeWGUN8rBVymybmHnSbzk
qinwftbjD0NqmosnXWdwMvAswAX+K5FG2IjbV0S6KxsPKpnoVsoZV8sq89UI6CBorKYSEiA7pL5F
nc0KwHJUeGxRXZL9kIzv1+NCVwJ/E5gZoUoCRkjt5FV76smbf8pmDqIr/tvUqd2uj67yXfo+OVze
WPt1Ia34A8xCYQilVVbGtMEMKpymAj5zjrcasrjw1eoxER3SXsJWJSn/nTK9vbucCkFxNaLwfkMf
4fD5tProG0kxCo0QCCu4eRetAQuz8Aqpnd/b1UOt9/WqladiEE4zvzMPCGKrn9y1F/Y4A51MA7di
nk0GCjqYwl1YRqe4uXLQ+ITF0B9AlQdZedCGrhu+y8cySayvcEsZzVALvZhR7Qa7b63zcKHtWGeE
W0r/+35dU9bQiQU3dBgMKDdE/UxJW4mY4a3UkfFmsX+U6BQvz8JGfAJPBFc0WBjNwPc+JlxGoaOb
7ppwNnDkBUBuOOSsYTdsXcakJsqJk+CRMuyJ1T14tgS5x0l6GjI1ll9hma3YzAn1JVNQHt7zA6Uz
ZcmvetUNdDE+qikQs7TUisQmt1ruXo4HGRQnr4yOo8OIDRIAygbvKqVW+CYYYKYVlWL10Cfr14Z5
KnF/PXU15Rsd8AcODy405DUdm/NBMwu8Yq8uTUW9jtV0wiqfgT8ur+X4QO0TQg6lg8AJ/GJNNSRm
lyuI+l10Sbqo0gRe5oH57gXkgZ/2Xfnscf4Cigqo6jE/AXaS4kaMVIz4FSjmWi8NSkCtdJaST9Gj
ofZ4m43EgS/71Mvzq07DOJm7lJSqW/8sx6/t8wlU2kUE8VnSZoEHFzfsNxcRqAFjo3DZIlFWhdGP
NyUeNcfiytRLHwxCuLCOJ8NjaH4kZoK5KwR+nBprITdQNFcFbLtn11zKjfjMAAXxcjKhGaE/eCwl
xTB2QyWXC7BQJvDv0HbThUq7f/RcxwhM7+n0dywqqk0Vg4PiVHH6Y9364n5yN7K4KZHf28llCnPY
e9QyDvnhdxA/ggqXFkDdbWtjBrWnQYE6MerOO62REfrXkkDylBkmN1cvRlEjvQ5Wssjm4kZ3Mdw9
GTqI1ZZM4MLgpLZd4PE+LQsf3pV/eKXlOqs/OHzcQ7QZYN+bme40b4QE8UMNWb4i3iIXuNTcIO0c
rWXsPHAJdRRpL225TCSB5RpCE0cyyyYQid2eOJxzw1H+sb1I+jYbcTbuQBgsH6bIaxn8DQR953/T
m1fBFNZx5d/u/f1M7EkxLo3OuQHXOP9Hrs02WROJS4iZ7o4J74WIfAKX9L7cjYqH8yy7NjWHGfMD
+LNMTNJG9yZYGeEojWCg06BQP+k97m6wBy1U24YERapjceNzLY2XjZCXwnFMGV7JFSvOndbt512l
T/1vbKSlzxOkbG5Wagw/MchXxQ7bg42JrwQX15vQRrqJsjujyXFuZxiiKkV+KynDZOD+/BS+GI0q
jC+szfjU3mf1zrmTmpk+BP8ImSjuEwmYY0wBrK1JrLrseTNKr340wGU44exj2BX0lAjGM5IY/aFC
eytihbizI015fOPxmBhzg1Eyz2PSKQPqnFDWi0ezCjlgZ6R2XQSSBcn87tWPY5c7pcCmdFlBh+wn
Ibnd+h2QVp1NdcsaTk/Yu0Okgo+sv962Xg7DvJBzvY+vBTHQHzQPnzuJmnGpsuTTofr06nr1wEkT
6OgjNK5dYwFiTh4tP2/sl+pecElnQeSmQzR1IEPULxtrc25WVAuRePUXaEnC6OWEy2AIduJ2FnSn
jesiFGc9aH6xInPUpZTCs7cjK6GMZcJ6oDif93Ms40yEfho7kHIMgKzhGS6vUvwxFzQeX1uy8FNe
PyoP0ArrRa2qqDnugUzQqutd1rtWmTZScC3nTUHDCVZdsfZWYP1EwURuuBsQqF6MSzRm+tPNmIen
kJ4KFi/IXuz4DGHtACAq41jWr4L0cdiN6E9HuM9nWZ0lQSDW09PIbpnVbCrNwmeOGFDV5i0e35FI
JmDALs7K5Mh+RivIJjjCRiCCqWP6LRJlMV5jHp4MluBFghrpEVwJhXoWV65xna0ETrB3gkDgVwGd
zyCDWqK/r/aXZqpKEQUPltVUuazo7l6iTcDF4/AR8ttIGeV5CG8uP+dxQUOp2e58mz/OzwT9s5jP
JeomTXWtdirWmKbPIrMfldfIjeRU/T52OthrwtugTRLOaaouVmrJ9nKr6GPR/7DTAzwIi9vaFZBH
d6R7IR02fAdgFy2hEEJi+mvq+xoe+PDevdQ7DEw8F9UfxRL7+Jx7I5xwVPpuYfmkZnSxo6VTEHrZ
z4cH8G1Pi+JfhcYy8in4ouxNzsv8G1roVLHrPzEwTrOJQgGjs68o6pVD38mIYShPzRvt0c/qtByN
6a36No5kAKrFsXkB+BLx0z0mE909JuFaDeebjX4b41HfD8wAzxdYhESBkNCvtIEM7nMUeaM+pXlX
LA3wjp2nY1mP90du61zAdEKHLk+PiM2ELOCvKsIoGW4x1yjTBrJH75kj9JCqs0bVNJZmyV92O9dG
h3TTvUzO7sMb7Ee1dcxkHLXFdZnq7DXLCI8iH3KCS18L6tS7tBteB+DWuNAfkF6cKQiuNUi8u041
7I+QXCDg7Jd6KEeM6yFmvhM4LZLpijUpJWk1lpuMTy36oQapteA7Pah1maf6SC6hRkAkEO7rTq5n
qSSu2iYcwQYRJVxOf+IU1fAqUDSaz5xwUtONFKXywB6ZQ6CVkXI+gbMkc76Lnj8qkayleHchB66c
GhejiTfxq3GwZ9B+0847YgXoAfvqWxfP526C4eqfrvpcsDbYMstJnBA09Nm9uvzqCoej9L80qtvT
1epMe76n2KLuVQZlDLn+RrOdZLDUnpDy88C+kSB4ltWSAd0u71jrQmWHDTZgoTF90BP25AMhniyL
otrMQz4NnBFDtHb9by6m8B8cgAB1jDINxmU1HiiZ7PJ7F5duldlSH5ryUu2DdIHD3GWuYwBFD9jY
6YL10VjPZTf17h8rtISo5TeLGzswj1mK+btNixdAB1gk1vxxQA/4gTnGs7jG24wNYL05ZRpBAevw
waNAh7M92sL9v+MAAuYJnahRC2mIyvtNkRoIxiZlbvatIofy/GIkIj8x8bH3g2JKcmiBCLF0dsV+
QDO8H52Aiw5PnW/3DelyC/RfgX/4G9DF9INe98lywSmU4OBHkI07sNZxi24IdEET/FxRWoI/clIU
WrqVtCOw9SazYolIeJf2tI3hPlnfsm4aLiOLHKtAhF+kOYrm6Kij4U9IFtZA/XKiiASfkLjBqOc3
kTUVfMWBhvwEOsONZyRxSk5xaxhiT5PB1cD9cG1PLu74tTt7MG20rQ8T/q+vQuVmi84Z1tExzSC2
yRrr21+YACChtLFFY8mxbE3zbf782CMy2Knw5nBC9GMHAmhUJ7vahmuRoASyQFhYtskzi9+mZhHC
5eUoGWVzKNqV18RYKmgr+hAPqhvJg3OrF54hczLqkTEXxWh7ePCV5VbVTRTP8FkuO7ZI8nR8l8SN
UfHs51L4EiJQHw0jvmYCkWJnpjTTn95G9byxtPUHvQXD0OiAvSbnD8WCkpwrJz0HeNrzK/MmMS1c
6apti4ncP/JfXnkgHm45RcJnCdRC4vAjW7skjAUSYNf5LljoOzVYF5fNdwh1iOBMEvtcBfxwg13J
l6lKOcwSd2/UFb8QitrfKugdBic1z048QdWtNeE1Yd+oFb+neW+2kzVjALooX+OPn/juDDE7wmrX
xmZtdZ86Viru+D+JrriC39WB9FyKNevo5/ZXQfwm2QXEu6cHRONezB+PMcj7/9iUoNYy8p/oXwYq
xj8qJB01jX+0iadYjeJKFHbSxpqPdkcaA+hGwsqa+EmFJlrF92VzGklFhyoDoy+APu+3guaTkFKr
nzHG/vgAOEqLJ10ix0azZ6sICIBpeajzcxY9FF0yXlH5iLTuEbYQyWie3g2oS4EFJVyFp5zpi39i
hnVVch0sGqhUfUKH3feXr71TN1RrM3VK/HRu6CITENM33iM/U2Mkk8bAumGULaYOFPEk5V8wk4Q8
eLVBsr2yE87khWebZH7fsFJIDxcdSb6crIvzijzkC4hNYaI5rPAgclAnwvrFf99OD6nQ7TaWg7zd
ZM8vqlT4yaP1FYWKY6+OMAbHcZEAXk1pPGshmc/IUnGhE6Cvpe0OPowbXlfwgYTQnVRM7qEjzMbe
UqqT5bbcerS0vJ0xt4woXYTrsC/0dcZXP+WsRIjNphrlRCxr6g370rY0BbOhAoPgcUyC2mLcB1NW
r+Tw+nTk62/jg0qY29RgaO9vfq5VWpaCd4vpgxaI0S/Bb0QFnyaeKq6vABBf2RP5JouqVtq5rUBi
v46hX7QlFSzG52Q3W4dTG6QtUvfgiOiUqb/qmOFBWyOnX5simnvJntmEjoQTDQw+puMlyimUO/NV
QYBGwxey+kBXD1cDQWdypCnE+X1SWzArKsgCkaWoji7dKB9hxk4BaoJqV/YIEddGifUsm922at35
QpXovm8FHKkkMpQgzNZpYMF33ybhhOwlbKwFX3i553USmwenV+aMKMzxW9FPbI0a91Vew+xCjYbm
IX45CMyiCNeejP8WqmneLgetnBcM5cI8XDLm1pVjFAPKeVsh6u/D4VNgaWwnxN70ZRaG0+lAiJB6
X4BJRpjP66jpZJys4D0bQs2hiRRd9aOb29IlVy9CMWFhnMoRIgXGxtR+eiNJxJAvh6wCdxa2c5d4
Fqjigb1F63w45BXVasgrcm5KBk1CW0GouPrYNaFqiL04a4RH+UtFJUu3xrrsg0AmBpcGUdLEQVVe
sAgxzlppsfiD5DEg0gIWm8yMThRfJ3FxfQmRAlqFHwhZ+9X+zRlfdVBYhpiGkY5gHw9B9GFJp+4X
HzxfktiEytWHIY6uRXUPfC9Litzcu9AkyVjrxC9U8WAJ0GZTGFllIya9SMQLySdkZ2Lssp9iWVEv
xJTC7vAJJ5R4COvv+aqmyEcEcXgBRa/AAxI4A6MrCqXYyBHE1gYnxL27zOYF4NYL4Ft3b9ull1xx
71BjjrXQrrLSoOwmQEJ719/u4Fqv1hO+yt6Bwj2NbHPDxXeTm8NnkZq8Dc4SfQHPDNa1vN1iT87U
1+hHMeo/ucSbSMUyVKbeZjsBHcOgjn7e8KIZ49xMv4Y3A/NuVPwTy/5VXF2F/deRWmX2UZlyavwO
jpXHiEgdihjOoOWxcWccfpe6OzBJW64km4HlciTD2h2bpwrymLxjTJiXBGyD0fyDb35ypJftk5+3
FisK4N57ahpv1ax8GKYZua/yWyIjxJG8TtpmNMgNuLi4rA3yJpOo5lv4FYsi7XjvIhwK/7L+b5fP
Tk2o8DAfvnNBLUcLr0/k//IYy2SCyj8BfFbt10s89JqHfp8Nh05zp2b72PCR/5j6hpNG1t52k2OX
IavtXB2cGEy227ZIVO2eBV1JnVn7FHoyFwi1lx2xEWbsWZLIA+KHQMh+wJ1NT9P+Lr0AFFFboTUW
fZ0p57mPIB48/ARmC03b72M0McOlWVKaUL1opEY9sGbzJdDZ5Yq2ek19pqNquZ6S6hR91o9nBCR7
QQ2bwmSdGhFEWBzvH1PRyP5rKde0s4ZESyNiKknqGnNkFSxYYW57fHyoc5EPSOKu9HSPzV9jJQHc
l5pN7LyHXQWzObZ2aTwspGkbGwwj7J0iL6BzLsLFjjEV/vSlmLYzIpevJGqxO8nI5bALpiBlaDZo
lpsKiIpNtPpuzlb1Oe2oX4iAeY4vtEqnR0MHOBWwq3Wjb/qF07kk48oyqggjoaII/fWBlrj8IqVy
0gqbiwSQlOCD43SssQPSLZQqrBGVYh8m3LRcTeUWQ9ExaFq/qjpvoqq5KSWONxPEbvWZZxvaxJIg
Vsu4+KHFulb9As4lWfbewD74Z2JfiuQRI1LYEAam6Q+sNY6k7+yzwQybrL+u9HmDNuy9l96wQRtY
xeFkc+THtxjT4CK6bfmMBBQ2fskXdoDtQLriG9DVkyjOkbM7dFziU43LUuZD9eyk+/FS9a1Ip23j
DeIj9ByvKlO7nOKLvyNG/a941aeHhu+5UnSo5SydWcRKFaTUY5P2UVeuJ8y0m/8AJSvYwHgEZZwg
4683ANkhypT6pB7JGbAiuDJtdNLZCyzinwaUjj+IoflSnlPe/j0StanWVMUbezcN1hQ/8ntBefQR
Fxf2GnCGqVOEDw/Saoy1+P4dyTun9+ak3Ywc/NOShEV7SS6khlgVEIHt8ywKJpf+spC3QTiYYmdy
K8cDneRDfBy25ngNkVCWgf+/NL3ZbGunpJhpbrTlaoKYBF4dlTVNOJCcOX2539t9
`protect end_protected
