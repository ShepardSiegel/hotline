`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UoAlkXOR5L4zwsPIXS0EgvLPpJwQOxzDb1s81M7U4dor5lkxBX0VOr2kr8064yqutmKsFOEXbWqm
flCwXf1h5Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f9L2jKI9OtEfnJnlhCQFlPWlck+XLODmx2V6yj3GW5PisXzx6RwQrQUhhDO4zJ8jAItqq5wPve+h
Fybi/n4skEtf4vOPGgN1N0SJHXUMZc5DS8QYs7HZ68bukKqXBoCbtbkJ80cE0q46NSToVaDEmDdb
eeeXe9uwW3Plxb/qubg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gydBinhdmIKjNWa9Y8WO3P28UR6Nh7CXXMwukET1tJUj5M0WO1w/i2JXg5ctasZAnVHJBxjq7Fbf
WeCMM7jW1l3X2xjY5XvpX6vb3f6QPbYZ52APE2UNdFGc54TIuF+Lmo8DquZUbtgZNlcY/mQUmMR9
On7y26oqCuQQZY6N3hJb0vwMXDy+uxoinHblYF/GYTWZMbLIgCmtSbUjbF6cNpxTcvjc4zHsy/Im
eeO7UYDzyaXRFNlDc6MSnkSnyla+eQ7SyTqBf0CwqfZnHPvewnNIuskaUGR+v77Cql05Lbgu7Yr2
o362pGNZfk2C42lICs3ygB7z+ZTN8hv1bsYtnw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hXwT2qdTZ5hdWPQD94JyqaCwz9/wgY0Z4B7WQnr+TCFDlC1iF57k/iDcNMrJFKWo9AdcEoOtUpD3
B7yjUAefWfqlALW1/K6oiWCYpSfWI7XLk5D5rXULB1UNDM34jHaSHRcthkLuCJatV4JhexHI4Jt2
pAy9PlCwQm87lMxjt9U=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GMtDHa/AvOwTGiJ2WJeyw8J41Ghcaj63twHxs21OemKO6+/kCz5LdpYpbNdlWQYHzrAaaJ4ziUF5
0QhMGyTWpr77NfRhypJITnKqd9/9745xVLPS6kaubYPEG/oEwaF4OnoWGR3xzz9K/40/Nc3bB45s
kTTHYCYKhUA02Fq6Kj4SPqA7sC5ywJmG/IEHoB1xJVd86YhTJ02weC3atkZKIg/ImKq/cNKGXyL/
1KiSjGXV90gikgWODS4Y7jnn08d80FcEqXQZZ2BPY9tiTWkonhjy+ZVGZyvNaf1XQ3mCmvrvy0zl
qseCaRoq5oSds/8un2JY8lYu48su8O6mPvoL8Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7040)
`protect data_block
D9xGwwTjsTNbW7WASjP5r80F5p48dSVyK1+1qlAWnKcCs173KYrV2/q5rmcZOWjKe2gpPTj5vQ6I
XhmabGpZS/oI7tAJQp7wHBI9rKwcdW/c1vX9pHDNpPmSX619b1KkKeiFpQr7cOXdoF5q4231Rjgl
tcvYcBRhfNFFam4kjPWj7pWbO+3kQxTrJ3N8Cfbw9fai1PNwKMl4QvoajW0rUEephThrTlbn9iWX
VXOLJiDR7RgNdTgSUbjZtmKOeamxxHXT9CCDkZ1wkSDgiYX8uD3UhDKvFyBrmavgN0vKzTUEDoby
CzgWaGn/81LTVoilTkG3hYNd7wXE7YeUQpV+c9o9I5EmnvxiB5O9skGhhxD2F6GcyrAiFe/jC8sK
wkDyQhTjVUAsS7WCVlj5GCnPvjHIIwi0NW0MiYAKO9Nhv5e+Smqw5N+eeuJnz5g5Ptn1eqRKpIN5
liqKnlHUqzDPdC6VH/JZaOjkry3hM7sEuK7wx97FhcGkI563xyRN269Zscme4FE0nKGGn03idDcc
aYcRTid/rh2GhxQ4Fu80TOXBGYj5RWwlnz8hqmWNEuBumQTYqakExJxVSnWgvONpqnH4+0mYMjtN
L+fX41TmG1AmR/s+lFJkP/HjDvFJBCgvW3s8Nxk3uVnRtsGSCrZUtl1I5DdhZrDzHvd4vlrERRwx
osWCdUT7laCyBGd+hoN/4L0+TrtB5Fj/zTCiPZKzWnnIZ40V1LHGsvJTaEsqH/wtfx7SWI4M+yNr
dXAUqf0npwBEQKKa6TznUM1OMOAQZwopQXKcD1Y5G2Jnf2jTADl5GOA7SHB6FAtya7TWiu5ZleLr
osViy0xVGtC4WpQ6gtpAVn2JBgtq+xDpJt3abIkbsoEAITJW1Gy5f4e3PLYPLJwcJzCWIswvPJWu
0n3axCQRD/gTEvhDMAWzKbKXQy9uJI92PlJuR/xlufGFQnU/53umIY/husdXinFPvuy3YANTcARK
A06x5gvf7A/xwKZe03pBOXFHg7YN+LDPEnhzBpCRE6/pDY5rx1y7o3BL0ZyYZAhRHTeLU4Sh+tpJ
ZbZ29wZR4U9iQZ9ELXR2puQVrwidnVLLC5fZ58y0XN+mfetshSwtT/Joh6YlR2DxB+fgMyGK1ORM
7TTYoLjSGPGUx6C+oW4tmDAcBQquFmjdhD6/qntDyna1r9xwALoCBC5xaN1EHxb5zuw94vgmDy1u
3tcojFO45VjD0csEnxe9Vlp91+GLp2cqgjtjqaxhpu6e+RlBVN086Ssd60aPRbGEsypLKzhWVPI0
HpjTMM3RUMqmbdguj0+TBAM2tYN+/c2oe0sMq8OiwvKO9RwhPry+LKg/xht3U1PBghHP/CCZkPFV
CIrT6qF069mtji1dXfqS5jjLYtfDAWBIrHyhSHDOqtt9p4oMdMxGoTHNyH5JIoJiCIxpO4RRENeu
AX28x9W9cEaO7p8+Z5vSxCk8vsd/nBYyZZDcSBrBJoRYYZnu7a5vyXnHWYDdfwKNrIPYMalHkH/O
PE0AXl6wGimH3Jhl4omcttKOWctVoIWYatFkNbLYKIAzRhZ2UAFoUJGDj1HbhCMrN8KLpaP/IDxK
qGjoQDUUlR7XR9R/m+lkn6lq55xlEvqJz8wl74TfvNmYB/z0RlhIRwmx8RA4m4ysIGDpy/OxE1yu
MgMIg3bcKYi6V5izGcLmJx4ObWt3rC5ejtwCk5sSWbL8WBOZ0F1/a2I+9be6SpvgsjSuEOQHXLx1
2E5oxGgpQpJMLwxJ1wbT6p8BsoSZrZekpfwjX6uGqLW4XhTyjacJaXL5K52eS6X7dDd/fvQ7DbDy
+vVKC7V2Kuk+82I32+hcOrDqqoy+q2+zdet0oWVT75Ty+32lIcs/s0ILpWbQW9FSAb2x+2rpIxjs
8raH++YIJ0OtUntpYFIF1a+S1uqpvjxHjWia86RxV6/7fwtHqgG0lXY6Rie+xbR3rY3FLw++wuAR
Cy6Qm5OkeWu3Rv7tOTwrMYp9Qj9RNHghILbNsHORW1RPIDAoaSvp8d5n3z//v3qZ2XKJxhkWWEVC
o/lzcLfwld1dfaxuXlxCVfDg3HACyUyGti+iwAYx2WyKb28hjcyHk6gIzVL80aU+IfpWQSJEX0jN
UO5laNlg3M0pHbljxep+o+2Li2umHsV8fNyFdVnIhbvxMoGucoU/JqMW//yxyA/n02eYVcZioYCf
yQ0Q1hMGxt34Ri5jfeS9v/BT2Bx3zQQBXN0JmAunWRulN2C7UzlGdjbf7/MktPcSJhJ022/NATgj
qMVUFsZvqolfu/LTtT+gJuJhSh+hek+2wUhRWXY+13+/Oo9x4Iu7QP3P9iTuCSnkBzD/jSOC73hS
qNvI4Nz3OgmueuR9wGMnU5qIni+F+BodTNki7NfrnFzbIeZmgNTeJAknqbFe5MpfVkKClvuxaRzv
byo6PDdsjbaYwK/UfmPfutqMcErEBzi1/oshs3WLrA1UlcH1SMOjmj2wluiaqXUYGfN9RdlM4/Cm
ajnZt2FXCDSqHgT3N7lfcljwVGZcm40uk208Glr8xSaHIYVKoSGzGcggrUOx2Oy31suEDYSJosko
ieVTXilVNlYe0JLnJKrAE6cuaBJ3cnXz+liXjNAG70dky3lHWn5/4q19Z0SURWux/2ypnjkg/1eI
PxTSt2pudmQOGPmGiGlfbADgVla7du7tawsDhOEWOvHumvZ1axj8APS6LwcHu9zaAhbAfYDtequ1
gKWn3TIupjI0zFs5YsPN4Ulit3YfKJwfn7rXMqTT+NihbB33KULbgGrqJDuv5WV58qKADe0CdbJ9
WB/kOeua4z5gZfPQVEsZtvcT+Mo8EXpj00/0iTdBiB708pfaHpd8nb9Ar6lLCpXnZv/SOOhQQZA5
nRZP6dY9F4bsmgqRcLmxx/azUgzP2MwqRd4Y4YVxC494l1XxPnzF5yEbCzs9HcXqGE15mCUtvSG+
ER6qo/x6rLkTlwoPWyY/7WTNaX0/0mL4dnHlgPjZJ6HsZxjnvF4tUdYWiFgkt2Pr1pqYDpMyAfOl
ldVlbUtpqenRMYQC+urQq4buJ8BUMUkCvHOsjAlOqfj+3GMNn2LvAG9bTHVTZlRq+x2zhyiPsAvx
DRkx2il6p77e7oAf7fPrqnVH9OfiEkgXwPrkA4oR26C2i86o3PeTYIRAoUlUYQvAH+3a1vjm7BSF
AFgYUvWCl+Hu6eIkAOxs9LEjCpemfc0u7Zo9eetoIs8MaMAVyg6/LmhQKirdkbTrZRKVLGPwUUgS
TVqukfsCAXsJIdPfgwvm99J+EtbIFDejLeeK/+R5AvK/deuCFiFuzBp8oYwJmvPJA9twOLTijklg
i6P/HDqJJEp/Q0RbWFLkDBAXcxcLLWL6avBYI2DJBhsQSK8BBCuOt0fzjwAeAVoz2mxK/8DZSK54
gM8O5RDbAczIl8865OdVWUU/Qvlzc2tTpllhdZeZ9O8fKmlc27xhqP5OjUCPaE9HfgMtbi1BrvgW
FdKbRHeTKtToO74L3iWwcuhQgu632t4eInUXqPKqwb9UQpX3slBfc/UMAT2rGhHrujtEXVhGiBMD
TmpTAoHhsesiexRkOfl/CZrJn8xVbYcmoLTFiuHVMjg1OdojGDIcecSfs3MKyaADGaF9Ce20cPse
AqGbsTF6wnQDWSSIuIhPFHNsvNL/sXxuVHA532nlxjAKs2YHFFtCFLWoFXkWKJdNlG7mGsMHrfoN
bJGrnrGb9tcoWI5LsUPMhCK7KfFiLWuS1VywHGyawblelzxkHLVMc5WcVLiWHpRkUFusWnFPHdQn
hb1zPGrAvguRq2B48Eh27+3jHJahagt9eyDf8j9GB+KonnUdNcH09InqdkV29YNBX0m4jG//0G4a
TRbo848tjsbAVNXpTXdYIPriaSkuTYUutZ9kOuJ3DKMcgaRT2QX6CcyBQJ8rM6ue2S5yNz7U/6Mr
qLaU3ZvPFpZVWJD/l6h5qqNs0SxagHV5EcQ6jHf7izgX9WvtDgqQZk36t5EpsUe2ER9ldZ9RY9pi
9PJAS3GZ7Nw/H+5E9VbQDFH3jKWhpJPZZLqU+3+YYEEDY+dRS7Mtam/pxR4YlTgv16hGlEFsYgf3
EGktEJTSPAHY3I9PLAAz69edGOZBOt2iN4upjA91/gKSGNjrqWTp31fjkqZAiTFfPq335nDpOKiC
oUwri+zGkJtm6unBatOAK0APdYC1xlVlTlaUcwQfOYzULI+EiYsQUw1kjGVDg0ac7vOFOIScFhrx
9ac8DA9+m6IcuNGlg4jkKj+B387xNykTZXaBE9GlUooiPtTDlNy7RUFFnSfmpGvFXsenisB/9sQr
mK9jlo2CIBrnRI0D4nRXdVbfmQbGa0o9C/PGMAvM5eFXm5madwY6rbUSighLT2RWCUeVDWetC/Qk
0FGcazUQInyeV+EGGwR56Yn2iYbUSUksySXkeA9P1jZpXHdIqsWbsNWVwFUKIH+soxq334KoHU1l
WMYhT4yDbic62e9wNglWyiA4Q9DDG8u1tEXQP48a9KdsUmi2+WZPB1pWNTT62+yq6BEp6clnQ/1w
Bas/d+s5gss3dwESo/Qz1umOtFwDg2KjsTzmU6zTEVTq7vvU5Rfx7QWGJrDUZrgoQgdWSHAm8e11
eOiJYsRFxK8Q92vqJnRN5rXbbMThG61pAJTP1C/OJyijN2ar82Hiill+r857SZAB0aAHJ4MP6an+
7iu9ymUMoHK1iKulAHhvWyz5tSyjg7fya1nqKdJsztqEDwvw5Twv9VdKEw7/fFtNbFPZoz8qSz5t
q28ovOOF+I3RX521HlyKmwsJB7MDCDvKtiyytpVK2/g2GUAAWn+tms+F3rZbF7/UG+eyjYadOe0R
0miXWFFNKj5DCBA0u5cTVFmDTmEqqgDk/NJXKndhNDVnCvANUeWdGlhHDfhNyM3SaTHVtQaJLcM/
jSD9HIpFbIxnnsIB/B47hs+fg2OmIsDpAsdo/7aRKhEXvSiJdc2NFFskrwhnwWDzh6lKE6S+aMif
tsmvrUx9cEjSB7odyLWpKynNstHSuhz6XjS58argDIp4qAUBm3j2mhzSSQCZdieCFirpBaJYw111
Jbj9VnpFPa5MpiKDvoQgpgy2exm6YKLkMgMnaKYJ6oWx/7fewwI/mYwBLR550yiaopkMB3NLcj8I
uqnGOiweAb54DFev7hIKLWdJN0ZZUDRXmltEE7qlWTSMpWowPZfK2PRzkJRgnQ83XLzaZ0EdLeKQ
an08l0wCJUzPpvljuejCw3LCwTGZmnX/y5m9BwC9CAfJ4OK1mM3uvVK78DHLorEh1dT8ZLhCtgML
ITvnZJmDiaLs8xzlv8UZrN5Bejo0AXoQDgGvmBUiHwomba2zGvwO7RUg1da3iNUHA3N1CSGUvjt7
ko1B+Rv1lf9mgXljwXz4MeAAs34B3Bkxh+GKK2n+8eG1KATSYMppycaiXhgjn89I4155gvY7JpIo
nuzlIbOZGET7FaXEzPOaUZZ3kSqvIKh1ZsbNjWrvlHWliG2ZbE+AuOXoxfwUULD+y46cPP6IL66W
ml2WAIUz0rdU2S65J8UVkOe0QxxgdD/2SK0rB2XA84ELGSpaoTszHkPUut8Gvtx4Fj6Px+gfKBd1
sgIrqXo6rGisXatRM4V4EU279M3FgRa4o0uLdEoRjoqPTbGtRABOA/LGByb9hjsNVbRdNd+hVKDQ
s2GoPnQuDiE2cq5D3qZua3Lc0j3BJZyreiVj6HATyw05cBxG77lGN86cTVcf+Ar9AurlZLkO5Sj0
9A+l0BVVSnobgXifjzIg/bfbHTp9EOnLcKBoM6rzysIwd4/3lixiTUe2CHPL2hlMVZ/pPHWGEKKA
jmgBQ0e7DdBoT0MwSWFb8L8A9NItxig1y/UJlqQe7EZfcIx+2lXq2oACx/7qu3DZNf39wX4Fjedw
1pSuXMFlIRTk4VhO9Q1P7S/Shc1C6roCjaoBzCfvBFRZnqh5PMSLrCgN0HixnAkhsgMn2aqi1tF3
k2KrPhPuL6Y5N9C+/uIZIcMGu084FerzZltbXqWFrVpfMqFwGn/fbXW7Xvt08krZXsh45LXZjbia
1DbwQRMK70oJwYXS6wFPSnUFdOAGSq/O+/gfPWwNzWaNh8sdkcYfXmkFEH2QfCUR7juu6MJXL/Dk
QvPjDBkqdsaG3Ir35YvGhvNsqRlmO66xVZ/EghmrLYBlk7J6+rXuGTshRUNSBVAQavkNw3965L2x
SzpSlXnIYaTOtQ69BTgeEkmWhDjj1j9y8MJ6XiE2i2d0pVShClfi8Rk2w49xA/u0oQFsvVxvGNoB
3K+JIl244tk/IEAmO5ZTyQproNr9mJWWNCC2mwtYgegVheCnY/0q7Wx0GO4RIotOSKVreI9xUoso
mq9VVoyA+z0u72WCFnTJ4XRH9c/sNTibeH+ev9LHYDclJTjpecLeQy7gMfEBw3HgcGvfRx8TFFP8
1Vzr1WAGkJIammVLoERajogQervAOlQviMSitYcbIZi7ygYqoyYWvSfvyRPSeeKP8uCvCPONIka9
afoApVLV8eTGQuXgeDGpcQ9J88kJzhwc1PWEkSiOaGZv5HXasapACEsL0F319rECVegzSDoXTZeH
h5ajwnKjYjgJjetLtzafIAVq3DmBcUjOa1qLULMCv3CNUkyso7UjXozqD9Z5NsfZX3DKxAimRODp
C+BQIIPtco5IqmNDiZkmErDki1djb4jattcT6btVtaXjIPbVp+MdFzlzG/TSNvG6liYxUv4+gGoC
tciNjDqVjhK8stWFnb+uA3qCj6DazOCWX1/HAdutYSZvElpuxE4QFeSTB/WE8RdhH5BipFYYeGMD
ZP/3Z8EyhUyZpc5ArIWN0qJAXyQtlQ0M88YYhgrie9/T3rTUJFETtOBiZV4ZAXzqJWqFuRTOwBxr
5TZ7pgJO/2WIZH40wRYXLy9u1E+b+9zI0uYEXWk9g2MPJMtTMPpG2qDtTnjRfBha5GBv3E5xqgz6
6KkKntHmC1TUDWbIh0T3XZu557FJzxXG1tSI8pyDQ821waIulGdtTHnqWU3xpWMh8XjDeZuAEQ1O
04oDLLtOmnHDCQ4wyePSUDj0R8/G/WaLwaworEYnEjldSym2XmNDWCpJxruHH8mCakkHT9rkIIQa
WeYaUYj78j+ByORZjDl45UO7Wc425cTrlKqj9W3d2CdIf5MUb/SwzV61X2X82IeArybxl3otVMI2
Q3coiTt40enigAxQBiBHgvslXLwmfZQx4IA4GshKyzp6ZN2wvYelKLML5Gm2SWLiA7s0woQpEgcj
nG/5+MztnPGJf1HVvOkhdzMG+47zmpXrTTCCC46rtVufIQqecRnJ9YJcJAQGWx1Epw7oDuUNJDlx
F67IQjVHMtltfn6Gvlx4JnhlfNPoe+pus+kxBO7Tk2YVBhfMr/mt2BlsATpXtTk1TteI+Um/Fj0/
Zcds4ZQcizzcntJZGqx8e767SiqgRIxdqJOAv5vGNkuS5JKoZgMIkMLkP7APgcE+B0OpAv/a/qCw
970IUFtMv2HX206+6r/G67lAD6bbK/aJNDhJPBzzNv+KOQSWZRhadaAQie/pRd0IdwfqT/XSFYV+
3bAK8bqNIgoN1k6a/xdhBKXkSYM1gUYikiS1TSRSb/76DQ5IcOtbp9VAKt3ZxFDyqc2G39agk2hy
YaX6fly3J7POq0Jwsvkd6Z22Z6DW6A9Px4TwcC4FCvPGZYnL3MSULWWdvb7LibgLAUf8yFewdJvD
vrn2uqR/xzoo6Wc23yCJRjT1if1by1yfQ+z9Lo06ZKRFovw0C5AGAXdVcKd1WYunIZDU25pAemYg
Pna9XMn5FkNnMYOFlE2in9YoBfj6CR7VCj7zpHgFxFPxuxPvKmzl2bFaLL3G/VFjseqXNIfB01lv
aH8h1sE2Q1VWD5mGsRWUdtQv3aAqPkjQ/Q/Qn1tfar9zDy8u4xI7vgVYKtLU/kAT8gKKbOOfoN4B
wsesQ/Y4yvrLypmhCSE4je8yd9BKeI3y55xx65RppoW0Uix2T8Eef78/RubAMWbympf+WiOvTcjZ
WbTg0V1HWSSMA/9xFijfnFxzaKx23Ud4S2Qloz8OY56MwkpFNfFbmwnSlGNnxQ/uWM48vtkGTjsX
4w7zPXNhwxELRUcERxJPm5/AzI0nS5M4JNK25BQEN9s1Mq0zJCI7h2qMTZvjtKH5WAG6FGSDgufy
AXLCrZevdpxQVKe6CsZPZBzRXFpgSglAeL6NTH3o5OrpVKCwyM4KDy8zidp3DmOffeEXCMxxJrx0
Jn57bVbvHDFiT1OAYJtcqnOiMkooXvHKv+IQ6IanerXV1MlvpeNqVzLrac7Xyvg0XC0mUJI0/2fn
Z2XSKr2DsigEXK+zaK7SewnopE5mAamP4M7Zh2iRd16dQdbRUvausyfMsdsRpRJ4w0WRHE00wim3
vERU2iJ5Y1l23F6pKZ0uE9vmjqdgwU0dhEhXnVDR3eM9Up2zCSbWD1/95chaBNG1z3+/gL/Z1nKo
kZZLJ1mT4hEBk4pOl/YzFCsPqRBZZDXanEMr3jc3KNs4G6MPgUtlS3KE8tnAST0/atoWiBPk7OHw
W7EwLdB5rT/mVa0MfNPyasy6doF5dHM/BxxmgU3K+DPIoQS60//83DZYUKDEPShHTLiKWflldYYc
5cXlkobdqlB6fRVsegvhTdg0RSuzl6XSxT06Y5UDpf1zoIRsTbeeqNNnst1TJBG85EkB5G5g7sZo
p5t6eCy4JYa1cQdtSzexruMDzfQz4eldk2a7YT2SMlyCd1lLCJtfafAps/h8NpOC/nEZU9Hzg6bs
MG8wHfDeJmVbmYMkEtiQ3AmRSkCPzYs9nwFa5J9KbUxwan4uMVAIuA8H2pPbECaynrAAXczdJAyO
Y/ETe3k3ZUcp1VZiHKm2jiPu+YV8/DIo/krOX+oqaFBgvHiujZGzchSfY7bx9LqPTnR4DsBMlcMf
OCIjcKU7AP6iIyLz10izLiRTK2S5lwKKYuOvOCLSmFD4ihlPR8IGsKyNnj/3Tlrth9qlnsLxhpdO
5XwEaOmg6h84ffjRzBpJf8oDbfO0khEJIbwiR6Zbht9k35p/skKdk67HfhMdzigHyAn67g0Lwsjq
RJLDt5395fytr19Q3anTMdkBkKqJm4GPqWD4Wme8HyIs5Pn82++NOoLToov8H6jTE0qAcUtelllu
Rp2ydFa3Rwjgyp8qORp079Qo6l/0Dc5EA28o9L5J1qtR+BUFUq0FR8FjFz0miUypdEWf3yoajrOZ
Mt01M9KXOybQa4IT9mLWcsHTdqTY33msjN1mc4C8R7yTxoEXH2ApEv/t4XShq0JIavJcFn/VFrKL
hJyaSvjz3gj2QTGgLKNX9maW327M5ffKM/PxBo0=
`protect end_protected
