`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
epOXkq7PuifqmhRlWNtFEyDBDrVtE63kjv5KsPjQV4N6yQNTRPu7iM0uxWOy39qQ3DyMqsO0SIk5
yJAZVbdsjQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
h3LilNsjSqKDq+EkL7O9eKgv4JEP3y/TtEBoOLq7ZcgwxQpkUGcrhzF8rZmr9eY1i/76eC8ilTLE
vOAyAQ+OcVCWhkTZk7nFU/fUKwwEW+Qq9X7jWiL6WuGv/4cJ7alXHVL6c/gb3O/NLcXmgd1sACMe
shh5w5xNMb9MzSgIPEQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RywZem1r5jKhr3aGvNrxgWQi9G/pj2yym/1lGyrQN5GH2CABv8qFS4uotqAkJxMDJq8tGVUUUoEj
wtVOkyAB1nUw4gc/1AWpB7/9IwsevM0pp4P5XJg17V8gpt8zpUI+483WRbJON8cqJ9FLyMiZ29hg
OsgIBCicQLM1qVFSwyCmz+tlDx1umckETjkqJ7aecZ4H9D0D0f3riN3BJHSmx5P8RF/Z6SNEWCVs
bf4oXm7ayjSvNcd+9/U/RamiPgXU/H7fBtPlKxvFlvCYy+1b5gieXRLfDQcapZm6N0CmT6YuPqSZ
VFqvURIXPhUMarnPN672sGIfB54NVQa0N3Gmzw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Mbj5FA5sHsVwAW4VyW0GIjUNZ+rDYU7430AFrflHMmfaMGO6N+dUVBYhpckg2uR7LPIFfddDEahU
NIYnYIbiuDQ24jMKBl2n3Db9/Xa9KbcxwoMRMRyTfOMP8zYkvGl+zFWAVwKu7bmddbQWJ9UW2h83
OVwjpbfd2QZfUbPsAdU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pXJhynDCVIf4rx3hYj8R1G5Ww+f7Z/G5zL6o531ZszndzNFvbnfrJuycCO0qFCiLR1hTOuWEbkBs
HdrhM/BA6YGQfRieRhO+/t0Bga/b70nIgZZ5yiaeeJwcZQXMORq285Up7zr2veBnXI8Lf9slHEzQ
Vg/qFXI8mNuA1fEJJCew3vChnCYh+iUIHMhq1BaM4k0qpDap8cJKd8QF93XJ0FgR+NOQalFY2lTp
qfnpwF0BW2Q7NPxSCRTLzZ7/mYsLz43QPsKz1FDYwsEwzjz9labuwYsNRBJjvIWa6n5IMkB5WAY7
KCgr6kqqlkLopUSPhblPvqw5EQ7jFWyH40wXnw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7040)
`protect data_block
cAEILfI2uPVJ1ci3b/C1i4LFEe/zsMTqfMQL0ZCpG/SHNeG7IeZR83clRJLMJzvqO/sy6hhcgRgc
xQbQzF7a6je8zsyl9pJwYRNsijmiLSUFcuBzIim4JOk1VqwnpCRQ3CQTbcqVqXwi0+OdJHOcb0Bi
MxAax3mt8zJ0Pbwx9Itwowm5ReRyW1I3pf5reLSnsTvNmuvgFf9MS1Ay++vBCi2o4u3F86xfwhrC
j3qGMGPlh5vFyU4oXUd4d3s3L9zUpTlk+SLR0pIBgRaS15Crh1t1Y0qO8Vq4QGI+ZhYzGntA3ei5
mDi4j12OAqOClWH9sOE6mEPnCxMrunEk8oD5Vd03evrTU6K+zAdje7nz4UhmKL1pEt8atwGHR6W7
o5xmj6p/4vwKzLEhUyWpTcRXTaBP4BKx+HH4JcS7n7jo4XL04hTsQhXgn7PS02pwOYsaCJ1es4v0
uKJDmzZvDZoUJ4PqZBpDLyxpI/PLI+RCh4DEYL7HIs8ao58V3RQsxW+deuItwRGc3acirxlAxSKK
tmd2Hd421QbTC2zMwWlijaCoEly1E+Yreg49wzXAEcgPxEARWIH2dcEIGPfR4ahDqxjurUNw+JzK
NQR6x8UJ94VuaGsq1EOlgr4cq4UiU/VBKENFZtJ4AnIe675pAKr8IGXIWw31H7j4HSCcaBUTQe4z
H5NCMScctZM0Y1Z7OEutoLC+hOGoq9e9csmbT3hx23aohbKLIO5bD/JzHWTBMrs/XpqNlGArYfVn
+vNyA6dhete7lGEIIQ57ASFoVluUAT/MvuFNBU3utpY3zAsL+e/D2KG5Y9We8eWKVvZIDvG5B72Z
NF3tdM13UMOb3g2v60o1eWaxRD/Bvu7RxvT9+rREjrhrmixytIb3LN05NyH6nplpOFfdPnh8KxMR
PraLVbRDUH5se4skGaQQ0cXoWG+qHqGQh5pA6PW+2XbvnMWvIFOgCZTdsOmV5kpg2J2BUna1UUIe
xXc97wUuRPf+otz2aqxgDDSGEuN30L/vqwk6e1iAOYm4PkOy2J9fVvGvTN4+wGf+IuMTAEZ4s9op
ADEmwLT4GV5WHEB0NUOj3vrZiP0a0idiaOthVj0oFki1tHjq80EwfAcP95kSOBrO5Hh8nkzB7PMU
ppBpg+LU2VgTIj3jVVI9wl5nxdKC2xl5Z9+C66HH2v8+KzZIn29A4/+QEWccuelR62yVJuO6M1sn
D659zI/Y0K+U8AhuXdn7bx/umBsq/L6HZ0vFzkBLmERiuvS6ONd9PxIsLwNOgeHVyQ94IKXBc/Z+
xYbIZEkvjr2E4EXS1YqWk7j+aChEpFPkNtzwpcr5KsqHbHE9lVxJntl4kLqqYcwAPZVlq60rSxkC
Ulji81KjS54IWgUCYgKPHlVR8expHiuUYqdz6+9ntrstQIPuiDA4IKytdG4VT4J5QsC9ltQvv6E2
6X5jnjJzBCpwzXeeEu0AGofpI/KQOAiP5mTlF7RxHPIaDTOya74yT80SxV+b9gkR7bfFP+LEQBkt
gPfXfxHHF1+Z2Hc2Z4xiHXysbkxF+OHyAymPY3FXEQLwzX/+5CRFCjB3K4yK65jPx/ULHWR3KLBB
HPMNTNZ/dokfR10SfTVNapOfSCxycKVkmf6HpxtsdnjKkZOkiy7ENPVNgMYNI066s70HP/16SH8g
WV16EBVyQQy2eS6JaDXEa/5wP8BFytE849KVIVaGnvrxmOeXqVeP+ohZozh5xQf3IBVNt78kAnkW
kKclgKAe3hDIhr0obsCoQrrCVyAzKCjq6XqC/ExdeQ1l/E3ixU+/pwXUaalkw/MutqtvIUj+jvJh
+Ic7Tu7dMV2mogD+mPT1NIRQ2TP2IubscXUYg6s6spUAeHM36wzCvc+n4FTfAgIZ0mCDKuVTDzsw
79jBWILh8rnPC0q62Rkto0d2azo/AyYm0BXiXRdjotEm96Rp0aBP4y5RTT93v82l4V98vMKlv9ei
Sl3SmE37juwC2it9Qr1uDx1On3/KQ9pvi2AO84642mLuZNkAdLOkdGWbpkNiOsY/a8rV2iOBM2ii
ZHZ+Ca1HL/4J/DQf5Y5o9EnGegG5idznB0DXDbwz3yU8185r9/llkrnvtYUJ0xOjSDpVQuRc5m2E
gD3VanGywBredQgHDsl4Yif73VVLVrsRVIrdJTPRASN59/JE48kJ8tYaCZYy2yI7SOhmY8/HmzLx
OtKaZqcA/dGKhO+V4gabjC34sQS2uUu36vHiYJ30/cSNX/14wjhJzo/GamX8n8HUabNxkz0AD85h
OP3WDyylRnSdj2HOJAQPDY0vsi4TO2nass46IckmwQSuct0po52xE7ZMDw8xeZK819zc+2nVhf3Q
TMTv0qSPZs0g+dL9lBYuUexnHg/zef1LCKpDeR10Ov39okUw6Q0VkPI/LfooHoE8YbcCdFuy/eAm
UKBPnqh9lT1iWBHE/SWUUOW9rEM83lWbKQftAxCZznP35WnQiGbT3Z+5GzNhpOJPmZZnSNSnkiDL
EjEq7Zs1cIWbvmZ+sjOBCRkLYD8dgCQaOUYnpuPQtQcHwVZEg0Mrq0DmqqvX1iI6DSQinesCaRuc
IN34jWM4+mfsW9PmcvdRrUYy3rC3f7DRVQDP5t+TUVxfdZcj148rBoe+BERaKKpKj69zIvBLfK5r
r2cjsaekJUwSoautRs85zqjNaFpYiksPnvi8I8p3HY9C5a29IkoNEXkugRpn9t6KB4/CzuQMVdc6
0zP7/Lsq3aXwJZQVb9rr88tFclz9nchqXpAeuqrVmH6lOfebsqKlUZwxDZKbQupjRq3cAbMUq095
K1pzvPsfJT3kvLf0WeZqFYwqcQS7UthY4KT9fLavk+tNmg7gbfVQGgZSio1URKH1tNnU9H0K8W00
OjOoboR8T4qSVC9bnNkrEauIi8MzMdylXsLrw9Waf1cQIrrVRN7cIbXPNAZ8jNldVsr63bBrcjwW
cU9OYM6iPvCUUpdbPxDb4TZznF5OWi8NeUOTz6DRRpTOJV/4K42T8yibrawi0f1YYJ8v8f+k8qzj
pgm8r/4KRIQ5D60uAREwe7XyG65AFVBgPd4usQE6u/wW0SOYOzpCLYILwXqvHUeioBgIusCeXgtn
sShIPbqA9rJUSzZrrprRO6YhTEquqbst1LOYjkt8VdLFJkdYkW5aV0CNGjmyNE92EkRRGhsvRhxy
xJyfJbYBLzbbWwfb4ti+XRLg/b+1c1caLYDJFxoO05uB3R9NQLB5NF3htwZFRH+9AZyD729aM1BK
jUz+ops4P+wmMl+b6m/UprW3WywQXHbXiYTXfgm0UUYPHt3udCRyeGaWi/Qi9uYf6KElm/QtNloW
udSX0eG+02mM5sXUadfM6g6Qm+87CzDgF/rnA2nMffR4G5aGOaMKDDF7fPDgebYBPITMfjgb3TA6
k2UYVqEzbYq3dlPXQR8u9QvWzETA5ES6D5oT8V8XFRU7c2pzlrxWuAMEVpgkO8TmN2EznyQAfdZb
XWuTnRhUeAtq1nWEVWUhTRjQ/t9LKf3Ypl4uUfPfCnUQDx+x4r589Rdq4jN8sw0em9ISlA3F93yT
gqwx58pjU3uif/l2TBqx5o+Sf//pavn97i2trCY+5rQwglXzhUw7o5qKExcWOw7Kr9c4QawV3fGu
915LhwOGK2TknxYEABMLVNE0UCfnL5s6/M9XG3RCCbCjl+J3eKzOXC/Y13JJfUYS2C9aKCKLMtNp
QExVpWuZlwrhCf09hmUttnwYofNBOEz7JY8X1DEiK7i3mZlqzQNTfk6Yy7ekCUdav7GO1k1dnfF6
PxiOHW+8xWZ57cSjldWiplyC7JxS8b4ysAjkmwY3ncalr+eVDl4GO8XHe70B17dPLEaZiMoejIQu
gQRhGQBsHNd6DDXFS+zA0Txh9q+lRwWtbGtyP10Wcb+OnA9lfDiFd3kBEaDoboQdjZmIiAc4wEkv
NuzZscpPZt0GVIRyKJTxkbPI5W56rmvHwMVADVlZTZoaeD+hPRKd7JrPZ7ar3rztFCzMS+lnMxhW
C0g564fpq6/fSU+j+9qlf08ckSVYqx+YL2LoT8sd7QEuG2DiJdJNs7ENpkuiXmUNX5qHIrYpdOW5
SiMxLxRgim9KSnVMGkQd0J5R7RfWvRlhZhVmJPs8x1Qx4zxZEwlJ9MolsJRvmkRVFWFqhiseSGMN
R6AhtBx8t3VXGRxtYJHlfCCgTdENA7pm0ZBzy8wuaiC7+0E7gIOmf27CgOvZ0QpLqkp/cx7YrfhC
fzbmazIIp59qbfUkMOPjLkPKAxpe6Hh1Gb2EUK3lw01ZLQwHxPS3Ek2yFBy+yODHmr5u7tzb+s20
5CkmZxsVXEEjfnM3denN0Ep1l4Ons7CX5MUeoUC9dVCQBv0kjrUBSLOVlmKfqQxBzEIk8HqV3Z+p
8XNxh0GZTYnYqdZA6KEWYr8APnjZG5948TxwQ18QtZqJu2LEsrmtFdytJbDSxVgQJxTNDXPodnUF
a9vQEGktgt64XOGeut9jlH0Mxs3V1LsUrRcaEhFEWxtwTkCLMgpHJwEwAeC29hjhPK8HKoT6BQ/d
+hdanQ7Wl+mXf3/bnv1qi5R7Im9vDbILWpfz9CiOgLRsLO1G1O+X4GOjuldiwx5MfsGRls3O5/iV
v4rFN2TQW3R+SRQD4rUg5A1AaPUoKh9SiIZobrliujaI8aaLIrY3dU5vKTgQCCDMc6NcxL5PzVMv
URr8ebVmx5NOV3Rn4pILfDtg8pa+hz/vvKux+1SlHOX1MWW35EAQNcCbYvqBScSur3uKHbR595Xe
tPmZtJoXmMS0JGBbBGicwcpoork1xEsB6fjy29UpMTfEOTR5/MJIyHRffRvPK987z+mgb91L/vdF
mxMAqFH0gu+ELkdHxaZ43C9Gilaq9A2CRUMeWCdLjlc325GbLUQTiWt9T1Zgvje6mvUTOxLHIYxr
h54nkaSFmsn83uvYqxOTIT3WoODVzyGGPaJUNmFptM62QxEUJWxVnaj1Kv/0flZJ0ZvFfIC07lqM
7iPYLtuXSsig/a7BoH26dyl83wiV4RbfdWqB65VoavvYS9ol552CAX/4maL5HAC59DC6Z7FlBalL
osv2dkrjnheGRdjPs19p0XBnu9Snbu/7OPz2DtAsXMsVqv4KdolatjdrnIFYIuX5KR5q+qY8TaDV
nOxmVR2voxisV1ZMWaEYd0C922xWSv25uxxRucG2X7Aa0F4Ca43wq2G+m7+rwmOolq72SZx1Cxxj
nIa1AgzfiN/RK29id3psGcNCd7ajaXijEgmY5IBh810uX5+CU6Guw7M/n+ZQ2jld62mZp5nxDi0z
RQuHZZYbAnTc0BzK7Aqov6EVWistmRX6K7veV/DvlxuFRChFuF+LivvdcVEHghHKLU3JFVF6NFcD
k51sIHkCDAs0gqHpaTuZad3g+ElbjmWR8KXt5hmxBhBv1UphtKweLa4/dZz+vws6ocp4UfK9NYRK
uV11ofPfxessIAfjFhrmcgqLV34Ji7OCGL0oj0MVSgkcFs74uqmal7XXAgb7yJcxtN6vHpRQ8nkM
ftYpokZJgsdri2UZOF4sfsH4cHaC5OEJtRdhtQH7sZCihIyO6O+tVx8X1XV+rU0jOh0vO8bzcSut
T6JoFbXuUGw6HE9p2eS2/bb5wOFDOo9Bx2LEa27Q/m10Hxo4XeyZT4H5pn6BSNgNC1VSRxVOjvgL
mOeQdqL+NQWmuojnjUHHZ6/XKSet87EOCI2MZRJm14wlFGdr8QW29NTH9C86aG8+kIdj6Shihpqi
3WIzD9b101o7BRi30zd0q/SU16dCHA7tCDeDVDe2X7L24uHrCamzUV+Q2ou3xbXx797jnE0sCJYB
mCOMxFCYpKGdaMR0lPwEuE0BIVFwmaQzfNx3qILcHGS2FUYVvv4i0UyOjCc3dJmqWhQ2sMIuOST/
EtHao9vCL2x9UEH7PC5Gd4F+6iHDgDW679SSe66fKjP1QwEiVH05vxt3KIA1zX8zslQFXalaU9px
gq4oX9vjRd79rGzDStl0Bk3zUomodJXNKFiVw0eFfLWl4QJ8eKby2TcqBPHBGS0Aa8cNhIdchyWy
A+6fTbrTxg8ljyBYBBU/QjgCoNb13pL8MbcbBXcAy7VU6OzrTIA5MbOMKNAH0KHLcFPMgLUdxMh+
LVaIjPSccocHKQ6QP94mIS67VP4BMhB8LFQoahdR8jsSgGFLMhNAKIWiuf76cLtD7b7Sf9K6xLuq
yduhjeafDQiRUznqBa4czkmxxf8djWI3dhR+P83S2vTv8Xneiv5FhN7UC6XWyi8RCaZw3dJNxkDv
vojBeDRJ4SOSNUB02aP1DQUNwGUlkGXOLa9RS3SDtB9QlsSK9dVDzwSls+sM6lKegZgVtZD5Ambl
0i5a8hFd8xSnwEXyfbeHxL81XRk57XpMW4lQv4MOOCw1fezXIkhRjvALNKHLjQ5EdjoKGLnHHFiN
5awAfjSGCtSdALgrq+1BtCrNqNHn0jhyuak5dkSYbuXukejLKRu2IilzvWeAragtGa6T6bNnxvKE
J4dvLYNJ4kgmVfkeViaxsGFnLuhE2AEOQDEXoaojS3NEiYRTl0+BiYYeAssjUt2bAxKPnZ1EYoOH
5BmvbEP/XjmhsYM8DfS01SMXjCWXvqOfUb9uTiLAdDpg6SGh24rtZjNJ2Gf0pZafk5H9uYimG/jR
6NiFPi4sssPaCKPXf6BB4LHfC5Su+yaQHV8ppFfaxSHHnm4kZUwe1bomZeB9ELBAYJkNt0DzPL09
RJrg3gMyRhkx3lY+S0l9IWDln26/c7ognhnY+nKwERZOIuTZ5nod2pRUM4uWCbd9fc6D48LECWMa
fTXg8k0BCYL5kYLYh/OHLgFIArBXefbO88n2PgAy6fBfoJ7Ni7fs7vvYDnRoqOVxzTbPN9/mavj6
tt/KmgpbUa1K86MJHIRkgiXDWMKiOdDdqnACubaVezGXvgwN/TFYjGoTmwYFmlFhjz+OCPJxal7Q
1cJMk7xuG7ml9njSMUp6Fa/nfrdRseIiy3BjSHBd2uaWASFkQt8G781e0Fsm5Wop5fbYS9wvrGKK
62hlC2kkIzKvy1z29B7YpLytiZznn/2pMCC8wpFky5t+pO9xswU44j2JrpJpUd3xUbOTcBUqgCHK
PSMqo5QKz2UD0CHxJFC/CkZG9cjbwgLypZRcCaHYKvhEdhzXsHxa6ImWWWRFWr+nJe+BmJVWItSO
Tbxy3CrUG2+JYFFvnyTJhhZXB7UIy8nsRXbRJ7eg4s3jukTn0AWM2PDehUuhuHQ5MbWa39XjSN3Y
K8ci8gzZnPHuNUbNOPGGvmLr1Q7HEKxXTYjk/2odZE26uHzHeeZxwt7B+mKxM9cKchVzWCmUCAA8
jZmt0X9Ko2+NFi/R8YjSobLGePRJM/A9IPwwN3kwDaVrpDD02R3ZzAKUbkHbCyHl2TwOYXYauQIs
u8TLGbZyHP7Q6hhhmQc1Qej6EIXy1odffpjqQcFCED1y0moAor6j26bgQsGb5jCTtooInoyDgtYL
jZaoa8NKN53r0k/vgr/VvvzPIfrXC7m5GiR3sp6pWlDkY8f/hnYuucw+U7lGgH9hCXWvrkc+NoT7
gtMdDgCH34w6Ku6jEEM92QWvVCx+XaYBVcswhwMzfyipL2pN9HpbXSlW2G2XwUE1Tp+Z3oEMzRAJ
12/wPQbJOxQjg4WfepfIp2zD9L8abLegDdvcbjDMPMQSNLvXS01jBanZePT3zGRWihCPCFjqQw8T
fOBjdkdkglfmzNHXGKAg7d92RuTk6Udhd1G+7zct1BMuiDwg0YeLIjHRZn7f6+aeNQEy3Zy1enVg
wdnGjQXDALB4br16PpGG+nd5JgHQKN8HZj1aAxWB3HWnUkeDFqENkGdPbitEfolO64lYEY7bp4qO
G0nWSpkv1ywxPy8UGd45f0bhAp/OeXRpaa7ax1AUYQ2Vv07HiXEKAYLys69QQgBhro2ZH2+dtqom
iFmuC4PvFDLB1r7Iz1eoFH1jORJqrDgwPHD5nC4e7V9fkA2nHOuHgSx/J6fxCAisHEU3slbisB5o
f71hlibbisi53NrQqrLJDkhWP0zVOgc8dYjyqHegTNnRGAGht7LvYtcu/Ogzc6YvC7lodQS2ITBP
trdiRVRV7po5UyTmTEGpZF+YVxMe4O8C2qgDtkL0etN5Tl/c5Ly1pOeq1pdKfjn5slpyhlzGkYph
ILvO/ftDYHbX86IAMc7zhNHF45CBcF3Km0ILIa0Yk+tARDWCWYU5Gw9ICcqZ8u1OAIyvREZP2QEC
nobjepiKQVGqfShcTIOeP8czQArOlKUutZokuhPTdiiLreE/h9TwuqvgvBpi2LZS+9d5rW2VM2Xn
18gFGbx4C/W9h29Y3d0qGzNztVt1hnc2o8Bt13fIQ5IMvxJvu81dIuHVoqSLlctCRvUCsVTulobU
0nEOkWGEQ0QmBupfT1S2gaGK7Cbs8rTfNzY+j+QcHqCT+ZXEmhvs7yyCHfWmAHMlcTyE2ejLpIQ5
0cGEdgm29oX6lEvxksXcpyVg5P94nEv+glMZS3FVAdqwxGP6twQjErLWzd5NT6Eg7AL3frh0Pre4
zhJ2v6Yn16JPdSoU5nBx26yco2ydpczRCnvw8OZTz/Ou/G11V2R6pFVMMi49yeXEJvf4rXi82499
cUn7PNVYA1GW1etTrukyZSkaU55MC2KhVMEfVxTz3hQHaM6pabzLSO/Cj8ouCxcmNICpaUjmlwz2
c/nTer/CMuHnIfkejfNwodhuWMhT1JE6m+bHUJGywYmbGzph4EeYYMR/2LsHsm9SWqBK5OtKNWN3
lSOK7abAMEys1/IiaeAk67WuiBMfixbtI0HXKEcjcaze/ce2IzoFMPt2rHTYF1c8NcwKARDjmK3t
teK0lEI96TESqof6usVaFed1PefrR45mbXnh/qepgiUgCSQ7NG+N5rwfGfCsQZKViYMsQiz6vCJ6
z8jenP8Q1RCU/PhdK3enOwSTVZ4Ke41FPiV0tTQuSQ5leloi//mRXj05UN4pLt21L48KVkiUTJGQ
hfurGl7kSMcFI9Mf9oeS0PJ8ZLQHp5nCmXYP/ATq+5/nl1nIUzLySSzrv2TG+HdVrd/iwWHULRTz
dpa7tadlAoCgtdzGfxlxAhfrYBODGF0wChdiqSFiRjgvib02CF2h382mscgCsNi5ubUEX7050RmX
0CnO2JRH5wt3etRIAzrd1BYlu9hMEdbVoec45EpIIGZf843pkRx6WnoAKf6JALhpaMuXba1XJMuI
ezvCm7TYtDvyBu6NPTJQu9RB98wU85ABKOryrpAGCnX06KsPw2cijv8g0Aa8mDdjaj5wRBNhWNnf
x0J4/Bm7SH4xOyGmf8PqJDPE1M6hhoSJzUIX3TY=
`protect end_protected
