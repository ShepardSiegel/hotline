`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ml1ERECJFmI0UydwqCNd4t9ze2pCKaT/YWzSLW/JYvN3IBo4Oet7wvvrjXT/Hg0h6cBJ5GlECJy+
cPO7LhN0tA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SnaoSWx+5k543SXKxeGnkDcu2Xpw2ILDXZq9iYLYnZsbjGkgPSOG6gGPxPl8M6Iln1RPg47kuBNs
nEERJfUvffBatWdKQEQxiLJjSZaU+pf4SwTbWMuhb2LKP0WX5HPPjJtRzakR+NEXZYgYXHcQZ+Se
7kR5VzhgyueRQEZ3RSQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S6Qxgsg0by8LxlgUbzbSYW3N3L7m3WEyI7f/dd3qouaAHZWpYA608ZZHAN4x4HgbTIWujVVn3ZWW
IO3Sy37mNl1KOZOP9Mxw+6e+RXEXIm2abV8DPIkHHD1duTg/kcK616AvwtpazOxWBE3MdcN2ZOr0
OG1vQT/IYApF0TXDdHwjKW53Lu3wTSEsdfPhzfK9oHx2HCMQsHPEu84zhpxkNUJQhnrTL0nqL6bm
iTP2m8IbK6leQYwJq1XbdFjd0A51MLtC5PwV6HizxVl2ui8Ltit9fTKhFhxkDigql3tjzrifKWEG
dcoEf8mv9lwBMyf58/MROk5IksqjoSjJAsTwNg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DmGwn8T3qKb2uYESL33L13hf0NvaA47HkbfygLRmCiFh1tUuTqa+gg18Fp01sVqYiA/Dhzczvp6+
Z8nG+i9jZ0qzwcN72N84RgYqh8GqN+Z/YKJ2kqyj8vMJMGwv1lTn8gq3nYAC8mXQ6GL1ectzyExx
5sgcOWP/5SqwLJD5/oQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XyKhUDcPx2pzpxbp/uxIUWPBtbrIeZ32dQi6sWb834lniqMgn/euhbmbrSyS3sqvoXOTZEG872qX
22OOX1ete6vH3OY0Ixv+bfiQtRCeoSV5Dk8NI7WVPeCR2Nq8GAEDabhTjmBQASbUtD/oX7YVrsg3
aNV3Js8aJVtrF4iWlR9AxLtOdJ38Give2B74D3Xt489uHeDizMD3u6quZkpnVTN0GbKnEW2bauOT
6r4q8Y12uVIE+2//lazDk2s+NFXOiuWDTOZ1DT2TDhZ/hz2WP/ATvEZYz5C7Pq2lyUhIW9R7ZKmu
gS68o9CneSSxeGqXDSnooUm/LKqCwStHAsiFVw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9408)
`protect data_block
EYXjaxF5kE4VMQvUm1kiubYvy1Ohx6OU08lxnriD/dAwUkneqaT5YpZD55koO4L+RsQejqp4CDdL
b9z4r3cxAqPp3g0qf+X5pZ3pJfF6sksQZvINlthIjS1WW1p0ZWldaemy5famfVNvcueq5RqFOtzC
8VLtpGABcBx2p+whmGGqDZxDHU3+R+nDGA7WECmnqPbnCgC+vnz7I3pnyYGiGWpWozJaJWC0GS2v
3786WpKP+FsrICV2iA56FHGio6jff5n90ONyCr9cTwgXO9aw6ZXgawAh75+xzwnXi1Jha9SA9oIA
ljGWE+IZQcMPiOr69AJaebYXaY6dHF3Byi2kzu1h7ccO7RqGz/M5YAAoIcouhDRRoGo22T51l5le
8Vt9gl5htcCC1/UCQPGBFN/iDGjl1h/m93oH2tt94hY4gFptlcR1S3jOqgDQGP8503QOdJalGeWS
s7DZysXC4EVOi5KLyhlPcK3ebpPyYhzfvkUbseyR349Vzwt7z+sMBh4sjCvLQpHPZN6QVlsTAwTb
I3b0N3n0vmmExIivl9dgZp1Y4LHAXBmqojdcqi8xVJ+fLK3dmTki0s2EUjPMpGEop+ayI8ZsUKX8
gutuhNKfEtzPlBjQ8fiVQ/6qWnHhlbY0rfJEO/mZ/Znbu4haUAOAoMt/JCZDyRYvtPtiZMhNY4Dh
NojLUDZ+XUN9WOf25nayE+0dTiLXbZDTF37sHjDlY/bs89OH+BKDm8A8d17kmVRdQRFT/KD/+11e
G84DPAvhzr52xt2gMrWGQ5J8/kbFyOAFm0HuYB/a6ic9ZD9BUkgrRwO0bv23A+tsqtrLVItpZ8KA
F5OhWPRO6ltB0WHiOd3V5LoPX5ePMWPU0l2mUUmdBeaooA5jNzg0EVhx6rNI9DaEGkBKyy0/NU7R
O240epfctolICDLb4Q1OTBHkViG21xSsAM5m3v6ocjDP/LiSwA5SdiWFhDYx88nDTOAZuPFpFDch
IfgKBpX7WcURXHy6POFdZKhn1g2ss0JuCtquO7Qkq1de+HnDRy1lzQiNjKinqm7B+svSSLOlfEMG
1cmA9Jj7xJ+R9X60rwibfL5anWlDZU0gy5N5pgH3FQg2qKVscoWrhR0TdIX9YcxrBdYPCoPmKvFL
AEwDLTSfVJaT65pOL9W1Xu2CPS23BMy8F5ODVfE84htuV3xqOeDKa2zR5EcmWCcNf04IlprFYCVb
7+sEYDDD8eS5g4K74rkwRKmOf6DhnHuvYAz7+uDIrBtBPCzWvSv1WfWCErZBgECx29NRvcSqBCVC
l/6/A0B+B106BJZAbKcBWHjSNHopXJfku14gBBRmCARVIK7xCAMECD8PP4uy5DGl6XvICD/OGiW4
TuR9iXjcOzfZiXOh+N/zxcBZMNZap3559uYLFjOxlLqpbiN+GR5nBrRUzLv+XmZW8BSWa1cnNcmd
W8Erkf5+1CVn266bFYR6Q0wEapFtd0fBFpNGjPm8AIItaDDVuUd8BunVFWCbh/McRFbrNDWmhPNC
CbtzUshwSFSq3Hkr5u7vSKm/KZIulOSTrHlok0bGcgZ30f0Y6+RWZqEaSTn02KR96mSexLef0c5i
Rx6qoqBAZejNzaQIfuuu1aWx9MyqSiQ7lWrYBgIHKAgpE+Iw9ctIpNMzCRClAd8ICaylPeOG/WFj
DrvKmbTIkwqfvqZsA/8hy4N2Jo7WwAoCH2OR2JrFdWOPLuYOoxONESfrNJj8IlaTt6FZxHM1dXDw
DH75biR18+PwLUhBKMHAb80iqiuXyWrAKmpV6eEVeA0d8QU7OEY8H9eKaitQ5VygwH2PbQHxK96t
WLp9iakwwhmD+aHsSZEKYMnDhyKrBWnVJ3v/EmiP5GtY1IillJGfZSbJqgyy3pKvpzWp49aXyUin
Tz384Mv7K4hOMBNeGqn2InQ6NFIYjyT/Hx1hl50ItoYC7QoYh70PCWDJHyiHLqKzo9r0CSfTMhsp
mVTomtP0AaquUSqm7kqVArtlh/4IkbetpPvh0mZbmqc8QDJCnH4FLXv6iL1AlHPg9olEs42B4T0R
NEuyfEBVDAYUNEsR56FGdBGj0zh3i+Tzqo4+LMDDGhtMEGJW+sOlxDKYREn3m/NO5VVnW/+G12hj
ebOz32uSvVadiYqfXsZjBXfcMhWcuxleSRa/UyGM5ud9hVsXylXc8xj/udUsbezsrK1SDi+OlN5g
P+OAPg2figCM2jiW5X1twCZhXEhcfxzIUKjvZWPgHaW+LtKuTWKY04hpEQXqgF0N1KFOBVqdTGX1
kwBxQdjetd2bFFySeNW3+K828pp7VFiIU73xAj/evkJxCc/8Pl4LIVSseRZuTXxc4Q9/Kb8lqd/d
BED3au/FcA000eKNR3cZbPmURW3lrmo633HG6nUTpvIpufWgI/4X22EUpahvha3103wlLST2xlak
mKimY8Gq4kOaBSLdstOxAV2/Qd1cHnNRY6bv8e1byOGOwhv9MmQGgYmVJT4/IGpS0T8SUtyzVcw0
xrRZxpqHuuHjo5favF0ep4XCFxfNzk6nOb1IckMf8qQiLA+TL95qlJLcHeBFA4ZVynbFHUgZz97q
erDK5p8g8WWYSMl4oC3aCjLduxhcUqCAO+lknF7rbFXiH27hr444WlkYWRRhwEwIq52nVGb6VBwp
N1BeTKKKhElT9q9MGqqFo0ncPj+xiCeUoYVkA/nTE903Wp/0VriqWg3VevS18T9slZ4psGjZ9Ws7
D3iLUBp/7aRwflf2NXQlP2c5iwMR9Aa2SPAUjj8F3d+IpdimRHInftENbioM3vRScgHGJAM31u/j
tXk7YUj4Is7wKkZu4BW88FmPCAEPJ2l7w2+NnihMqg8ZCWVVQVWVGFTuEukck88EYIjCQueQnWEP
fVfaRArZCIPYQHP/6cDB5toB0eXTAON4eKIymIpsJVWYC/ah0v2vYaRlUdsCvY0HB7tjqiBB3x2r
S7oga6Z/ATFx3hzjSeP01UknWOlMb589u10vedB9IMCwnLHw7qAX7S1ybJOEtfrGjvy02QHjyoa/
qstXq5XcE8qtz/3tdkPQ2OIWJHp+cy7YgS7V3iziIr+evatsCG8ciDCkBaTGztNFNmtdA91vrxKk
YIc19IetF5j83EmwJ61BxMfK4x84GDzLJ/wHZr1C0CRj9ve8ZL7GSGPFA3CqqxbvP14qIM95HjdI
dhftozIgm69cnzmaUOXiVf9THuWSamWYo+x2XQ7rLh9wYY0C+lqga4KtmPT2InR7ONEqs1omSA/7
qTXiyXaW685wHYdl1amHNQXQJOsbQDnFNs3lGd6HMOv+gPkALyFxButyfaffT0YRgoqlMMGQ5puH
uNjSIAHoUMKUfVL+49vRYZyJqjRCEtoIuPWWslJhFQuBaU4le0JsRLb2elQuUuUEA8/Y41zV6sy/
braQtaFu6m77GaLEaxy8UaMpspPFgAMoRjKd+ym9gOnNuLu0pX+d7WgQV32fuB/uOt9U4ACZ5Cx7
AI/Hk4QLF3jQ/y4t9/7jlTY/WI6TUjxcT59QTH+YTi+bdnxyRrAZ2pE/Nd4bwr18Lsue9R1Mceed
alG8xr7cJcpDXqa7FsOmfqHjpMJt+625lwSuxcam/6/4mWSj2B0Grhe4eDsLe9T61mHUtCsdvZRe
xNtyizpDhhkWy7OITbzuHt45JrYLXlxNq6gBNtd5bI5TDJ+yifa/y+mEJTC1Por2PM8M0SwckkG3
ZGcSEEAewpejq2yGVHMMXvXqWe45k4ETk98MZjs7nVhroKvKoINl0QbxBYwzm5G/E7n84a/Bhwdp
4rti7g5MqX9+Nd/3pBt0wR8zA5K+3qIVdopygkR2z3ZGOUvLEzMf9yVIVyS06l1sB35mk2VzW4DA
ZJzQ8EM/1xMk8jayE03HBWabtud/04/f5ofK7a93nSxLBGknxIaVVMAOObSKGPxCRIvoeOTA/JGB
+7MRuLZRmcEODxf7lGZFwV9DAR800Ez0HxGvdW7Ypg6zBaBcoFzArhU/WhHTYy2WpkL5fsdxy4sE
W3eSlWU1y9TZvKHmNuX1ApxhgVIgyQ4uAKCgON11FA+1xdDR4rAJEWO983eJ02GOEbpMuXfkGx3E
nGiVtpQ+An69tw+nehGtrDlH5qFHWgu8zI2QoECJMVj5Xgbf+jOLwvVlEbwp6CinnUVuH7oVx0sR
izPZBb3qghEUu/8FXNINHRM0NOyed0Kyg5wnhsFicMj2g6Hq5SntRKbJnJtlJxtWfWziBZJjMJ70
aA8Kpddwc91wgH/6JcTEVFW1MZy4x/p6JEpmFLbJxf6gLLho9xn4xmepZgmW7cEvqCOlK4buIgI/
FBZaAkjUhUE824YoG/Cdy3tOybROGdQXITpzCJr9hdsO3YAWzOXPgYLLh02KEtnjZFULOA2oT+cl
4nzduSx/43uFnoghQUapIb4oLx8FR4umUMguAR1wUGcKnzS3d/X/viydnE4oQaR/m1ajiCLfQhGq
/Q0uNVk13QmjQBAhzk7u/xC21OJVOFX0GZbQudUL6QMo1gF+b5IJ1IBTIXWOl/xKkBwxLXOWAJIE
I8H+XqhGFnmJtrWq244Y8vHJlnX4f+OVn4KPm8ubbHXShqdLUDvHowTlWBuCTN48KiI7RpNGa+7D
Xek05l/2/e1oNCe02frGXliIWyH2zdRLuQIehl8d74MX7MqexWe/w/ofdsHWwdf+m7wPiD/Ebhfx
7M1eQsEsfwpsRguKgCHyPNAgyrvYj9TWJEhZ5Nr37QBAPuF5sZAX/FMPrlh3nZepfBgyY25oI+6R
6lLbr1BxyzaA5jzo8qniQQFR12fQpF/Cw0pKNlj7loO7AG538JkXwI22dzpjv+pCm8sdwNxfPB3Z
45e7BZ94dk/L7PE1y759O9H4kdGmV4lgbea53NJV9Xk4SXmtdxuZV2mtD5nN4ty673fieOPmoCV7
oZd/rRdg4iDulrYla5vFJINMp/h2zCoeJoKa/h6FPQiNv02qyZb1TiEzDhT3o0z0rh3eEpJAmSCx
xWS6JOqW9tv05La73/TENv1J1f7qQ2AXUzFIyp7jllvNZsuCjyUH+r4TJH1oj/VnopBUMzUVU3K7
G+sMLaruMUJMMJgb97oLgw6un+D2VaHBrNFmTO0y76mKMpxUQSiqxef7TNOY9gYPNhaBEykxc8Ro
CsyKd/oSvbbLwDxTYmK9VuKQ47fbffJudGFN0WxFCpJ97dmjwLZ7IOGqr2kFtKxwiVOIyKTzKqwm
KRv6V9Ow0BEIMo09YNLSDs48wnBvr94JR8c1KZ64MjtNv4BcO2872V/2WMAYzS4tY8Dxjxrj36VS
n/RBxJueWaueGgwluM+KB1AzJZjp/F+QlwZoQDlt2gq1QMolE/jEU77ypaLcE049367L1DOyptLF
+vE2FugyVKT14In0RDMF7bh5Xe4sZ00PhTjamZAqbvHh9LeqyBhIYQv3WFIuQxMEvV+07qQbCtXT
XXpCHSCY2IBeCoYpL91pkXJ15i2cg0NzS59zA+pTGAED6qSTGTJnrB83E3+uN3uYC6KMgoXPb6Hz
qd3LJ1x1dGdjhTJy5qKKgVdLfEgt33XMUyqVzHMMsEaeXfMUsMRaYUo0kW4KiIH7mJbwAFYzgFAj
ScYfVqufraTJmsjVDiK6qdDDHFFXnK6vbepTHJRKbBYk6n/4oC9yh8ScnYv9js8Gq+W7vMeQvUYF
3TRjU22znOz8TorsWoUmxhcwTAn5ZzjlNBq08EfvDDAlwGtCZpvOqWcoZxtZ/hMmLJBmADx9ePFn
xWsfzwzWjjzEktxfpKdO8oYfSQFMUwvab0EwJmGJwgTQcVh7ZZrlT4kvtmL450pKqcLbrBn+TQuh
sc1hreRUSIcg6V5N5K763MlMv9f+F0eLOLvTaTKl9AJP5hSHCDPI/E7E0t4SNw5kSekDdrUTMb83
Z6PNNjbvkfrrdtjfuiJjwPhBzSL6YfcxD8V34JFeDAsKEYYv5APdo4YI4KZRLFVYVmzAmn7U2SeS
9SloNEsP4maeIC1Mhd7ZLIwu3xWJJg9iGAdz1YvARtLXNJu6/xlgyRvdC+TQh2ZRZOxt+/dQRGr3
SI5YTXfV+URe+RA5GPQ6gkXJjfbuIySImcIMJsVHElM9/GS5fIUbYyDqVRbalo9etF7zsOKgr4Ye
04QWb+dCUX1s5ySqUx65qpFUiX3kfqQjECT9oPdKNeS1RAxFYU7c9tKkXmjcvpzPpceqO3PwScj7
aRcfCPGBlZrgygkbCNdBPYOmWrNsphTetJ9pwKQsBSnpvZ8xq5zhduSYHeCxQ69vTi3xr6Ir/YC0
HAUdJOE4A7QRMpMniooaOaBxx5JBSsufKrYTsPevsMeP+ZS7FOlrH21uOFpFqLIYGba/r/dw73Qj
oewJD1XZiHU0v0SB7PiqRXzJnsD7icTVgEGQWfdFr46wAJmynU3z3Y4+UZnC3i1CbLw//tRsI0RF
3Hwu4FtMl8HbROCiWcV0AlLSxrkTdgxDTNBn7rln36VRMCIAfupMh7GyUXA8jtqMkouVz8bOtXZe
Nlq0VY7AV7gATtDIgKsZaPfpCYHIauquYUdBv7erPUgzsut6BVVvxP/TB0iFX0lxaPqdNYQ3Gpa6
SfqW5QwfCrp9Ii3Bvcu5p5U4VZb6v6oa8ujm6LGfXU7Ue3BRZ1q/uM6DpwDCwq+1lChTDn/gYZMa
qgLPUwnVEZCYCDAOP7K6hIYhLoFp+ldRfOni9v11DDnkdeDt4gAb6EFxRRpL3tbo74nRLwrSxpRJ
2Li7NyxccOXeAavVoT6kFONY4nRQ3oeFMY4UmgER7rJSh7G6NgYnndprl7OrumIORRlDoaclee1G
IUYThYw+wh+bR22+4IcEPTZkJF4kulqgy2HTOldHAj7lYo3E+DDFydP+RZF1t66dr1Sl5uJyieWk
PaR1qvEMcdlJDL5Pv4/O+5NR16NO5E+ysD+xfcowHq24gsTZC6SscAnmbNFIGpoEN+lbIyURqvS0
9crVBlh258FxzBq9hfywxvvo6Vc8+1P0VrSIbBc33SmuMwuX9xcFai1e34D+Q87X8839Lg5QOWRU
nRFAb3VMQMOmiF7jCi1xnJI3q9/8eL/UZOXsagiGzrVfQPNVHrxeKqIpTz0Z9HA8Lh49Q0yCqs/W
JCZqcQIex5NvMfJcMgUEA8u46wMQOmfJ/TtDIfYta9f9KUQRpSdg2PevioQQotJo8H7JYTBrQ172
aHx2U+q9JVQSOJMtn4AwnHKK6Jdj3JKRjBkm8+9Csp1Z4igE3h2MT+mM9Lpqolij0CVS9YWPtYXC
ppRQBvZHjDLq4ktunmDXxOfiEk6fqGvLA+ULRRo+z5SZGtT28kJGyZqlNAbcG57sDzy7PE1hVy9o
mbhgOe2kHTilMlRd4cu/uLzNMdsFUNtTGdMPfgPbz6YQsTaJRfL29lXgP2auOP8KDyP8k+zBPmb+
iMSJmY62DRZWDlO2fjD2GyvxQzYePTyE3jJCeDKFM8mWd5/sKIdZvU7UAXxPkYWf3/8sMgr9DTRU
WjRsrZNFek2i6BtXwut/pw5EhwB6UlkOvT57k+h4bjuTI5vCsxmJOz6sCrpJyt+q8ID8xBcy3QFZ
+QFtG7ezZBQt+hwBE4O/hHvrR+A1+5C2GsE6GVBCoL9urveKHhULXw8fcueKoq9W8kjqe2/ImNmz
muBVwTSrhI5Hu+6bANAC4jg/4UBJF0joZC3HhdclDa4KeRWxrpU4IbZSQwYVYMalbV2WqDlHhz/G
0xt0qKzCfz6dP9W7HD1jEfky7sYQSYVGPni0vqaVlICwms3wXXnBESJNfRnaKFzI0hdywAoqv01l
q70hBMDosuoRm5ycRBobMbZEYTDIaOlfw70fjl6w4BrqEEWBsQTdQOx9dzHpg6yY76cPWmKDfglA
VexFUl4+WK7hSPZhzQF7d48UquQkHjwuNLFIluwl6aloTARPZx+v2wUTBVlhY8ykRRNWIi+7Vonr
VtQnkuiTUQBNcazeNo6My+itK5yEJS2prK6dFldzU+kDKenLgGGkWaHsYfsUj7Ys6B5++KsyADmi
q7zDT3+H0z6gx45JGXXeX6vVxnbqeXP3W5EPnjdbEuESFuO9WptKolkS+Xi8bba6GGXLnBZdltc9
8CXydLdfGT748OuzkOEaT+0BZkHYzKoOktziIAKV3ISXF7vF4Kz7a+xcXlr6CRArp6/rerx3y7j3
wz5KFeyXpy/cXMnqq6WZR1IvldPrPVSshYGrtx11b1Nd61L/+XLS3qh+SruTn25bhCslGhR+U/No
IgcvHeZpil5VxL7pftG6iWjtSGHb1wRo0FBqoSGJkzZjXKQL4eeyDvyKfnh3VFVJRxMVhzyyzSxN
Hq1+mKgK82M75eAwoGla4lOqWWwuDBAXrJq3aX0mGtTVG2CquauD9nmGCgVqA1KPtysagsYa1w3w
jolWiBzqcK0A6tXZtGMD2+ANIrqOiyST1DSMSIhRmaF4lfIPGA+/H70BDiPf3MzpBmfu5yZFoJWV
o2bxVwEjpIG6V94Ovsn55B7/hoJgeP04PYqTS7GGsaOkf48QgbyK6VPuPYOFkrTsrm9cRgxP85a2
SGYEqwIwzjyjXCjZDbjBiXPlXzOYGvoVEQwVIQZpZjPJ+oKIFC/kLLotBDnRbNBWpYU9khmwfprJ
PPgxX7O6kqQJbZqyYqa6VDY4ZocRt2XMFUCH63JoS/Xh0AS8pbjcaJ3OdPE4PKW1J5scRo4n6sXH
rXz2q9hORwGKI2XrT7z57Mvk2/lyGMaHIBXGmVJ+PfiGBFaYDNqpm/+FhYTqVN+my5CGs4ifJoZp
sL0G7AsvKNizbZ0X8ih+5RVDyrbkGllDHeT60JGXnB3YPMd5IXi8F5wjMp3LO5TnEY1YcbsEeHdj
o/YvM0ThlT7mRAQDsi4MhanomXbmc7y1ydTKBsblv4Pw/YnJaawedn5Ej5RfkJtV9GepeRBwhtgM
IL/1Qx7URtl5X5c8olz3ALkff/+yscHxeuacl6VXRkKTI1PD02iVBYZA0jJu2mILuzdiK1UBQ7kJ
fMuXCKTZgacTiyrj1nGotlkppYaBs4ttkWqE+3gfZxUz3gNmTs4h5Ga9USJIM4lZQQYIHMRzqt+f
BTwEJO8/KLX9FwJZAE7WtamtHp0zDByh0tGUg7PJCFNxH5QPCTz/Qw6gG61m2o83odIFKYg+YB9A
X3brT90xn/wTV1nNii57TWIXyIEqG7rZw7X44o+adrMZC5S/ByJFQsrK874HwoqtB98qvMu7Nd8R
c6vJ3Nn1YpIyV2JD9G4I/3kfZ/i/omYVXRK6Efjf4I5iukTXaLRG6wVlry5Pr1Jwa0MeEvDvYC0V
IS3e3X73aV4taoQB/+F9F9K0L9w1WecFvtFi+oj4pHG5S0GOlWoVEUvFVjK2yx3BD0A/HQ2GNyXP
bmkkR0BfMSiskTIybpJ2Ss1NZ60rnQ148nEIlrhkaCAIDPwpv4yc27taBXmumn/rzLmfof1jo64w
1NisAtgLxeyzDCgXbiZMpRIUfh/fXdDuZPktCgGtIu/n109TG4wY41Mjf0DDPEfqieRTIXW5PIPr
N+H5YyoDUjRP4MC279GmvsrI6upMJVDSaQYMmu6pupy5yjamRa9T0SL9fHkBjXbyFu2Vvmiu+oa8
Uw1YojPs2v65l4Oi+ArYbY5ymoIomJPhMWz6K+I2jcmrlGLGJzk7C9JM/t9x6lROw0bqniZADN4D
FB3izbEnKoSTYCnFBGpCEiIjZpNjvUoBiD79YAUfMB8R2w9WEC0WfYCEby2cDb5UXiUTqmpq4JOz
+oUsxBkJzeiJ8NJh3xsimo1MEtdvxKOiZvfV3qtuBMm0yYCQJSOsjiCq5w09cZx77p1qyHhJN5zl
2YjsiMMwJjyw6uXjlnC6dQufmqqGccggRRnhahFv5ICu1WRcPeg30W94gPGTqLbHVVmXEJWdAGmh
Is0FUrvM3JSg3n3yPtXGj5frZXVfUkjATpOYHvfFL+XxvHsYAEdLBztZNPkn2NSVp+ejfsPAe0Gt
0kDuHrWYSHNAuYwyVbT5Wrr6ZOnPOHaT9epaLh6jgFxGLKIsbyfMuzTQ3dqVueLQJkRdfVA40gRO
M9200MR5MKaLiYXK7l0nrVNK0oVVOW11/c2qA2hDGbOnwrGf0fggUCNmaI+JPkntMDfQ5qsEfWQH
K5xI3F7FqT9ZxH5SUpzzlw7RNYJhLVwL0Dxj1/uR7ieUR8jaa9O9HYV/nKWWR4BxmUfVpqbG6HFQ
cBm6KyTuUd6Wy+YYkdBA99EpeP5MdfCMPcF+jKazydanD82/flAWViv/H1Jdk44pfR+/arX7ziVn
dA90Yek4m8ggVd0dTk72kaBY5XhGPi0fcnbPIXgUVeGekuofGUfup5aGVHes8FEM9mIdXT3HTzQ6
7WAn/UTOETCGMsOYa/B2VKY5wcbM4CFklum+rw1G2NTC00hnsvBo24edG5kUjRQ8siYQ+F/gPYXF
KTNBpCXplXar129DZzBvyVyi2jxvlqM+AghGg6rEPicf22flKS7VIny7gS+AjF92UX/Qi6MedWZb
cImsBX5J5UrbD2lf7VFehZUxETbobtPPSUhchVQaBLPxnM1BGw7p1mFF9yxNuKDkpVgdIBsFjFqs
rDGVJleDvsr8dp2XPsANqmMRLAxUfpgD0yZQfPKdo108QiHQYiKLih7yne964Ab7QI5VgQH2s1Fv
Np0yKjlyi8xFTSFOg9ah1A7xTYN2IbZMLY0K11rM2cQM6FaMYHy6hv8U4fPvKFGIeAPDxwoRwDaY
KkanZVpa2GwJ39zHHNxKr1x3F8GBaJtkh4Di/r1kyFSStDp6r/UVS52CITIjKbpuavUxWDHQbstY
ULG8/2sawSLQMj3s8OkeR/DUEzVu469qBDE19XF8+jFaLM3mFiN8Wc13Nn2PqwBHlgNVYeSwSaUZ
AHHyBESOE39u99/AMImRqWBSlcLvlX9O5fLKJm3CEKnc0VGRclnOktsJgH8Q54HerLdTRfmCNm2T
vAKb7NdlcRumgj2kW8R4hfFVTYkkadxpFNxfeKdZ6HtglgYCdogdbFpsOY+SmgG3jiYsoJw1NSM2
vmjveuLohUCKBGG9sQhTnxOXj+aAlPG4+YFCXkMs4iplKNYSsQ/Kil6a2fAMBnL6zassFTk83anh
DFbo7BCxaQW+z/2XGh54fm+MCN+l32/6V10n0Whp7GDX5ZLCc2MFdlyAV9NukhEVcaqOwzMTqx3e
KRK4NhNJrLJDdsYG8dD0Fyoh4vRLGIEMuFM+OdqCq6vtK0iOT9NKjc+d1I8cl9g92WkLGvnPmoLJ
uKuasBSv0A8w+EDyb24BsVdZUWkJEhRIg9LBMbvSfnWkwA39w+WVDjjENf2360GzMT3LpxU3SAVQ
R2OZsuskvIjIA4qi4A1PoJBK6ij3TqlYEIWXAPC4y8iXKPZ9GnmcRqGDOtVx3DWWxzrJYKBGfXFW
a/l5N+Vr++rAnIWisIz1p+zK7EbQSW6Bh0RpKnZrLTfpjUYQIce+wrGQW93Q5Atacurl1ueHgp+z
TdQ+Um6uD4zllTXZ8+bkSemrpssIRnuHIKFIOHiq8vGGY1zczihAMKNgE4qDX44bvGpf62MfSJuS
bNrALyNe0xdndD60XMjkqCDuenrOOHd7x5QIFdGdpQiVD097mcUhxLYercoF23bPqkXNQDSJbKGJ
fUiRG+oCCugNzjvGGeZqlg2jaoDKgALGtcj/3ui8yebt2sM5z5xWK/DRyIEsaSXJ7MGlHg7n27tL
OYZFrbH1Bh0xGWXZ2uOpk6zUWrVniE0q0UPa4xDErBDraT3Jb9s//wI08FkePnPOcW49AVkPMCDj
FMNbrl+fxffMvJRzpmoNX8z2ZMroQpAgyiH141ERNHy/X4LH4dQAZqhaLsHcTN+0ZXiAdHKgrFcX
+zSP5g3TZpKK+PTXs+QH7zcK7TgE0umcRbLwXXztW2b93yhR7N6+SmKkIL/BmuhMM7Y7Suk8MW3c
ay63c1dPRkSp9pPBtsx0ynXvdBBSTkmRp5SVJcHBEfVKdkusXelKmtVGiRq2cPXMqr761SP/DtHh
YRRVQcaIz8IcMptjq02iYnhb4CQ3aun9lhSx5sUs0aA+z+kYrxG1bzzumHDZFaU3DaY6O6JmQmQ9
hLPhUnwC38a6GgVRBzo/vMR2IFZTb8dLDPwH7nYqVQpjhUVh5eFW3Jt2PoxEZRO7eeQyrYAHCuz1
7T4QfcucU1eV+BMMfMg9AselYEhYH6fkvvT5iKJxwby3KXxPEje+9UbiiqouKW6ZQEUDcqF4zq1h
sQ3ruwVILo2da7YfYnXpJ666YDHaMs8acXSMLQRFDS/U98FeNZ3aC0rZvZPdHY3Vg7BTQ+9WocqI
7tIggY8Ool1vcH9tvEIW5ZfQujESh5grmv6HrAOyuIknGBnnKJqYtAlHUAswZWYJL8+AOwP4aGY0
NkjNswbr3IEM3G2aFZTauYsaPf573J5bwJKHUqcFloqaEA84p1sSJUsXyv3ba+JQ4ZRoqGZ3xdrx
5DPa
`protect end_protected
