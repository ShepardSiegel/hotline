`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Xe/zZgJvinnQrXGMEz6X3X01VOPBV++wdCDjb+eBTUzJRDHT1eoS/MlFggYKHB6uQUQi5mCN0gVO
OSo5+UObfA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
osgFiTds9fq+FHQtY9wsn7BpDIJayUymZbmUtmHH590RTivbJ1Oh9qC9JabDsZ6GQu01fj6W7ydp
Rs0SVy88QZ7jJSpdLJ6YQMqu17XaKi9dImfyo04frbi12ff2kUAFvY5+4sBsvpLN3XtzMUZk7mPs
AUJT+eObeI0OOFj55cI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
klWJwZFug7pNpREpHmNXqCvcH9+yabPJtsCozt6wztmnbt4x6Qm9y73NKNOXuy3fpQy61kNXdppc
G/VEPCwvDdWroOKcmLncZvr4XqXVQQDyiUxRqXyIAHWUEArryIeP9zjKOG4HANf9cdMq8bc9NnBq
iIERWtF/CPQ6PosjO56yD5LLqkNVPb8Kvf3piDOWIGwed4m+vtA28OIBzsjBfzRMxjTxooeyM+ZT
H4q8ckx94NpKXhVMjnDk7GbKEyOaFDYqFKLXR6gWc8gLYqjfsuJ7wopXiBJJUKSittbFL6PygNat
YMgHpD6fu1HFHti/1FZh+77JsMXcbqK4npEWKg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Fhfc/5jLchB8UMNqJHMDzvQZNLcuDshmKQFSwlknCJXigCIZ9WOCmuBoElD82bJoMGVD0EnmP9G5
XkBDb9VWqrt8IF5jg04lBslS2OVSTnH6q8tDgOAijS52+ZjijXxoItTPBRBjB9qk8Xca2fChv2Bv
ypqPnhoJ+PLHwa5XLMo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
obJ+3C9XZ2G6OwGodfED+POvGEqwOkqxdjwcbMG8hTAX4K2FOL+TxvpYP0ISeOii/wxVYFJVJwq2
UxPYRWvoLsZAHEVDxM0+B+VgM7DBDh6X9g+/H2HingxxUgWiIOu6CZZfNCGlAqLIbnX7Md8FomuF
k5+jpt7zOlg8DRfgFDmHP3freuTKnNq/pwl3uPSPMZoXd0Q6vnSS6AE1o5X7YIc3pYAzFvNmnQDy
vVYCeztFXTM0/+Cw/VEj8xaV0/E+a7/oGK+Xgw0Be4ktPDsYv/CnTHViye4b7dbdGwnuL0G5HWbB
crLkuH+Lv+iqs/TMHYWNf1O4N570RXNmQ+QSQw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 58688)
`protect data_block
rrqYTjZHLwzGjoGFI4nf9pOuCHwZ15sJSh1CHGo+GhjkX1IelIwOdunFvd4ZWXVlitvU2YzaRSeG
57JWmquq3ZjCF7r65o+MCeQAcOlPlykKRVqvx4BcSjd6XtkWPBC/mXWHJmbX0JdpGycknZlK3KHO
0Rqtgfz59QpmT5YUL3aKaHsZYcQgzJFbtefVjGM0m8/3F0igM6JzP8sFjY3ozhB9qmHVHWvt/fGt
g6lcJE0k7EmDMriOVrtCpjcRKlTItgcx3tdsqgexdWYB5QXssS7s7lKqjBStEcj2BUBWBRC2aKMl
sSMb+ExBdgzlsfnzA+BySLZkTomwsnLXjm1vKfOwKIG2JGTyEhcbmyXCtFcX9kx9O6z1kqR1m9JP
UMRL0u01cfmF+1Y42Xwa6alH0jp9GKMmEL2mo16gKGhAL5dpr+LsOV6/bH+Le7tsBMSdTdZ4PTYz
CLA39ZAU/7q/DhysmZLv4pbjFrQCJJJ8DIzHNF4xLuFS5b2SPEI0GblT9Vt1wQLnY+LWQd1rHvGR
HNkMtXhV9Q7dufKAVAAHpYyix7QF5uaHWONeWd/aaqa+nV+pXL/K92XYGhpJ4kg3K1evHhYHJp7u
ECkC7kC5Zm1Xb40riDphqHX2LD/P6WBIy/zYt37Pf5UDQtx9GWF8FISg3Gt99ZbWNtCz+V4KTefc
9I8UKF/ecc9+CqSpf6YAmYKwuogG9bLsQ0pmo9Dp5xaICR20czOMkGt6TNB3lZLGvBqxoMPtaynG
o6I3mMECi+zFxnViSktDpAkiOqv/URwVMrENnU61Stp1ySYYwK4+Zf55UBnLe2663HilvWHg2raR
6eIkDHAAj09dW3nYjxFIDnDJxHwkOgeFyIFpms/i61nrELjcJKEF+vFM6rxKLrt0QElDLxPxoi66
1F8uJyfKi0r1+4HeRpTwrbrFo+THYFnwt0qDgDtyrISme6zF7DBEiRgzCMmeOAIJC9MyyJM5ecwH
ehlvom1ssIQAtFYy2p7FzsnMphsMu3WUSeQsodyqTJR0NCEKMLUjU1CJvy3CsH7N6FdUK5bawO2a
KUF4Lw6rP07u+rOOm77WnXFidOLpLdNsJJRev0uJjAWzQHyvGmj6vHdr1lXs+9aMwOFmmp3+2xW1
WuzDTM1P1pTLsCOd9LMva0XexR2z7HAgkA0DQkygxowjukq7URx6JmQoIk/JZ4TiTusF5LpPqcJt
72Rteg4jgRrGLIazAbRgMbZN/yjt4mXmSliPghzWNYp+uxFRcSV4+9xiv7zA5KHUHsdmdub6Oav8
GpMNmNTM2463FEqXADn1Ywldm909jXDCuF4nB0laIDV4skHYRRp2fxGRY48s5d9oWqhPVXwiFTKR
z6MhPKwGHwBp90THpVNipc8R+yJgle7l0SDHmIz/Mi004nKXhV6VU1L0YQPEfI8E4xQq2JAupWaI
y9m8c8njSKEGpuSEHStg6rR+c9qkRYBKbRNsFDRWh693ScW8aAdKsVT8prmdlZ7xEoTTgCj+5L+C
g0RQ3FTeEnCqbVVx0PVgfXT9uPJbNPtAWCpHIXwQ3TZvN6YcvAvb09Ih0Gnm/WYpXjifX6JdTMvC
1IKrZcpnpFyUD3L/Y/Nmx+2t5Y+ZtLN76F9HnysurZ7V7rBFzXG+7xYkNB9stAWc8HvTxfdWEe1W
kj4VwMEn0Kkw9CZUtHXTHD4Fp0WAlKh3se9mlyQAGspdTdIqqLJvGjg/9754gLxLBKMGli+k0hUP
doRwik4N/ZlDvztEgKM32a1b4MKoSYq7QwrxqiXIbRMChDwULMcjOgzy8KquAU2o/FG20f9Dfkq+
AWco7K2o4hQg96lmXKCT2cHzmevDDTmPqiQ7IGFFnZK/H+Zkx6FtumAWicy1hIg0sRv9WU3SkOde
KH6Qu/wEyGemtxVhNQPYv8kJ+YWo19xWm2uQufelTtDXxQMzY0GyycXYPiwpyWEuSnS2fQ9U0Wrw
5rFGXPx3NiC1Lf7nQslgkUwpzLAykyUJunJ8y4vVNf7COK8GFG9boMdiRcrAy0tQd8aM8hdGx3mi
JxXWMuIHJ/oGAB0GPuDyYb7b8GW0vCcW2Exco7a+Jr5sWPo9CvNqZ1AwLImUQE3WHHUxc5nmi7H6
iHfJrCg+wHPxVZP/zjPhXzIU3+8KmDMhKnMTYE2ENsnVZkSc+gq1aAB+N7tCgk8DsgTTXhKF+aHr
H/+SF4OLRIDmwwWmul3vgyFx1Pdp5xcCoRLOh9G5SKRGzXUE4a4hQUT4NPGCWjJjXXdIrGo/C2Aa
8IQ4njBk5xmCaA3hMas8JetkRxxSGJJ5YjsZjUwjg1L3ZvwgHxFa2RPOl11NOsNTjEvZ0tTus3hl
tLTbP8rgcMVI9ws9tVQBL7RcJyTgHOfYa1zCkKqUM16rSR3KDP08Cxp0XhP0rm4UsPOBN24WCWEY
QFLDQ6uBWA7pZSW4Kf4pJQB1phgI3FddUDOh2Z+NbyR+eZ9ExleXbtgUtxIyUxmnoGyvKXb1IOFT
T6Q9GkE5bYzHBRehrgFiVXrCNkzV2Ri/fr16buEmdFalj6sbvnplOIVLYRtr5RpWHYNufCJBz0gz
Yh/282HT9sDBDgALFMEUYQwVaXgwOuIcvbCPc4XiWOmPzhjdFSFW7p4Aq17VdpT9V5pjC4JZ1sdN
Tcr85eEoVD3T/BM8LtoKrOMZRc6a+y1M5hoXleKakHjvGyDmyLevMBi4yiIeY0DimJnrPM/LN4pK
MGV93dK1jP8kZ0Whxz+NdAZW22VBBXeLX7ZU8aQHR+KlH/+yBJwZWx2Ks/FoUEOmLvnnVgl9V3jf
ZjvgcN0k7w9itYbZ/vZ7IOE7Vk1vDCTCQLpdy0Eu6OmyR/JZla0Ulj+lS6U8QcchujolIrXHw7WI
nGh1MbqKPYQiH9HWEY+RhEFk1lYhrf3aJg6XHOC13Fk6cpDV293OJPWpMYmyfeVfo8Bzw1wr7S7i
L8fdk3CVK7CJtuJP1T0QT0jIHcDWu3UzqH2ZGTIOEpAVpfDKT28u9f/NzNCePhUkPMne/M6JfZgF
z41cjwc/VI886r+Z5sUQ1hS7iI/wJqtt9m/wHqLJwTns4YtDPykRjArZBtwoby6sab5Fmrbv2LXc
p7n+bsGK2STFIhhGyNpH6y9n/68D5MzXc3i0/cC12LSCNGX4/Xz5JLHLd8oWfo3rCr0NvqWCveay
aoyQlCb1EwdL7S4sZF+el1iqPQKYTz5gleajqcGFkArX2ucxiRQipbVu7qqUCvzz96ToMQMe9ngf
igRI4Qo3LOq6jJhG0im7hiWlbqPWhXLJsnLSo/c3ZpPlugB6Yg78qMfqj3DaYKuQG5rca4iBAieW
+gVME0xY6rrm7s+SnkTZAfa39L7VsHwKe8MgafEyW3q4HFxnQtGuFXpNjAcMdIsKOxeeNJneiqzf
7za+71/vlsMdCNc04N7KAsB2gN4oWzw8jP6p0NvuSi4r96zV8d3Ri8B1sYCWZ/W/h42npFH+nV/S
UdH/AtovOEwqzqVd3YAjXdTZNikriITJUNbXtE5qhr+MUsKw8KEwH9V2Bwr2bL77fIzvGUThEoh/
PwVcgI8gmlaCF18HmefFbfGegWUZ1S5SPGC4qYNP/g0q3gI5CEyWkJ5hlOLBWBt/Yi94zNb9cvmD
ElclBsUrPwA4d/O9cTcAvEF0x6X+nfgfM0xtk8mej0e/GdpLTF3CNX5wVrZVgat1gg4QP7PaHApw
05zDTYhSFqSlKF5b6O/4L9n4dpVrevSgz2pljwfziJhkQM5GJ0wA0drEtpsh55vQQFPwCE84zP0e
Jzvwhv0ULheVDGgOgjwFy8CexqQLMOIXqKh7Q4Y7L+pP8wmoCah3gvC4rA8WPGjV8Cm+0XYs8X2t
bj1z8Dh91MADLi/2GhBNDkWS9XG2JsiFhFXoYRvd5VnkaX5jBmgB9ZIPSR6Butck24fonh3rZkky
p+Ra5qPcC+mhhC85m7FOYH4ZnrtPyrD5l03rKzm2iAdLOPRsJEdMwWtZ1bKlXCHO+Gg/7M+HQSIx
iXUan8yrra6PbXjKLDakUet/YOKjVIGRF6XvPYwhZHS8XpmzlyJsabwycCWF+ZnwRfVFKVwcsPWy
KN+1SKaPdfqTlU+As4KnYaTIRNjUZwLP/AU0d5NrBOUXqs8vxd7U/vIJES/w9+vfuD8QWvrfGYaR
MmScb7JSS5mcgJ37DUMLeSAOaMY+L/yVJG9X7chWF8asrx+IbgqsRVPK8FMUwSTO687vnv3MNzd9
MF4ICwnDYBxyt6c/8wMavm5x2oXABTowWJdKhH4rurrmnkttFk7woUwtlw8ui1qt9TqdjGQqaPl4
vKcwjMjHgsIIpwJJmKehbydrSypqIv/fG37VQYsP1XB8H4NQW7KMIuEb5S8i7RD2g+JN52jxThZA
mcxyQwml+vuTqykohGYxaTrRCH95+yBaNjqSNK3A2FTLBUKCBAJ3DW3fQb5BKa5npOtYUULVww+Y
WhhDFGR/N/f9XE5HanXna3pgmCfnykZvoO/M3AFdL7sVG73GFiVCHK8pYgzQO3wX2+7PJZBwZVkZ
PZARJ1A3m79feYNauek2kPPdizEJcilSQJ5zvgswQpclbgkU9nzsBIkUMtHJRlAozrkhnyF5xuWB
Ffdu/JiOQroA5UbeXLspUq1lgarazi6cWkIQ2kkvzqfRTYOTP0f249zyQIWg9F1fJmLbEd+ikQ2V
BWYgaDz4z1hIThBc0XBl10mwWRmMPEYGv+DZBwMf4F6rtAG5RDPXPYor/eoHd9lUGs889B+Z3qZP
Youvd19ziYuh90BUT5/AdJtW+f1A6xi2Ce/FY+s+ucvjqecJTsmTgIwlSjLBSJJQuN0FEAoYeR3F
6SKaZEYYI0iHBJkiIwX163X9faDbfoqpyHQip/lSFODlq360by5b6txs1EYP8F4exsEWtwwmV3cB
cSqeqEba8IDjU6cb6pP/jZW+0XlN5dq/SssTVaIXGW05Vx91TGyf9jVYS7Weq3+O8pMZya2iqGk/
/cud3JkNYA/dfqg/S1U+wuXNZ/0orAf9EamNjShzkyY98Et8FdaE6DQ8YIUBP1tdLVRQ/kb1O8io
QS/ECLwoqPLt6yorO+sKCy/0LMckiMRaPVFQDIsJNfmK4QltFAml/CNIYGotcKDLUSbkYu1HjU7j
kIxvLBmucz7+rJUZ6WWnhbGShciawFlS2q912j70WjiQwU8hqP8p8DmU+6/SFkX/X2+nb5ZKV9eL
7hWTbcY3SbFFXeJmzmnwsNMSmgRaFP3t4Cs14cgMU0vonIA3ytx3Kz+SebBd3o+Mt4qCef3oX1Z+
ObZnxH0YT83P4ZJR1oIKqRZ2CN/oHnzZ37+j5kYrPh4HJV0gmY+mlVQIoznUeeOfWrciMKxq/mVY
URSSYj2wLXBohN6xwkFIw5aNC3TurIWccy7xpB+MwaNFmKqvQiIxnk8O3olTbZllgZMQTsNtGNXj
eycw4NFdK4sno7k/zfC3JisfkSeMP9jIcwxXBZ7DjBNDUQlDgp/QJ2UoDUpM0DwDAArs2N1GFvau
9mC8BVYQtfDGUNH18WKmeEuvZMDMRiBJoISyC9w698xL9v+58EpBn+3LRRWjsanGjWQMOPXiLK/F
/H+wbAuvNrZ9Pv66HGJeiApM1rXOBOqN1rD52Ago4OmCBYsdWDP31QvC/w8hSh+khM0LPxsj0ffy
Qp3yZ4kYvID38/giNyb4sUAqYCPUfF4dLCLJDyw/V5C6KJMw1hf7I7Fc5hMap2pS2tw2LV+X3pHK
TDj747hyYzPAmgrbJs0T3N3NMAuFijOv6rIaZ3BizDKMBJ14cMUHLOXB0lMIpKUaAytIM8YNp108
y/y4mwx6+btcKI0+99vTVVW4mNeU3cnjZ8haSoiqkz9pTShnlXV8to2k2hcXCcUX6xmOSTo89qGM
tCIsgYt4iZivqoQEBc6XuCDGzgPRzq5NIwzu851TdbTGBhG03CWJCa+h7UQc5xA3rXNPY/vvwxQo
KgKjLFdyHG8pNbRT2oE7tqQvnuIr9gODqxFjHfu8jNo4TbUtDqz7dhD1XZt+ereRR/AHgqcXwW+Q
sj1nYSXe/zx9WADb0L0KvXnXDbYDObuBQJ4ObhFFuE/CbVVkE75NM31YD0CtFubbkYppu3QnntJO
L46N2uagHAW7mhyPdBpm04/wnwp2iG9rwIJ7e035fA8S9E5iWhqxzgrVVQ5aLXQjc+Ixl8OI52G5
WyWEpDQMZAIXq82eHbsACQ7BhsEjQqh74BObarUIyANcYpwest2lqWZLonPRGZuKH+++b0/DA4JD
4YZGnZwyBVCUC7OMXid+6YAzcIUdpCSHbhkOC8j538yRmA+vM6VNl7uC4HeU6VfkMEJmbVVd5wIB
C6MbCztqXwwdgWCAt3OXdBnFxWHDYOgPdHZCdO2TwuB8SJ+Ej9tXltJI7oL3c8Z7p28dp2h9x0fl
uFKe+9oKp6UB/n9Wf1Nf2iPG4SDXVdPUzowIQBWuHG+ArMw4mqYYWGc7HF8gbqVZ3tVh4T9FV6IO
rV5hWsYsEtUPT9TgEiuKm68VCv4vCDd/6cENfyLTGNeKQa2X1ih9xCzis85+pZmkzJvUYtLr5jde
f1HfZxdLN1YHHITrSCXqRkI23FPpbBDR+Fpl0wimf8TSYWI6YomB4IuKV+2KbcmIuzj+YrTO4RlJ
SVk2w5R4FN0jJBnhAB2CRBSZ8Skb3MNkWyPTOd8S3U9DJJH7uKpZcov8KwC/ac6S7q3loMa2K6ek
nyr+Z41dSP6fYcx27wIRr8A/LsN7rTEfD7E2K1S7Gkj90RYqWxwcrexkkoMUOnUz5KYPOEgJZOJ9
wpzOTQbWJjfrhtZmGSLR/ke8L5WZVFoxSLhQjnfyyYN5vk3dElSJCluLaXe1fuNQglILtRrnLT40
JJ4N+Byj/o+CijXUsCmPxhqDfpE7f8aGqMqNdqhlZxHxLpWnnzHh423ClvhdwLrFwQHTBuhegtpb
x51j12TQfQI464dpjKdppJrugPr/GFfuSgZWjpPwJXQCTQ+Qx9eq2DUXmE4mN04Bu08BqQKkpS0z
C8uEYsaBmfIhWD1b4B20oz9V2SWZv5yabPDC3Smae/rILBQdxThjmr/r5Q77aoQYWFevAuxRGXL/
1wJJHqdpkfORNrqlQppVQGdML8ISh4mPoqarK55GzMUS7ef5E/nDTFgp15Abvtjp4b9Sv24avodn
Gony05Qm1cGz+MyNKDk+jI71bCz21dVZBMISq/36O1OcS57fBxXC2rXAQ3s8EmVFTyNeUzobDY9z
zaxPpmnUCvyW5b1MLpuazojeFcgJnvh2ALGVT6NJ/7cx199xTZ51UwQiifzjpUMwNwh/YirGP+Xn
0YEh3srpI9lh5cMRa3kkoZJfRu+CZwmIRHmr/kftNQJyFum8GjZt0XuOhhRRblofAjW2z4Fv3YL8
VozH2Oc1iVtAAmvUVNbpYlnwkCJXN6B0CSouq9yyp61E0xJk0B24Cehv0J0khjHJzjfrlaWzxccg
avLoo6VyQaOzjUrGuVBhXNaSUPrRl6rBWhOYGP+pBegWAkYUpwxJrkj9Vd3y9aNbLIkRnFaDk/LV
xrUkIqOqhr8Mwl3XrwoqwIQp+Hu0TgbqKR2rGM6Xn8vIk+2Lump/6TXLkjfQqyjs22Z3QTNszrB8
18S9xqTTpNUutg3Kv4PioTWGE0nMCNAwKcabSENdUK0r/BHg9pe+CiXB5a1lDESviPXfhPTFjIIw
mwFsFtVCZqsSnmCWpOhXrk67OKN4Dt/0NGWJF11y9d48Dx2Z7VxhEqQv/9/qphCi6ZsOiv80JljN
oJ2U0JnpQCnECBsYnD42aphIGkqgvqfJpJQcdn7Ml4/VSZxc7cfFLhuuj4SnUFB8y4swS0chRmni
CHn6khWS/vPL7I/5aJmiGPP3Xbsb1MWwb1LwAZU7fYRvBbTRrghxnIMLfRjAotCnohez45CHP3aK
O7m22FupEshcryKo2qqAZ+1h/SbrMDy6EELRl/LswhV1BnPuyh0pEgrSyHbrKP+oRjWT8TvA00tE
5prewBw7F7+gHyzyoL28FPvTKqtfeos43kP7lobjle7pnGcGi/ZauJUhBwKYVrKti07IAPPwxGgf
aIEiDghFMLf24Qsaxxm5x/LhYjQa8PB4k726iah01YX9p2wjJbXhKJ7rNdtdwZogwSy4EG+aHEDm
16mW7NcF7jredydUmgvTqeWcpUB8FosoB6pTyd2RslxA9/kj0Ul5bvjT6RY/zbFAAkjQfLtGoBaM
tHODD6O284V5xX+NQI42Aup0/Fn/87bbnDx6oJ/dii8apxmriBM0FCPtxE/WXZQme9mzJcZd8fBL
IhBZ+Q6oYvnjEXxayFQSwEqkjn9a8NpLrqxM7pxtHQgynDvTYeCS9Ub4QQh70KCadR4dUJSVPktN
z3RskQD3yo/z02F4AOQuphrt2VQcR15J8VKjRKH2Ri6nkxqIlwGXP5P2TfHSU55T90ho/EzyW7nz
0sQBi23AK+Np/cfVjynSm6B0K0PmjYMZL895kmPaaWrGvabBnw0VdrDZbGx7hUI2LXHj18pA6Dho
gTo0cKdgZVa++POReUATBE6RlEgs9IbdnopveFY/DVAi5o211B+p3puIHjSbbF1+8mwE/mrFsOLG
JNZXj7bANW/wq+HM31s2KZl6ZmmBnjUm7i69zGs7d2VSlSQChAM49takGuwMx/QIc80ASR1gqJJH
Dw8QukfVto1Oa7fBrL2ci7oKYXWkpNDDxRa9csdX1Nsz5J4iaCM4mAjMdE3Q4OJl+G0kR1qJQXjs
UY3CarWE5JlSv5ajjdGBcLLQTmjIkHxb9M5m2Wz8cuFmpIY2sBI/v5YZ+tZzkVdpUd00nppLm4/u
031UwQemzHNlBpsy3JFol3NrBYr2ZxV/dcFu4yyVf6PoxPpYiKy3dcVtBYQyp2eiwC8TAuqUMCaG
zB6EaiD8qU9clilQkjrK2D7N5/DhY/FGSf8i/f45BcdIQ6yOUof9IP5VgYeAzaBz4MVTUCVJWPOU
v6wDJRALe7+FCw78JgRCwzlVqOpH5zIh1+5fE3EKlNfLAJAqNHe6b/fjINJbVAe/9qe5f6ZD+YEm
GeFRi7sNzQEGyWYVqX0CurA2EHB/xofxLSE98s6hUE6zC4h8yywnznqO2Ff7T3H31lvCWY+x5RAz
WPyrurUk/sIDy2DleItEisIgxXjW5Leza0JEPJLBZyUgjhOldwAlSU7t7FwqNTPpZbf2JazQ2Nzu
uE9SBwbZd4jvMuqrOePvJaynoKtKOTh+7YLm9vtwZD9+Omhx/5AYadfeofwAqxrJwbi3+HsGk3TI
E50fAtEo+OkyAqHQtdMGUQ9nVN8VRFTUp4v3o1qrK5RQRe3s2HSj8RiNRXzBsCpACqP6PPFSj09j
4oznYkkviYUFtF7G84W0tGBcFPtDY7OZpq2GBIzxfo6PfavAULXxKis1AaCrVAtUhcf0hVIPuNt0
aZxKT3n9hdV3Z3a1rc8nvyendOC5mxXToADBX1suQzewxN4Y5l/SvFL0CU4zjbaTST7by5j6SNW0
3NbuPixXX1CpOu9qxiVfjN7ozgpFLtVTTakKxHjTazwlGUP4zbnk5kphLeOz0NeHkvNv1zFzwCVk
21DDTqZkbq/PXkbcBfxI2Yt0k/0+JTTeZMFIhcj+FKSc1sqcyZ4zOACiO1BPPu03xF4e+h3tAwiY
FPaxW1IlrgDASpbwRWi7Ex3a8FfkFnG8IFdRwYwAoyM27ws6yNmJOLSYXen2VdPnO+gM4dgf5vZ2
Ck19wIna62zbd56tH1RISadvK/sWrtVjC6jyKmRGQIQEFT5tNQN2PyTEu1wJqiT8MpGxnJVL7V/J
cJt+4/5xua6UcqEAucR7UB/JQAy3LQ+9KyrBuuOej98VrkYvOfa6JitToajOJzM2IP7/hZY58lXH
vZ+WNG3f0M9G8NLeqe2Syo6TklmR5DQg7tdFCaUf/HMuTxkIqe2jfAiiR0xlPzZR8LVo+17onljL
XyzPqJVzUzPneuLt71tBwlixZpsZeQpBVe2ba9h73DIidoHrW+5yP51SACBEwDG9e74U4TePYv4j
r3lAfwx08fFEFsG66yyNPPuylfWAlga+OapQF7iJ2Clvj4i1g3NMWTesdYuJPq6n7iplbrwYAv8R
NRkAWYAN2fDFMgYf7tCfAePQ+37rLy8S1PvFIpduiVuFTXfBlqx7KNA2Ui9+JI+1r5X54V49XIBQ
Jm1RwB0OosBdN1cbqNg2moraQsPwqYEwyfkWycHoKnRaltSGFkXvXGuf8depYrHKmtDFHVzzh74p
YYRfF7YX3xMpTs/dzwBciru1fgzOb6+nTzu9JwPeau8qeQLPQyo/S3NbE5Oe1ZNNou5qDHugTfK9
viS6bVswtJ+4gAb0Jj5ImYZTBFAfQhzw/gyyTV+G6BSWDb5D1jsyG1isnFvXS8aaKioiPDenplrY
ieCESFT/8C1Yk0mmJpL91gF7zrTCm2euuuALuNTZVobNwUyVEmJsHwP3iHTp/4GjCb4ug7//vZ+b
xK1UpawKhrlqeA4aW9gTfAYFLJC+BwvORRqo8UVOroN8w++8xoiX4caUO6vNAiwqVhA74QhpzBen
la0hAeR2Y5zntAlPbQvuJi/VwxFY/iJWRK1Enie+Wky8lNrO778G4QEM7ibf/lJox3P7jYDkeFBX
73YhzlxKk7MwJUF7OwdMyzECCfg9yvTJI9WsvOxmEzNBGL2SgITh6fML7iqLo0okOIVw/zwjyY1w
CwnPJoRfeo9UXKXAqs8g8/l2APv6X/COaZivBOglvoIzSiWxm6lwVJ5VV4RBDaYa4Q81fuyN0F7C
9BDgqD+GnX6H4Fdy3DJuku+VvgRqmRzWmrJE5NmAEvu61ZfpWF94PbhYPqC1mzOs60xA/1LdQLcR
ihMs0CEzkMjJ5gx7qOg//4bqi4UOHY4QdcRh6KPdwzycbflY44Sabxgb1aBaIugG9X4u+xZ9OOSt
iVJz6um0M9NCBk9yp7COtnOnfrvfLdOTw10wIDMHSQw7MH6hhDRmBKqnm1mLj1MFkcNpdOYEhhcn
F77iOTtbtw1nq+UAPb+h4v/tn9I4Mjn10PjVEsVEa/cklLcHbBF9umcHwbh0znKqe75HGI5I1nfZ
YoAg3IS3SVFBOGrsNqSkVqMBgKiGzGbWOidZ3y3Dh6vqxWZLPF5gJlUwfao9O6dJqz5PF89OKvZ6
sf1o3th4kk/fKq99Q9k8wDsSKEEUBearp886WHDyu0CeVyHsM5yMTx5F74av8km+Os7Y/UmxuETT
IalCuSI2HX+jIULiXA6J/es6alijbMxlyUhPnI6DlkR1vlKS8azvt5tge2vX0MVewC5FngKcr5sc
E2fQnSm/QgVBJF/XBYlhJzSe0EF8/i+M5zC/zDgRuCE87TJlzTYk3rz56Hk1TrkzuSjM3GPx78GE
YKfnjms6Txyv33+leTOceqZKbpbqSKc1CblfIU6W89iLOrJVIUsvBanCpI9RxLf1AcjIb1BD20yn
hzIVaaQK/Rsd+IcCpkrRbi48JktT/XGUTpxt2NskuGmEmZUM/ykjP0rgydywXxXL+Ke2z9/ks1zR
WnsUvvZ/yQN9lJQp/6qBZCvCn8AjPc5+bnx976gEZEIkNxSeaKV1iEwK5c21bHUHMwPg1Mn3WyPP
VanCZVK4SGdMlFMh+qBoDrBP2Y4tMhlA0hYZJsi8JdB7/zyi3Pw4yzRnk46BO3F1b5jN+efsWdUV
rtlEgylmUO+OTcV52fmGy8rOZnnVaL2BexS5ntVcNXeoS/SutLzzYARQ9ktuftUr3vY0bUdA/X3U
/rB+IFZmPZxAsK1A6Ox1t7aqrVUzONlOFTzamU2lgh6SxW5aQydbLprrAE9lKWM5Bvx5KVCym+O7
18mqXib1DvzUiclOsy3TlD71mu5SZTxMROmYhCNKK+XlpWSuyyplO5YGb29PDhLuJdXJNwvWjciI
1XrsTouwNXr19cO/j/G1rveJPutxUbmTqypx2VdXbzsDnPYR3MuzblcTPRe6CIqT7qZD1HjzjENA
2TRM7pk+4jDy1ebXJmofcvY0jWe6L4+uvn5e99wRokMKCZWxK/wTans4t+ocPPJEvfy3c30cHK/V
IurtTXh0I8GcrB9FkNi5npNHU4V/WY711C7vybyBOQq+ZYpi96Tkp6q1LAcunJK7uYh9uM1itZRA
oD8zf6PucTBJ6lC8wi6f5PyuX6xZaz51Ppd2MbdZJ0f19P/OEOiENKOqwOo7kQOVn22a+UtpRgSd
yv4zfIBahhZfoBL5YloCltNY7qkfAiVCU7sB0W8b0Z8UIOtp6+/ADfnWTxFbgnXSRjSvKerSFkqO
NOcR4QrqMb9iBCFMvhVGK/MgBC9sZ3QbrENghdyoGQ16yY0EnlPQa7FHbOkkj7tE3gyTRxx3uAJq
8xUemurrGOvfo/uMfnSEL2xLHZyPMeWUST4uIdQJahN95J92HwKYo6hxgLxhQmvQLrWBNVEAzGf1
k9WknQx9IoEUUuqd2FMFzyx6UnoplQAyG3DtpFkSGanPCrscp/kAOyLvifMyGz6v0x2FKDVR+fLQ
g1GaBJnT/Zr0J4BzQKOCYVb0poUzyh8/4Zpncw3rw1zBKO5qCTX27Ij6eXZ6r9Ww8lLxB2ozgAAB
LxwK2MXc5IkMJWHyrGO5n9qtatXEEISmI4Yz5C0UIblgCLVoFl8XRgUD1uMp5SRFSmf1PSlK/0df
VVuuaJsvd+Y/XN6r08qoaIZvLpXDLJP1hjkIzrk9tgTcZQPHYMuczoCgIz0Sx1VlwOBXktLWcNuZ
c8uF7KL6/Yt5ZUi1PBIfoQTzQd96gTO/Nz4AVq6q1n7nRsadXd9bIYYDDq0aEd4P2b9cKo6sxIBm
lQsYKNnxMcENNSUZ8bnaAD4jxKKXoM/WTi2cU/HcGNOX5jxPNd0EX0Y2Lp5KfY+HGLXQVhWyIL6R
GfmuUc4Q5bD6XxBudz/PdXiZIt7vXAS0AAj9doLKOaTCucyXWa5zbLgIyNlEC3u2igwoA749yHHN
LmeFFINGXw02myYfGFGpXzF9mlYEjB/5QfjNOMdqp14cgy+WLmm2VyUDiqTN386OI0tHY0KoM8Jd
0KpgiyC0kX3WIT/w+yBUgjmW5pD70mFHOAeIZtSAWNnKYw7CMmzF3TAzTTKGlyYnhVm5PhYQoGwr
EEs7w+r6nWdmP0ddOLfiJ3TC1oCkf4mNtxwpAfrq7X7Gf671fUMojDMyPImLR8lwCFK/BoCXqD49
1kB0d/dKaH7g5iUR39Vwk0vD3HiXufXVzGDoI15xtJ75/QU/Mcd8K1GtErey7GqGV+zIAQhpBRHw
WhXAJDXoVrHsA5eLon/cw7Qx1OO9/5JebzS57JXmRfKGbuYre1Gpec9pQF1BDseCbGKKgAXeBk0r
ePXggW/BRb31Yo9/GTUb+qJb68oLU839QB3iCi9JZUDzQZ25XgxW1whTmMOxG16QEIdavD8AQhAC
gXiyHelim0i4DsjUgUrHmZXrSHjEiwnNj6m6kjrXS66PA52qVDlyD5t0QZ/EX23fCbmYqXxGIMaC
O9DeKuG0tjFMEEZ3tRBXtyz/sDzxITfHMaQcu5YMSKIUMh1TOFdlTghsEKzzfqm+PAN9vUSgxHtL
Al0YyeTQUa6WXNGOaP/9z4QaPlryOAC9KGZHrGdiNrd/pcDgy0s/0C0DxPXH4zdyQkTbl9tdLOv3
PcQWl4ZoDPsJk5auSKWZzw57BOJf9xMZzLYCS2CZxSbps7jW0/8oFAE4/4Ip8bz8ylGn92DY+BMZ
hSDllMo+jdJnUw0IqlIs8p2D4xEPPQNzCr8ksPUZ1tiuL78phJWh4ptl59cQs7DmC/B2AzfmKxbu
LMlxPYm4geQiO4kKk7viHQ3+sQjmKC49AqSbTAidY4J2rGD2DqFpMDQa4lDcdq6+jgs2NjkhYL2k
67TocNfvnEL7VgdlsBgEl3wq5FlFaD+1EbSJtEKceEHMoK8q1J+5nmySskuTQkkkJkylzupjxBYI
NXEr5J3+sql/T1vDZkHL2w3/I83lby/6c/RXy78RGUFot2AOzoG+1h0tNR4fyZjyMzwV+jpaUguW
rVPoupMVcPBLi/f8NE5ghB4jsmaCguU7mx9rrOP9QItcjYSjvps32uNm1g3uWsXa2ajCF0E2z2ti
RpOOvpfyIqCsOjD+v2VFl56c+a6qLLXhD1bV9syfVvD6FUvNtAvxb8+nJU9W83pYmhsvTMA0/Grm
lt7U0Iwgwc9qPsVDzOCtYOMqpW68SLDv5OTMiUCR5bzoADY8ANEhmz0O+MJCzGVMlv02xJ1xVJ78
A4YO6uzRnBG7j98aY6JfKKN8Odk6CFz1C4UvrXWZKINfrNw/HLchPDc+DlKzAdt3tiHuTFtMQJ0x
eNNuiXzAh1BIB55mgGkX6dv+9YgQP9GHILxFt2uHCdDJxmrwkLCBe7u3z4XMWXDwooqEdYBb8+Q/
PcaphOZlW3CKaXVqH9ZQAgGq64MPl0lJUeernrxfh51Pav4fGwpdiCnyZs5qAJAKoTEKK66Zo2oH
PNYyqDgHyoqpfcxIE+rzur0Po92gu0DwUjReSEo6XHQhlYR/+vpSA4NhbbXREpNasbysaaFsErHe
S9F6jshbAJfy4NtoEjZva/0XFAxmSOwp5T0pXfZw/DRs78MZK/qw41tRYBbFn9lvtqZqy6EpcEup
iu2F07yokGoAkvbDDPm/xHKveu0JflZPsHB/CJAbfLc284836O3N1r9rBO55KZeeC7wcOcof+G3x
VuN87C0OSAhHvH/FtVOwFJJY7x1C2b1nKXE0x2Ji3oU2r8v8aBpnoWIXaU5/ufp8xS+Rq8x+C2s/
6YOYSg+HUCLljprYJkXjpAL9I6K3PgxOVab6DL+dpe04F7a1KOwHx4rs/WatKBXihzyMo0qBfpw0
XnVkaQJuA/1NJZBRyy/xxjoOMydLvu++Gt7NAcGGAbfhKg3CsqR3iOF6ggmPW0AuoXlks37PpRUT
f76BJXyBrq11Fs34REKNknz6BZ2APHCa0U0Bea9aZRejtDyD7E+Z1VELWAwzpos13/Zd2PbyLhnk
98wxY38aTsStrcbDZOSaANhMe4+Ky0sGjstZeHG8BSBZAJ19YxW7c0jHlcWt0NADZQTlJgrbgvLG
Q55JC8UnRAEn5azTcHFwZm6m1PniVcHRoSV/mJfkH0qV17R0+HuvUqYutrAO46GQ9QxwVWBckdxb
vaE8rF2EPzX+VsVBDwH0oBMXQzB1dx1BsLEny9tuKFXrDHn8nX2CU/8/lNToYS1JdRXqcswMaB3e
zqNObyFBFpNJ5H9JJKNsdR3P92SBGPJOSZOgYMscsWtZzrS3BURicK8Id34Xd/ptz5uX0bf9ZwCP
HdPJnIAnPGr8piq5PWB3DhmzpfIRJD7kFLItG7VO1HXML/gCCKOESI0au2crGy68Q9B47poEyWRa
JkjUjDSjpH6uNIcYVK27F862b5GI6GMy2z9M5WaVMlMMYzh6QV3s8ZMLAJBuzqDGQaGD9N6R0VJY
8V2ANH3i+eUaPCNAXvDiyfRGQMtQtjnR01rxHnemwCqGBAUOK5JG7qIPLShMhkk/EhiiogTNEGmg
cVIy6EnVbSfJta7YXrvn6EY3VmuXxWcwNuVxU1gztSDDF81PIzJF0iPUTeaig/xOUjpatLqWcVui
29oA/7RlKwzjLuyY1/+bbSl+qmrv7vwXbkAcrpAG8tOVviPTXR/hpOvaDmgitXslC2yC0gJ4qQFu
2VutL+99NdDlZFa/zmdioOkI/PZhegMB7rREDlsUxgCFYsqxlo4Sd5O8l6JqQkj9Y9BSh8yo6Fdy
lEsWvaR46DI4hbptl1BkiraL2VhtKj9OsY0xasdAugUzqj1pVXfdevGSAS7NoD1zXVZnH5h7mEE6
CWVnlZI409KKJWwZ/MCzofS2EG8ELDHfKdCcFtej30QwW97oRPgIu4TNid7+SWgVj4HNEImnGsuk
O2k5/sFq0A2bYnzsyzk4od9ykF8vww9A5vnFowZ7hhgs9Bj17YLZAUdQmpnz/L2wRAlvrw3YlJHP
bxpEepY99mJ3YPO9pcMg6ILmvJeyRskkX99UTMuxhXiddTPV5YWJ0m+PRvhYzWyY/ipUlbC7Hj87
SAieZDZsQZcpY6q+rh2qVw4FfS9c2SltXFSfox2+masLS4O9vYj99SYOwrt2Bb5uaEGfUVgbJtwW
zCYUsrUqGW+eg/haiQ/tHq0L/RnWWVNeM+FZXiV480KMwVYMyQpvgWy6d0fnflYvL8X8ifftlxS8
m/9vgrKXcz56w+JxbylPn52yw6Pe9wqGY57UOpZgN3omUWhhrUNDkpKvoXY4o7zOzeh6cliFwbVk
fWXqh24lfnpm1QdGnqwaUaEbn2BHf6BvkvkmhOS7jvXJ+VIxqafobYzM8U9cJteatYvZ8Z9ufht0
T0kuyDn/WtI5AXtgMhYyhuDZ0MrJrXCT1H38AvDCbSADISMAQcKNIZBqN7yKbWlu4oqC51WGkIzk
gV/jDHl/UBSFVub3VuhYvUbl0MsobIrV00CXAffxyxjK9MnTMZJBH5V0zzPVhZOI2sa31cvcfdsT
683jM2qqcCWVFcOTlyVXOTco/Q4QrVeCBYLN7r3TIO/JgHKq+O0r2VX3GqHbZ/qscSFPq/LgXneb
SJKJ0UkBRQJ7GMggbyiO/G8SHfLbQdj5Sc34yZUYDPKKzYYFZ3nGpFTqIwQTBGuytGz23eCI8P9I
sM63VBDHC6lzdJQ7ZE/5RbS0x2zPAmsP//MuiZqBWs7bz1g+3lFwYqr71Xcb1cv7KCUTaR9+h49W
WAFBBiglqV2ijA+E4790I5FFOl6LAQ3rzv82LkHNI3ONwd23t5qI26JTOS5Imdj1r/HAJRirJIlL
N1jAISQt+X5AJuoq7lnr5yEEIFs0ESOCxZbk0uUulR1HHG70arLlqAQV5t8MT0SBZcFKf85QDoPO
uLqlO9MIDfd8LjUjrs/cRoQoaiTGawfWp/+Jb/DrShwxK+NwbsAIXStVRRNW0JIa9AYFgGBxRZM0
dds8WJ1cDnDJISu1/6as94Xks4xrAkn2xJB7Ks6BYTDYczFN23JwBet4Y90HKKlQ57HoJP2epX1m
Pw8f1Uq1sQufvEfVRYDVH/X0KFP2RC4QcqeefBbC0Y+dj156CEYV2YNCtjnmyizdHVChlb+M9miE
pDvUqapIXdgD1KpUAV2Mv8qMAWB/mz+0j6KLqJ4ZnhpQlT2zW38aJvpwrUArKA83K81arIr9vQwE
ifwBn2jGWUvZd+4RIX/PLoW23u9kT4LIQBqbUcQ3hAD6jeEwVviLLDMcyBxAjRH9E9iGKiH2vGXD
iEY/Gp3oHo0vUEu50y8Euoi/bWPujbPszX4pNpXuAq537+cyhkLEv9avJSpxBZwb5NX4vvqIYZhx
7YeXSJ+Yjmc12BvRST1ZUFjGIUu7sxtxjNtQiZ4WqEWVMJ7sOpUpzQiZq5Dbey2I1F1h0LtblyM6
/5VpOsMi7zQ20WGkjHgoCWl1cKDAQttgLCypx4U0JHehZLH/40Sn7wK+xa2ubzZsctqTm2d7KseH
PGV/Wn9bnS7uWC3Z9lwjNIZNpgnTIAFuuanHjWd0TCyoQM/8EXerC1b6/zaFVffh47uW64GmPE/q
komDmFaM9h4t9f/SoFykDH9JgB80pB+t37fgUxqgiW75z/sZZva0AZo6zY+aJHGJ4yq1VPjA5xlg
a386wYpz4CNni/fYRzAmfnfhBgfITshp8/UST3QTXYpAUhbL8QIOVHkCwUxUKEihP1RKg19k93NW
aQuuQ+DEreo/g7g3TMiLzFE8EHR8/C65PD5Yi6O9kUG6FH7Mspr9TI6TQ3RAUbLuloXRHt9IeyWc
i1jjagsHePtSBmJ5wox4DvgDbA4RCTmSjwGCQeRAYOAHcWXapdtnxiNNyMlr3yOBzIqdBTmwg4Ow
YtjlgVxWJ2g2DwtGAWow+3PmbVaKfwVEA+nrJPyl3mrizzMizlP4mrQGzQ0fA3IPkptDiPathaNo
Yg+6r/y0789y1tLqWDupPhy/As+4p4Lo3jkOBoyfY7c6Td2pbmJXd/R1WL+JZ8TrPYuUgyj9dVxX
eNksW94wtw76MMPNG1oiJJSRSkYSsK2/rlyxwLGv3qVWA86KAKYiaMM4kePmGq/gPHZWV/ZXVO7N
xNT4BReMuZSPJP/OPEndyOBflWRWRuH/PXNITrJflm9wmEhfoVn6ZrsDanKXIpUQ+e3tEN3O1rMV
BwSeZawOZUsevCGLKomZu5l7ejyAQPp/d0jqetYvVU+cSgMoUPxn/x6XZcyMiHgdIlOfwCQ8OqPi
/m+L42K9G5uFjkPJKRc7+5PLRgFs6MG/TH1HWySsggJymMxO2443cRAHEuTslvc7QUVedc4S90Nb
KfFyD18idHfr8O0QhhSP44AUvWLoKg7vfseXAMx7ihLCH+kwBlCJfMWtpo2QNhOsWSlRz19MEXvr
z2GG8GFYPe8TdpZ0AXzrBB1ZRPPwpPXYBJ9i/ZyT7cOrIey/wp7/XO/LJceFvWuZ17X9+HpjdS8m
JJU/6x+IpNApAIy5gIeUAtJ9yWIBZTFWFuV7Vxk3swUiLhqsBkMS6Ji0gUKBdgVcoBhqAZYPEw/I
xZogXWkyBsWs5xC9BqsOmW9axvPTp+Ao/G0YpEFqlQzcGP+/akVVOFNd/Q36ycy9O84SWhKgGnF0
emHanmvTDd/W+5q6yw4iv06ZfwNycktksgQGpN6h1lMy3B9Ihf3uPViNhpXpNb73uevClYirJ6dH
D05AoeYvGyj+zlNWmL93+bAGT7u3GgWjmRD3CRIb752KpajD/sJ3rEi8mFwurX8GlnzKvHvQsnXy
Wk/h7ytIPs7Kjzxyx5h+Wj2VM2XXlUuv1yXYEE9lGp87neLZVYn6VIPHaS4BH8wPKj32gCf4IHsP
Y2x84E69x7PL7iSV1W8ab2rQerEkaapnPLXGDfYRbevnKQ5nKFCcXRXeY06nswYP25CewFTIZWgg
EyB9LpARKkxDXcYB97i7e4OwnLIOZjfSbs0vN3RGicCfAo+Z/+uv0FGTPOMpZpdZ/woqqhBt+9NF
LpeviQcxuNR84KWvGs/pBjz7/IoAscFIAMyyVVwt3FLUgvmKZnvXJUChoEd0vsP2F+NzS5+UeFHq
jBfHv26xN7mNZvv5ksVmGcGtkIeAEYf63XBIw3oKwahQ8B4JIsl5dC0BuHVIGP3ffHbrhlCx6M7q
5waHiqT6uDthPcno5ZR/HSduoOheM1u+GbPFWZeqzFwSrUKSdiS7IfdcZB63Cj+Hy39jZXV59QSj
hEbCoZMeZENc3DYe5h+iWPRgoHHVOj/vn1FM1Nw+fRNM42YlNHpE0nl7guSIAka0NHuSuou3qyVb
3xgGuHB8hfnpvxjZC7set7lipe1kGBtqlIvS+dI401L+vVRuj4wrXR8xyJRBwGekluSy3oaLezSe
3/5nnQt8BNj6LFilT/u3eBofTc83eD5+ZUXwpq56YX8D2xb7uzsVBABjeSor3FQYMvZ9I53mXvOK
46izKY7aS4k4BvBghXbknnKnNeWVQeTiJ/K4rCWrf24vhI3jxbO+u/gdE99tcTDalpi1ZWkCLyj5
ySS97sJiS14OfFhA0be3NnfslRiU6+BLTn+sZTIq8zjYfS1mH/sj44alnBO8FsuS/3ZRmNhBpTGW
y4Y7Y0EbnrmAwbMhxH5PgdcKq5j2DirCeORDz32NZ1ZdNvb9FbbY1c7rF212nHwcJYPkx3IA6E/S
Z30nHw7KKmTqm22g4IKAvNzd5z7WOVS1o0B0oAioAZrsY7WBgO3tQqpvPVsgCexTn9nRAhKrytXE
IetQgco+KqwJYV0lXPcNHH0iZWAgBi/U2pVo2zuLfntfntJV6oluUZiuLTFIqQlGw+6FDLPWjKQh
Q3NTyH0ax/l7hDpt2xG+zpPr5k9whKJP5/CvVSDyRIyT/mtPS6Evlv/jegEpQFDbQOAl4ULMwzm5
9laVo5aDcDvUiL/cy6aUKGaMj113nDZ1xwWZrLMfjJ1cBRzDHpem+qNAGXZ8Dp+eIod1VqyyKB0Z
wz689OuMpdjwLuoWEcxFFqZpEJDzag1ZG24HHS4Qtrx6DzZB1rfsIiJkFjFswCxzI6uQCUq0NHwa
qBEKjj/QbQaB7vBnIcVtiitz9efXyWwGVY/gbvhLyfKyneFBaNTXy8w4C5WDdYDS35QGsZ9MQIVs
dlCR3jbz9/NhGwJNuAEbCX6PTb646E6n1VucU7vXdr8lBSFmvYuq1R2EwEJG9u04N6E5bELRJrGD
pkp4sIVb5iek6dRMwfWB6Pjb3fHqropyk0a0RH6oG7yGDTYUyLndYfmNKfALEQCNNGGfn9flejTT
i7iI5LZuawofBOXazjAdvIyJDKezqOZ96gGdI/Grk+Fe5SqbFOG2Nqk++lcYUutMPciZpC2T+WtB
g0IC6wSvQKDwB/Doo8MMHs7OwBTC/tQSZmyVW86PqghKPjAtd4kmjOKAkD7Gkdwiq6tS8/J0OTNA
C2ONH/cKApPK0I4Maxdg8IUEkB/JLnVVZlCDejA0EXVSWhOEPM2i9hyZegSpfPQiTJlpXyreFokC
kd5KpXSec/Ot0pw1zY/k89tEKy3zxf2NonFmn/GSZfYiPnileJHLbjK04kgNlhcvMqynPWkDe9a/
gI+XXYOlkJewHKaXVUBAJGENFu//90/i/ZfZ6xLgh+IIMwq6OtLfvqc7bhqjDjwSA4Jw0rU+F3aV
wyYd04T/3GYk6ykaFMvygE2AgldwL2bfjrLKJpH3ul1idS9vEGO6Jc4OF6JRcDMVrUVfyF/aFztu
auziAZaNQvgNruGIhP4LHkPPR/wU9/Miqerk/91lwLTkXYeqFD60G+lzivSoTTVrBitA6ou/1cQU
fYfYEA3Z+Ge46ghRvoWM26tmc/dBSnsfjo7EDr/jBboqZYS1Ue7NPU4jkIpQ4dhuUvmcVj/TQ4Wz
5eGqcQhQMwF26/DLuww6xoZkt4XXfQD1JgfJ1Bsc8ncABHz8DuIAMzOfxyUcgCExJPpbHEsKPguA
pIssmKzIY+Dcu7T8wc0Q7UkDP9ngrmBYhHjJ2tw6veWjDYY7UWKc/ku2viBqUwnkQcgROGy5dmMe
AbYQrKnldz4I/Qyf6MF5/DKG7ZYa8FER+IqW2ejgoBON/IHpA41u9HFzL7Jtz3O84hwrsxtKERcJ
610h4D85XYdpPzPN3awHtpR4NmyP24YyOaaFgyxQ/b0Hp+Mk1Hf8nYOYslxXGW3g23NQ77ZepQbs
dGBZxAQ1gUbpCmZoXmr35PKhLs0RSNgyhtDTxHyZp0zSZBWXNmh/kmdMXUIstZbICAPckjehhmdH
bZNAsaTfkub7xyDwMhFvukJLqGiLjAk51hLEQ/f9dd4TOYjQ5cyYI2oICvfEu2jFdyXfJQ7QhwEP
kgH+9Lqv9opI4gQkTXkMZiSAR2qGEVDI7BLqyrJjDWZBaMj9cFkp3LaVNrbmx7a6TZfR0EXS/0/L
MbiNPscB+lVXx9CFQCyCx/oRQB5LhXRur7e+WFuCput5JxhnjizW4RKlNrU4uWqDcxuPuLa1DHEO
nSNVjWY2lmpzYPmXYLR2l+IJ9z5gpioXfwNa6rb6TqPhBuk37JLS4w9vgzXi1w2tv7iDZHjhYV2/
THyjjfS/GBjPGUwE8/kCG2NYewDrwif0mi3yISiWympmL5ITOVSrxZgH6eJFxfX5OS8x8dQf4vyh
qc3UE44bEE3wUKBFw5TVTw4EtXrmyn7pKtVpbaFZFoyfgxFMnQur4Zj8NkwbrbFtZBxW8/EKnKtg
h7psCmlkGLT5HUWHtD5VAUND6VHQgLB211c6OEIhsfmAVkyDlOkT7vSXSRl4GwPIXx/e3h1HGG+h
eu9/CSkTZugyrE5Osq3Fb+Eo9CsBFvBLx9J7hTNJtNtp6mDaTPpx3JlIdiEA9pgecvyWm3gN3vim
NjPgqmqWG7tBQ/4L7ZpmjyLlEZQW42g2j8Q017QjSnpZJ8bPzFGgKugUxQHbU59HI1GGqZhknXpn
D4sN9l77OQoXEeSAomQbePaXT53/oN0TP8oa7QdA40FEvpBEiNtrr8CtsRlHaikGaH3G2Q4VC5Qa
ROIAe2Z2e2SHiEM+57nMB2JKbiHAsHYhcy1RSzpmF8XWwMi70Gz4k2DaEVtPkoigdJlFxNa3mgm9
DYTH7M42rdmtDdbjtDCfvzqBaLhqq9Fu9vBYivurV/ltGR+w5f8SoqWg9zyQPJ9agl6ifh4Jgfev
6XM2pJaHp/2BgRYx/cWS0LRFB62qsr2fiUXNN0Q79LDfIAx5Md+iftqBSywYv9VkcGt8tklhyMZx
D8z1J4IEQHmUBi9dKkF+pv1qELCDECFkXetCcyXtK4rfaFKJiCyfYMJ4jH7Y6/vtW9HlfaepTltt
cdivV3ivZFkbbs7D+87F/4lOXN7AzIc/70afgQuRTInRaxb8rhQy00jIA54BEQrKWRGyhqkM/4lB
pTwWehttY6hKnUC9XGo1V5CRpDvB/Lr17C8dM1AUDh7ryeo8E7gXVBhy2AxpbVnq7ZDK/lvKCxZI
LxFUxTCei6BDeKGA/3yV2jnGRiR5SSdrYjmOn3vMwOmU9FnxSEaxAf2QvA9CO1ff9dOcD7jO7J3x
OJc0qS/TppFz/F3SzNYrm0+YayrZIpmtkBFnTIO/Iv7u19VmBk2DVoOfqZk6GwCjJdiOOHTiYV8q
C/X6/mLn1g9qsZWpTx2gV5U24GCOoCo207aAogrIOEX51/hmZ8LDYLK9l84ZnBsvwWjNqpCJECjb
ZiwsiDicohgQwAn8ndJyjXHlECzM3qIhWGMcdpgBWoLf/uGraDlRQ+mwzbfIvrDoH0d/PaH58Jnl
4jspRjgwv9Z9bGrp3W0sdZtG8ga56k+vMkaAv1fhv8p4acapNkvLC8bvoALxFDGS44mabH+BhNeb
x0ngxaUGXjdRLmeaiAAbdyhQMwHjIzLB/mhfiDpJ4mj1lWyWhS87OaGjKQvFnpafF+4+qkuEV7ux
tCS0yt6MR/XRZL5nDaGezS3Y1h7AK54eXiflY1InTVXz+UygjNiAQi/l3lys6jt0vnZzwAnG8OLc
NMQqzptaYV2ee1AhAJLBTcLO4d8pcN/ptw+Q7Y5StnoJqoOb2CBIv3lTlRMGcg3h2cjht95DSdpC
RmzJxkhWmwmwlmJ7UqxOCZ3Z/Z0vM9SAFE6gPCNuvQfiH7mcrPYkVk9NQApEqstJbTSZCzz0O9Gb
Rcw5MQKzatASzXL9AvadmkfyVGdHgepLXqZyh6lt9kJlTS/zP3AUIjGbPGUDrB9nvtTtIfsea0eT
Zt7aBxcLdpIYH/4f6VYAVImnqaKkU4lv7KN92xb1S12mHmGCnKx0bNptXRGaMhXx+Z+x9dH3VKvc
zWiwKDnzHGfGdWX12H+CO0W3sF4ZeNKfkBSzO84zgg2wVvMHQ7uR8jAWDpr8WlL4KVeoZAAcITUX
0Sm7rkhKqVihvhsuh5M2FWvGLUQHCLMVsSCoJvoyMHs6MT0pvWguSDuTGHrow/5XAjGTRJUqhQQu
M7a1rTCLAt3QI4gbZ6jdwC+e1jDCXL9uZSAxmI5Y9PHo70R6yA9Q2VihtnF/U84I6ODBGD3ACO76
XFeXE4pmfEeB51LSowURDaUa0/btOc+PcF6FlHHtBFqjTi/dyycSO1dlmSR1USqk84hGfjwZYnJS
vYwc4CwzSukB30cm+jbOe3nlxksuYZnqsEzTZ4imHZ4FK8A5s2r6FiRcKtKGsvIKQMdpcWJRpD1J
lYMuuXXMbN42PB+7yI6jpEMgs5+R62ueL4pWRIeNmw6XaB6VPXLoGc9lR/TkonqlvDoQT3IXl3nR
LQ8ZEOr3TMtyLaBafyLYOpK5Oe4WAKb7Dic7LMOeEjMs7fq4TqYhok394F1vkGIKQ4Eh6wmvxOBP
4p16HeYj3kItnyS21KbshWYA2XKxhKTjygTYKX1jVB/Ol80YZlIDyVxaUp1TxXVCsuu2bir2nNvj
JTx5iZG2yrJLnp3JIh2ATh6PpxngES/l3TXDw0v/a4YdK4y2IOimA7FP6PyS3n1wSdSSy8odKJUU
zCeoEWiBubj60TmdAoyOC8VDAUpXAXxeIs8kVskVhLI4yKFs0WtJnd3D3nzuFdBaT9wtr01ILJuh
8wGHWV4s2MkHW688PrsK63bP7dir7KIZTkcieFjJ0VxRzcWtyXVIK/XhFL7fEEPi/JHCQ2xw4CDj
+ox8BgXbHWmaJweArFfCQ0pWPlKH9QFGJBdyEssmUvmdIbvPRNTMQkQtjBi5wECqJ+1K7ryF8TCz
oXxZatveHwfJU71MhF6YQRSwLUWgnWlpV7oyWlds3VViiQ5xaGT78NHxMyhmAw78GJwgRHnMjAVA
yHDQgJAlBl61qIDTDGniQDGKcSWztDedvhGhG8u3i1lwQnLfj85Oci9MZxXnWkI8qFQujKCdY681
wZr8sHeiDx0p0vMIL1jcoNXRyVbdnN0VWq6yU1S/1E/uhZ0LS5I3wkvjOArqBIqHiopNFT25Y83v
DBIT9kRyE3Zds12CGMLdjDMJ0U8W0CdgmKFkgKstox8msNZtOa83iNSU/mE6SQ9Hv1gZYVbL1iaU
wvK66F+InPBRp9EBj+cFITjnCZkJL18SpqzycZDVJarfndjLQ/AydCnc5LhhunfolKfEjmCSKQHC
MoyrXEU7ZUsmUfIG++0Aa0ev8NTPGkpKSGUSAbYBUbPJgCg2Ou72YjB84ucnQpS8f+32OiVBFSbb
HIn3p7x6rcXAxfz7akIWm1fCgaG0YHaK2IZmNsnP7wWV7WH7BMDpH6GecLI2AHsAdVmk2wqpVlRO
VgO0CINUrAcPVKA+dK1gxGvVw6DBrsTZxQ0V0VaBvBmSlSJ2PncpopD2qFtS/Y6rpRKA+LYzbXVG
SJFbsivETzW5DUd/vCI7Z0AdMVIxqDruwdpcOWYWcZdB4fMG2GLU1b0rhXHs1MqVZVMJwekWR4iw
tYWs+6O48LmZWd4dJDdByY3UG+/C/w9tJrie43ZoH/M4LeSgkXD9DDsVVLJSMklZplh8Xk2xdPcw
S6/sZyTn+Daq2roqX8Wk5ICD5EwBsZ3fr4r0LPd7M0i8DZT8G10JxnmkqdBCBjXD+9zzpnErzyIx
z6p0W5CowuOop4E0ozMjzF04OMzVSLkuj8UYt3nomboA0p/ErR1o33FQCfcV3RYyrHoAT0zCfD8j
Szch2Kqo+l/iiy+ZBDvBHl25/6soCczfzH9tAsVIOn75MTXEN65MDVukrqPOEidonPu9xFLZDXxA
S6pThljK7ON75qP1FVcgTnOFAk+InCZFLCHJ7Q0rEOdy3dXy44Dx1ASSJDtyZy07DtrlWjU0vO6H
bKgmXyWK5kMGvBDsnCcXnX/SBr6iaJz4QEjJ2Y1R22im5GIvSfXB+imw2WsWHkik25rSuPlkVo+y
FMg/K0/P0TUZyITYBCoME2/loaswMxauXM5rV7gdu2nQdxBC4lRxzZfIu7ew+HLcWtpOy/uH0K4x
Y/d510esz8LDUZLbOKyn3DtDkyg/5zpbcDegiZnyBL1cX4lyifqmNEVkad09G0Zq0X4PTJAVjOMm
nYB8GtMeGglGyRAQYJcBkkO0ytozArQp0+rGEZpShevX0UqMHFypQGY6Xqkw8FiPCzBUNYm4frC8
+5tpP73/lrhdiULPSnm5Tkhqp94mx6/g2G1B8XdvHwAGsJrFdvDzmkQ98vIC73QR5WazU6pYsAtK
mCLd1+Bdz0oeV22Wu1FJBBV7vCaQQXZxaQrSa8oU8oMjr8Z7/Js3a4KMtuOYm6vkC8wOipeEFDw7
OvMBUsyIfDamE8HINs0fxqxcLXTKlz8cFyW6pG5lsfQ2U7SGX8Mmv5WNV82ScA5EJFO+WD9Ly9/0
o0RXYxNQVVv7Zo/CVxVJk7sTeYW4wEBvUfAgf9vba5R4ohUgA6xwRQKOV6wZAU4eYWltf5hewfB4
4z/AQapXyCp8RJDIFAssde45OgcVa/LCeNIGKg46QrFAzBeGZUk/ItZ+8GcGxEhwgHqMTlybfVju
IfslAwxuz4qLbAcNIBQDoH070917D9TWtlV9B0O4pL7bJELlaDHxN9c5Az417+7D2Qk88HJNbmNC
0AGAfy6bJfR3R4Gp/kvV3/g22e5IJcvAMOiiZmTbOBr2taEpy0byMPk226qC2BvH0QVbJomV3Nu2
Ngs1karZxLIl8gASwY3Y5yqhzm1C4p8BxyCsi5cX0bfh0KWJ5ya7B0bBMHPPYf10Y1bwA+OVTiaM
9xdGM/RH0b2MHQwMFkv7xVMoIaXvJCNSG5v3SIZgiiuKf3sEBKQvo3pT5UUNCra24yNUjBYLdZsJ
GopSEL3P98Fj3nFYoSBDc5AJWhtDNvH7J/Riz37/gFma2SCG9dXdZdT1p6S/zCLmZzJTD4Cq4J67
FIrtU/CkUY9N7edOPjuxGwlLpyldx2TmH+kEa6z1wc2dfaaT8izTROmNF+qG9AICsh8pmfXWgSID
OUW5DmryqxEZH80ItLMEKVeA5bLEJSXvDkD3B68KTN5BF3un4bf9SEhivJnMKu40yO/4VYFyqTPT
w4zUjiIREMnMr4ldDw4HwXzq7bU8AaHJqbpoHvj5UAyf6eReKWXOl2iPbmEzhjZcvDNaQFcguIP2
iIu8XLUMA2ZwBFNxuqkMHtjY/gxCwj+2BKXDKf1qMe2CuUWcnTR9viW5Ei2ACxkU1fLi+cFMV8/b
4uwf/f4mFMztBFvaUogoW2iomzCbW9xVwYQqsTbMgZ62Js7yJDYwPEb3BARXnUBX94jiNiJYt1+P
ld8cbd4BcadF7L3lepbDSG3Nf+bDafUgyVIajkaDeHDnO6leeIzTAOu6l8u49FbhUtk3njBzmBC4
3c6Q0zN/tFJu0nIl9+F8mjnlpNUbz9o6i0nsZr3yGg0DFDhmkDd6jOMhroAG4KtA7fxiy98Tiu/Q
kSobZT1gZvvfB2s5D5t2GpYlPLJ2gUIcmrU7MsCK+NIcVrU3jBVDxejZ17oXp9fJaFBn4Wg9kfr0
7HY7sYM8Dci7+hhfkLdxFpv4VMYYaixXd5i+hcWN1MAS7VlgCULtdFuR8eBFsqb0ZjKtrcaM3Xzz
rpGOkqL8+hi0Wskru2x17JeoAgGb21ceOelsxeaM7+sQ1qbGfQAmiYNGO5X9lzRJeNBSBNzTnPmW
Y7ypBQKn+B5n3N8sxYZ25PC/VFDBz84TnaIsTKp2n5yLmoK4VCu4YX6ZYjJuMZcM20sqbNsoTfMu
MdiSYYciwIssWXbdxtpz3mLMzfvYcGZYqijjYlN0SbS6UDRhxmHTE9ejMkLAQyNzmjGfFASEMFwF
93ri5ejq5JZRPcqOJ9CRHlnzk+5gfadu22PTwWzWLYXwvuIdeSqvWhkTlLbNbuc4qwdUW7GzqfvQ
eOL8UtwcNTs8JpPYBoNt6ruuMARYorlSfrAOBLI6l/f2YVWZbdzFxHcZoROIpSASZ55YrJANgwDd
T5BMtKwvmGExWZ/LHSB2yiIt5XTCqLjV+gDMATmvr72kvzU7Qboa+dyzcWEcqvhNHSzNKRmd1QQA
sxvuy33MOHLpRd2hab8urh9xeTiVzGiSJPoOiM62kQ2zsXfAKaSWcgErRAFAaq6KjYrGAb3kmqXY
nbfd2ISWrD3dtufLtgQ1yI4l+iUCGzfzittF46UyEo2w85fGg1XdivCRYPAwYizRI9J4+qHRDA6a
6pqThsDDfgyEpaV7zGlUuAK+0Qgi/NX+AKajVxIrNFAB2fGhDXDXQZfoj8Lq4TlFRncsq3Vr70Wu
n0B+J/f1CePtV5pdYa11DUB58SL8Jg0eYRTiDUEiJVm+t4H+rtNR93w3M8n9GLA8VhHH97kwwI+x
fjkvTmmNOyb0oVxTCtzLDB0mAVsyioICAgSi8itEXS+dTm3htJ5s05hLcRG6Ie43mB4dkbSwgq8l
1cD1yvscVohTP9WULMBJkVnWK2OEizFKZeQKtRLbiXa12iEDQK8i1m046qZA2DhTUFwv20FCVpqi
rpl3+3zXOs71mcT4Ms2420Bugj82KTfeNDvjPtyPreJ/1IWcYIfZff60ZXfj3uAnJnK/SJey36gx
x1YmPW1oUsAs9x6FWLqN6jWTlE3jTEmKjwm0AOLkuCWJe7xsLLPtZXTc9izseFc36zBpc4N5arv5
IvpByid1WJ5qSF93bJb43WYX3A3NQf2dkHmax//XAFSFw8m3RUkS/oVOcFFud+SWQs77dz6k/lOb
jdMc6qxXuIPktPq/vU3oKWRWvjXfkjiqUvxu5a9D0u5CiuJXiKzOUmkf9krsebDnzTFunldXKY4e
pvbiLgcLWdcO2DP2AbK4iRYgSU7VJD2kOdh8PC5br89g+bJh1I8F2+4bW6Nq4ImdORava8uhYQCI
yiw7/GKX8Hi/eGESFicx1dvdG35EBGvjE0Tcj2SuTsTnJk1FKrUoT+SLT2EmzJStLUno/WzWKJoA
TXbpChqIXAOGvn5M4VLBStjrtAaIS+ckYEGuipCtwdSPmUZVs9nURc4g/Zsp/HxRgvd1tINy9zh7
DhMDiq/Bx7BAI06xlpGZdsetH95HbMTo0qRnfliSvFVRC/r3Qlys7xpUjpXT9gIUKVVdgBW00K83
LEvdD4oVz2OFu7LgAhshHFwHh6SvOBhxZoPqjp8y3iyxGNhTZyIlJCD+UnnfF3hhpeuqJuC1nERg
sRxxh5qB/MI6dqesgbG3p+hHwzthb8OmDLcLUv3SnviN2KF+yBQRFocKjZjoRrm8NWCg3nq5TyHe
UQjX0XZLmV6xON+makxRGGu4nEKacvWwEutZTuK+ZGSe6RRP8YRXPy1ZvIwCsPva4UwSd4xatlp0
uO0pmK9558ZlvEnGTDcwKtHKsSee8YCnnxRrJe5ab3R9DhCGMXOc0Z9CWy50X6dSUZygeIwSsA8X
CgJS9/Oag+EaYc/aRo7JVqzWQY3oZ8D9G38SZSBCcsNC4qQToO6cXvd0Gxti5uYF7w3IroAzegqO
vCPw6bXFlLeFXF19zpC5Lf/wIbWOTO6lgvDmdjWdoQEmUjzyjL5r9H0tYEbHxbuKAJ6er2g2LHUs
qULqUhWuRdg6tsyqYnh3DJWZQYP4qSRe6Ya+Bmg3mtSiodvsIKvWDQI223AQO/dK0j3i6Gpno5Ie
4UdlFTk46n656jmH8OLD87q82AmvxOKrLgSgDV0W7IlL/UZemTS3uwZoiyZV1U72QJyPQOfwf3Fw
L2UG1o6FZq4SVUqoLU2yUFATrBiBbCrXOLR2dUQjt3YlQQPwWRPVLgFcM2f6S1UdetXByQB2a4JF
INS101xGwMIhx2+48Q87LkmePevHtjupL3maURgFvCpSX0jkLN1ojtL96l5770HBAyc1Pl2wTOAg
FJt44+/MhOhmG2lOqSu1n+1Q9vvdv0CB/8BlqXCFJd4HZnc1EURjgRDf9r/5tPc5H9K9YMbbHpLz
f9q8KGpXzkLuy7VuIWyuCo6XKqUWZNFmiwut4TxSwFyKgGmRSr2DCNI5mRMNRRuejTPWTYrSO1fv
GZlQcQFEhnzxDib78ec3QDzDBN5z7BBhtpuhyaD40PNlAuaaMVbG0gyEOd0c6+9seU3empyOBsOx
ueFNaBw4/bvVojqtAkBjcpqEoqv09chLho4j6eN+eb1G566QYYT0p8/AITpuyOd/QmcC0Xsx33Ig
RIYN6w6ytTR6yU8HZcXVLG+lv4X7DOWhuORRa/p2qYpra0/T8C+lUvtB8jS34sBCgxUwjY3E7D3h
rkWsJ/RxeCB9z8DwvlmEto/+t6dSYt8N4m4vxW3E5yFZxjLvC8o+Fp2N6KUl1n9CdVrnJSxa7zZR
ni3sVe+vE9EB40Vvy+l6gvfrwbMnZ1iwPk6yZAJxfvsBA3T/+ehyx7drFDpkmn7lkqa60cIjBdrd
vQroithfIAznrAnBfmZp+plYQeymSNScOotwhDjL8tvaBcWSZ557BcFNpaYbAF9wQW3BMfSRhnQa
1dqP7mmnDb0iAk+1fZjMLZUh0Nm0iXc0At809+iz3Jrxf8uPo21ihWWVSXMVIReKCBmqw0Rm/mj4
OgTegB0pyRYNm0fYHJ+f2f85vXiRBKd/wvY3kItMI0XtcJHyQ6y22oLETs6F1zwitgegz5lAH0ug
H0sBewoqQ+erj25IepLPOxI2RbXNqFmWvSc49GRSwGQNoiGpWvyUZTbTwyr82mvAn4/B7GEj+vK6
3Gu/CUhvat9xCXzCCpGEKDHr8kciIHfOlKxaKFOuHAXPl6SGNZqjbtnpnWf2MPAN42EBbxDjm3Hu
eevBpNhldpME7s1IalVnAPi+jRL9vASiFn6KmprTDeFTVtGzNEaeM3LVwdsv5yclefsXAmvhZ+HC
iT13rB1pnZa8yh247jys8C3flAGIbbJTjshpblv0ZnEyRtSni492zQejY2t4zf+6yAqEwnRT6G1y
Nq2qcO+D24yKl01dBOPXrtRCeEVPGuoSjolBaKocO4Ss0gOHZOXDnzjhyrXQcjtQBT4UKdiuNDPq
omC/rHBk7Qad/Qrx/P/sI9A6sZxRIhWFolGkYULKWroFSyy9IT4E1woQMQKneDrh7qYVIv13Mo3B
17KQWo31Rb8HT6gEHkkJCJeGY6seZgMitv0vjbDHywhQwjCKBSwRrFVttS3uQ1y53KA2JMBZWfSX
iTLhebh9HhEHU78OGyhr/AZtRY0Gu7t6ZpwcAni8LJ1BM3MvdqqU5wvBhx8fzB/XKASXy2dgfSDN
4ZTSZQugUYIBPtoqkKTHCesqaNh3Jclm/Ll+tcgdGR/cOgUeTIBqnZfv/zUwaRXc/8FhbRU0Mzvw
HzoS/9Cx6N/AEBtFRojwSPKAXo2UvLo3o3Tg7sZiUTWwg65OkJfVF5GsbxwFLOO9rkAvxqKfaaWT
/5aPguTPvoijLYaCN9VTL4+bZAqkMHxRUTUM72eZwUSY07Z2e1q+gBp7WZO1IYoMq5HqtkkzYm02
Gw7tCuWwq7zOccpI+yvJCnABnu6h6XlAOKyfeB6ftMn79W5uPfzyHKOsM6vlHiomV9luvfY1I9m/
0i9xjAWPu+T6JVHW9oIaHtfQQ9g7Y6OHMcrFEkqpct54wNuybc4coV7poP6SWtGYK6TYBcmBgfwd
7rOPUKN7pe0u3G2noL6NT5a/9qY6wsXGkB44AzWAazdbjuerkSqCLbaZW05CMtYFehmbcT019zNI
K/roWin4L+OOXwk4Fwt+lq1W47sGU6BwgHrFNlw4RHYQ7ljHoW2ZGLFTrbXxJIPvIShaLgBDbAi4
FsC52RV22mY4oypMb0xPGA6gwD4m58vVC/FCxK2Jz4jviwxZmwnKC3h7je6jAMSB10CsI3ILb7S3
sf2qIOgd3idYH1qx1V1km1smLZ3CS9dO0ruHYz32EloDafq5YJjqCOPWLcHzOseo3BINIcKF5D0x
0VLiCFAfcS/Lujb+AK0NM+QHAb6aX1q6fq6SVLor+09V3TPmSCcHzvN74/tdo+IzKjAJaTa54TZG
UAGawA3EyskToIHMPXnbghCyjHScGufj/O4OE8kxYd8NroNPL/sbc7K7DaoxN+Ag+SZnarQImxxf
yubngQBg/rgPUWankA3YxQ+X0nYZXJ2Vk57h+p4Pzn3LSOEdJCaVaxHTM8ZVFLVMW+pN9bPIHDLK
z+oO9cPj0woWLyS6G3rMJRP1ymYB6umzKPwe0ofavh1eCOr74Qf0aiuKpQlKt4pxGyJqeAkDx5Hs
yxa2keyNf4mSHq9gtDLw1+pTriMi/XCZCtT0GIsWKOfpNzookmnPU2IWFkWZEXgw6S5AYESt1q0h
tS0JOiIH0cojeYvrYAa6sz9rKR69Ms3OEkHTuw0GbRYEyOCKs3UUwvC4OuSJ7FD5PLkaqfEfM/AQ
zA2ywEgD6zM159/NvIBqFQv0aCKSkM5B3boYucjjlcjB/6Jhl4/Dmgz+D76ZFwg+Vu+5Lai4rCpg
44PiIh2x1qeEjRs+aglAiZKUHQbuWd/AwP3G3Jx/7Ru0C11s//GOfGV9x7xVC2JDoCYMTEJ/T/yC
p9fJDaX91T4DUuJhsWggEEbKFqrmba4sJA3hAsBKTKMhADmMlkkDPeQCUNDQH2+yY3GRJ5JVASYk
+TpNVo2rQq/9dO85AIG3YWHV1kTiJA6nnwTd+FB54dktl5HeJ2fNtqrN8JXS/Q7QakXOqlxjqMvg
AKvYLcKTmnDyFrWFaYW9PyXkhL+iBwIpXiqSbjbJ3K8S3coMckcE2+F2Tnrjh7nSsJ2bNOyELO27
a04eaMq9ffHQ0TmsV7+ZrxvWBL1Lm9B/z0G9mzm4hYp+nB2Grh6uRrN6v+Mp+bZUEpUei5s9fKQr
05AkCD1NhIhlvi/uOW075fn9CMyKToh5A2o5KoiOVUs+QO8HryiUtePdgHGWJkKCyN+0Arg3MTvo
fso0SGFRYE/Tq3xbSmL8a9Y/Iv2n+Ligcx+aQQ2ffjii/YclB3lr75vpXMOoXAv9CY4WcUYvDrdC
cDR0F2Uxmg8NJAfe2uKz14iA9AhagxIPUouCRtwysNNTMUKbnE5ahrnqBHiio+U0s4om9ukwB7DB
8ptgk3puAXymKM6UB2hOOBJAJuDCpjKgRlRpdIr5o9aAfaU4Sw5fL7m8Vd/wIiZ2PqO5LI956RM6
UVXFjVPRdGpQsnu83AsQ1nYqdMLNHgudtrtZ96FKtTJkYB86t4Y/SEnuSPviZhmc1XI9UkMcEa8B
mdzOJCZBQDdFTW6ctc6KZaogSaFm5mK2+pesa7myI6vPg5ktCx49pEeNJF4FoaKVM5HO0c6XZfGB
nMnscN3C8ht11NDwaRHCa1ybbCACa/3g6oXQq8rU2fm698Mkd/virzisz+iJqsSrkpuul8Ofrvex
y7/mpmHW6qbs82ELc3ccp+m+mswTO1Fei4pW9kPmdG/gNnBPfmyCwVKV0WgrZlz4q8oIO5+Elofl
sFWbWOWNJi2ol1DlowLs/l6wJaG5vBC/UJyuVJux9W/FSVDtA42e/1M+HYQ6bgtk2dVOAmWsLtnT
W28wQKdGGnHvGRvuYGpSXFGpn0WWEn5wYy9ZmsHkbFCZCQwwWPUA+32TSWbWp+skSxttDm7fSVBB
aHks2S4B2s60ekFTUMYuRac+3A/UbDD+8tHKssiBZYTIY2yUfwWqEmYWZnWtdPhPGM9dkKyctFoO
GIfnag4JSM+h3JoK9I9dvZ6pRQFTt+XvzKmhK8dGmwXfh6PCxojdZFQbw61DFnrlL/y6je4jQV4Q
QlBZP7h3ccqI6DrS54CbavS/TqgP5p2hBiyKyz7q4UfQBPnOW48PFhMkamZ9IQDzzUC//PWjvgtS
sJ+eqaTvp27ugVO90rm1rJFpqcTOkFBwPvWLs+qF9Sr+FWoOUnu1HxKla2K4wobK/CcZTzkDlkg/
nx+Ax4JrcjnLVvolbFAfEMMwIi2YUFywKvzcFWi2p5CZRCtg7MT6cvtvQMZt84YZ5EXCLtgDHR4k
2ydpmL7YBhmCExLvr/hTs6JhW91wepDw7fNQXGn8WVVeeK3oVI4I5sBzCakztXILE5l/SbeTj6YV
6E4pmcXNTgnW/0I7PiQbRzzJbpk0Cs3DdcDTOEz2wJLVw6YAGxI5eNzYk/wcM35le4YjO0hglLpa
Zc+DP4FAHD/GB1gQzuvntUmKWG3PTtIUN27quBlTG8m4w6ZXS2JsPGnRh0/5K/Od9/0TfO6GgFON
kbE2cAM/nQvtgGfoeu5emNwHDg95YHCmp4dJWiOjM+N7wrLk/ukxkiNEA11/9IeSDzamjHCu4i8H
lA1B7QriMDAhAKgqTb9Y+KntiIKbtMAOBRgx/D9CbnVnb50u2lTN1THe/gArGM/tyAECyHnw/2VF
xv2pU2P81DyyNijeJoYKhrwKoh8uTldoDfDPQJCStIjOzM5Ncz5hy3783IpohtNMitLmCcaRdOim
FtIHr8tpCy/79K4bZZ18FQMlut46c5QY2jX10oXERa6X+X5wCuNfHDyNgi/4bR7qxH/aOAFrHPjC
JVLKq01yFaJnpaq9YZM3r7a/Dc2PYBX/DG9UnTgcf78cJPF/Kj+wPhgz/1GCskt6hReMkmke71Eq
a8/Uavxl/itgj3JPFGoFMCHPE91BEJoPFERy26g6mrU9Y5E0j2i78wwy2cXxeTEtOhilE4s1QJXk
5vWN6k8LgqnzxC20Mlf0x+HFC5rxHSC15PV0ZICb8916D3/xg77bXCTpTkBDjMRS8Ha5Z5PGkKpy
HvAhZFiDV0qeXrHfmYqLJBJKUIR13cqay3K8iQvwt/MuyTU7p5o0RdIZ/qxrppdzdAiDVn0ntzNP
OvzOgHZzEYqsqSEOz/7vu0UUsAg/h1mNDu2SlH1M+nwXqFcU8KEuSN3mxt+3EuUSE/pKlLbVkPKZ
S2t4UuvjZ4lMcdmi811C2f7l7nJvH+A9sAZ1fEG2BMRwLI4GxIvaw1lnVhHtFNVtYCby50QqPEtA
JqFPSWpSY6dxxDeJAVX9YMFeSq7ByQ/j+qCSbZCJHfc968LIq2o6WgF+pfEU6QXDmxqcfz23arqM
Zw9IXEkDK5tNHUw90Jy+qpBk2HqhLvn6JVqtTmM/tGRMJgrUJs0rDsgCUcIpSGE5AehTqqjbzVY5
DMtj70LaBwYQSK9ynRGcI7UT8ZYnsBCZ6/GMxlsyXnasC6avhTr0bhzXDlWIBMy7dnZ6/h0k7Y5v
nj6vfBSvO12z9od5PFcpiDdAJ4HhqBk717xcnzcYJiGdFZwOmsn2NiFjnbWa/CoXusbzWTsAH9Wd
ltrDMjOITjoRRSGYmx9YSipNa8aVl2ENEBKkzmDArwI7n4/mZGdU/5mCOlx+9l2vPw71Q40HgeUQ
rG0DaGLPPrqGR1UxQd3NmR5YgNtiG+OyH2pqtDfLfOHm3qj7Rnrb6w5VMQ0+aDYRyR8PLcya9shG
KJEpHwLHA0LzM/M1sspSIBl//eprjCkx8m0lao9WnEDOxmfpwTAtFmypAwRuj6xu1it6rhHxUheo
T1yly5dnnDt4ZBPXQMF0WzjuaxAoStLMDmDjtC1u05de71CbZg51bp7S4YHwGsxz5N/3PdwWrXUh
nPmqAvVse65XEA0CCGQII5xFWuq6huKCZjXOdvl8KbtqJ9u/4+2tJcy8uYshIjsulwqeN5TMxuiZ
m8cDVHfdga0bK6cXrS3g911JaIFYJiiKKUXW3tvF+MO9U5WN50Kl9o1dBDNNJIbNqwXJ0HcsJPys
1gWnP08eayuvh1wknrOUkGpEeX9xPXECDL90Fbz3fOncfh92yEqaYBwzZkbn5tYULlrbkgxjYHXr
8VhComeLL1dcMzrgvzeSybMdd0HeKvBQHiK6QcnoNV9GWk0GjIwGZsRN0N7dU1yz4E5s/T1GCofu
MBojjL54/5dzcTj2wNsCiTRa4ry7sM8NpE0CzQEtsFhu9sJl/hb3L26J56kc+8EGjhuwQR+TRZ1O
HDtyV38vYtVWpzeW8uwVM8l2XpICY8KnbPG/roi2RYLRMI7ulfmGyR7SKcfsHBkhrN3pSGQe8j9r
xwk96gVVYj1/gatuXL9NwMJF4Q/Af3SH4wmtBGDZ1cyr1gjNpcfpKf1PiNbPJDkzs14Cs//RNWux
YwbaFSyHh1L/xHQ11QFoz7iK1GNdsICwlgS8yN1ERaYpXkgque7NunOHulpZ5qkuhMm5Ni7k3X4e
ZAFhvcOPO4trUKAgZV76LSe4Hj6vpEbXTSB3r6+R8HHvb+6pDkI9ZME3n3ttaSl2L2jjj3MZXdQp
nqePswWzPNt6vVnS5vhaIxGljFC1HZM2YpBfUb635hP+6drsy/a311P76U+U+Vq5OwofhN1Q5NN0
M5WV7BMhRHhbA2BkDYTqCOR3NlmcHUmKZEie3wzUEckcnHUkv5M2LkbkegeIvANlBt4Lqr9cE5Ie
Ait0ajRVNNvN1+twx2W9219ChV9IRXGA5t6bd8lK26W+UW0T46knc90pg2Esu0mBC9FSdAQUnlhn
TIRMtc3t5oEey7SXYYROMZ6UrAEc3TurirIpPgwLmC/E+7QBM0ayMjmTLruHWEL08BIHeKt2Cmq+
1ZuHNs3aZpXV1DYAyqob7ope/3OekOX48y5mDzejGnxsmYD4UcwDY0sG/9J/ppz4gdYm9iDX03IT
h7EGGmdOGIndqEmIepQlRrl09rSsbCTIFjaWGRe8Qhpa8eW5SEEmtoADocylnjaTCmc/aQRVUHYd
81Jwx51Rw2LlyXB7Vk6alhbY+U2vsvWO7NtMjO8feXQ7KEN9/5FxyDOw8aYzmkeSonJRISMkHXh2
7KEL2pVt4rJ2ltPmWIU53sYBq2UBoFDX5ZhSqRP3LSrp9PaaIgriBpPuF0yjjluZcRKlsVHOrTvK
DsWKZ50DcR6m9HnI5kl/9Bhb5Me9PMkl0QW2+pKLn4GHdQll/OALjqzrYRQ7lUF7WFs3Ju5OH2I4
Uh0XtAX6gAt6z857Dm7cWquthXdD3AFJ5gm5WvXBw/Ow+KzkwfjpPyGwOApq6ql0DXKZrPxiBU21
T0Swc0F8n6pj1P2PD0BWwQy4+gC3YdcXtYhPvM/5ORLz54kDR4Gynb9pOH6FDWRlxmO9KzG8HviS
MNzrMi7gV+XtUSpaU3/l609dSnnuIyqyC912EFQA4rOAmr6cfjNa7LMAR7qQThtgneAzGNbLUnnS
/TXar5Kx1x/VVCoqassx92paK5bhiOY4V1ksfJD0kVq18akFFoNrCy1IJwqQwNnLrOwng/B2FA+P
RtUIhhNone+SrkKezLB9L7iy6FqG9HMIVS0+XPHdu/udwSggTF4zBGVkBKeHoyuFNA8ZRRvnuZ40
1CWmKy0tIgvkfnZzRrgKfQ9skbN1bKJUefppQ4VajG53obYf3th/oUpPVExRffen8c4vbYIL/9/t
MCdzl339220d9esKaP3Co2ppfJuzUzU6Hl1xgFrQ1XwWTbQ+v65ihzlV2PID520mafxO6iXa41/M
Lb33UAGY+x5lkwJmLkWMMdW3/oEpRHzMrpLCP5KtC3UCw720PK/KtRklXuPobejeFlz67UPELHFZ
AjcFnaMMk9v01eRr/fpDlBU5tz1lDl2nW5QGLd9fJxToW3vOkoc1lb1LNRUNpvr8YkHPGY1G35RG
O+n0yFOfaDRAABLdx6peTAibIg8v42+aWMTneEjb8GscoW164M9fBy3lhkZNJx+RVGC7War1kInY
8hGbzgpRqBdpvPdWIPVEmMjeW/47hQuAvd6lciQYnj6p+RBk9Y2rFjD7s23mzwL5tf5fsHBUd2Dx
+VqE935s0MgAYWSyVEOFKXDJNIOdRGuIyCTqVo1B8TGuATixA4+7vI1TvIskG4NoyMIH97TI6tgB
CbCR5UEqSrkZPnle4Bx/Eu1Ce6xsukxDA96TkfS66QpTzDNHRORssQmSd+vdpXxMTY9KRdIDUhnM
sCbNdEARfx2pI78BjTbDGWazlKADLHKTc4+9235b1ut7ktJCuxK38Jn/+ePj7ZBktJucwmemefOz
AKH84kWnrxyL6eVgpbRRFEfY9BpeiUsFHDs1SYWmNwDNDQ370yST7yQm6/Z47E/wiIgl3poShAc7
7IN8MoaqWYQe9UqURqtEl8r3v2FtPmg+wMt8n+rP9Imx26oBeEToNTWnbnEJACMFMRhI0YMhXBJ4
N6mmERtTp4Z+tZIhbq2hnUSlRMKbLjbxeI4FUuNo57wqRlZjqmTebL/w54CkQtqotdzivggdu9f9
55u3XOKcDiYn/6z3uJSZGWkF1YfRFdKt3DDPB+ZaXSsP4NjqlQY8Bt4rM/NedXaP4K5DlundMEUM
FUMMi2Q8wkq5vrnWuI5EfmjwcTSyweUlMniM8H4T2zaQon3dz50soII8hAUH9S1v3+wyC2zsReq2
cl0omOWOnLylFDmUFHOxCENxwOacSG454MsTOz4nWHiWR723Zcjw7JOapc34bYSst+KBhBxgiGrT
alpncWmORTPBQ+aLPsG3tbjsyqb231CezLbWWH3QyUSYudLg5zXVLo/ObBAYKYJ4/v3AFZMYfriI
TGwCic00g1yS4/BC0Kj+IV0hm8FJjieHnjjeXWCmtliHJqY9CTQl8s7Gp4Btr+8nGS1FnmjiYyVO
JnSnlYOc140NcqRpof+FzBo99lFnyEsrI+fITgX/n51siIjzN3D+dgqxDlH5L2AnAWlvzZpluCSs
L8umOzvDSiSis2kVAY5vKcPvYu3Ehhg2uD3un8SoPo+4djohlof/a+H1rnNYBH5ADcj5QwQQpacM
0x5aXUnPTLJvsbtOY+ac9V4eF0a5mUa5tEG4YfMTTTdGP5DoGEJS+9CeSPCUINBPcHMFSz7f6aBz
kBUBGLnUG26bOeA2isoa3jWgRQDcshKfJMeoHpclzHyDZF9fBkvP3yBCuyYQqqLpIBJ4GLf375oy
5WLNsfExJjjhjfYKUMt9W53zex0gGpQwN//9115lXkJVoUkOO5e8VB1BXVTlUC6UmM7gZFcHNqYC
4KjpFcNx67W5K+rBC9O8lfFqtNjTxlc2Jb2rtfQA4FffEQ4zZlrd9VDtYJdGCAu/H3vLFnLJxuiM
WRfBWheXn13d/dDS2gTbC8S8lnxnKBGjX0VJ+5blbzRlMS7yv/z1cofxfAFUqpaphxCePbKgzA1e
egtzAIwOWkhyWwMs2UeIja6q98e2HVqBkPsA1ork4OyxDBo/4o+IANbbw3o8pJawC1+yT6kn520M
d/HJJGfxcgwyXnkOGZadmKtVEX+k7xKrt9sfrFn7mJljSLsKmsfHw5phz9M50z2rkp8vxwy17tMG
U0jmSSsvMSdtBXpKdn6xbF7AjsWLmcxi7dUg5bosQPzsOfgSfSORRX2uW9ByriyiAhWn8+Tjo6sg
3sisSX6pofk9WKbQOCmNj59BPiNjArjHFBGIbS4LQwAt9WsNhdTasb8wd6E/6IjbGF19EqASy4Mv
iLOZ+MdKS5KNpVmHE2Y0Uua/pGMPKjta45ngb9wRA5fW2+8HROe5QsfkuzS+At9VQm56uj6lGgxL
VIKMoJeL+iXEEIbFnIT/kExRM1UX/LOTznpZXN4DybC3ak21NyX9jaVrLyUdKz/WnBWpDuRimUji
UHKsHC7hDd8mmisolaOH/kY15CdY0eFhn6eCjdgMoQtfJmTOQ1UXuOf55wXl5QtVGGOEbvaHECXR
YwPncGVugH6cN8HwEzwfMQZz+1nVSRyYDG3uVks49KRRLWXYllIDprWnhu9S/X3EZunI04Ujt4kO
Cx1ZskBaVjVNTy4hDxrLfm78bn50T7/3dwrGDHWaSCnPfHP/jCgcWZEBbwYaD7R9gBBGzV/N2Avd
pdj/xRKgsIOxsfd45UFtw/V+X8p0fMfB8vFqkXFD1Uz8zQHuwMBWbB0DVG4JqSVY8Mq4BQExdLVZ
fzA8pAePM6rGoeJTC9XGxRaCRxMJF/HeQPtezaotHPwd5xYQp9v4NZcmtzdykqrJRFck9I2L1jac
5WrNzccLzVTtjW6vuWnES1QB8v397R8RW7hc9KJTcSlhTvp6hYh5TCaRRYv61F+D+X5dlXIvRzHD
Qm3XgEBYPxR0wqjOPpvtYuByNSAzmE0gjNcRjCr1WUreEX9gjpEL818iYZBRb28ecPBl/nyu4G56
vs9rG0CsmKUl9poPjaU36t0b8esoIhd/LBBZ1Ql8LkOmqGsFp+WbpeqpZYRs2CIMRS8U3+KNIkcV
KQ+j1h4SVVZ5eu4PaPVWN/XN0JXhFXYJk7kyjmlvkfdG3NlTpSr0rStgeBelYG5HsGVai8opOi/+
NYKArtOfDmJ4yVxbT1jh1I60ndJRTinN3yh4uYh7Qz9/639DLc+DB825n6zHLmlfwst3klmxRS6B
ulbqASbqAjd0OXK+fim2DrK6ZpF2UiANb0l94U2Qp4VRPFUmra7Y9cc63BALNCx43huSFC5jgMpN
ojQcLbgY+76wI/QRLX19mUb11z8Y4pbQdVtMrcCmOxC5mRBRpZYk0bqdZSBt2bHHWz6UnBCy2U2d
YZ79iwtw9nmgk+2ush74aEfSZZZ8/uAkGJlwZSWeI+hi8O+j9/oSAnNGQHGH7uaoGy4XR+okQmDU
hhZ35XXn8AU1av21HWolQptdVU/3h5+7uF5m6ebfwnCjz3dftBmxni405ISJCeOe+OIMKUzD/nug
pkaP3cB2Dudj9qvO/skqp0bscQ8XKYZMu3Gr21l0YQb0oUrm2eMtxSM3hP0R0eUNOuq3Fu0FKkCn
U87+P6v5xZfLk6QzG0Dp2ScK+a/pCL6ib6vuh2NK/GhKrePpwnZSl/bzlzwRBHd5jldNwc/IJZi8
XZf2d36OZFPvbTecOiI6DpEa9Dt2yT55+7ivF/bdhsqBCnbRNnAs2lM8nj3U9PpUAFsfqBzQFw9r
ZuF4Y/yXDuMVle9ybWBXqW2tgUQlIXh2+dF8Hxz8bWCmjmokdWf1dOT+vdnZGs6+FZi2fQlkBlOs
dkjoi5OdT+ETzxRV189EwKxEGl5UZi6fqNTdaPGKemwq6f6BHVVuZsC2TAIH4obOfBfkWqMS+gqv
eKZbRX0LFYogGHjW0jYtgANvlsXYWH4oIjNBXlsYzTBYkjMcVLOHDYFbnwCk3hk1YwOLvXZvK4XY
iljnMfHJdRJWCgu1b8FDuKuSG/Kvc7QxU+htNlFEHTVjiCb047XyEYVSvjqGnwXet7G5LrFXKk0N
Nf4AIF56At0/md0VdErjPmEBodDnaMTD7f+/LaBO/jiYgrvC3p8Xv+IFI/OTD5toVCkNmrXy2/kU
TpqFCZEebbCrLbTZCxuNwsRtwTocz8jtYw+ixHuHx+AfiS6Xv1eriIWDl7tKUY3FeZdWHtzrKerJ
VCOflWbccKYl8l9YsmkqzMQQf7nu2hI3ei8zIqi+whfMwF03Yp9Wl8GnPcBYgK7axTr/J9LKGtUt
gkXbQBxzz8zQU1m6bvnHZkhYikTyCKGeE4oUe0DZv2KZJG6VgzY/T5OnJswWMXNbT4/5LTDQ4TxV
Z+eGNirIOuHTbg6D8fL84DAWwGIoJGbJuV4i+2h2czXC4/EwCKjps9YB02wWyIlovLLopR6EPRBO
kIkO77gPRfh8QbokrIX7+puq9LwjLzZGtbmh6FpaKKVukj4n1P6E7sqBQ717W6UHVXz3EWM0EbUY
1Qk/8WvW3gJyebUVWzObPB46AQ8qtrsF0aHR9BEgUcKUDaQbr9ND6tTWqlXLmG97zDJM60hffAS3
s9IyCjX1wAUtXC9xYcPtsecX04ov4/wZbNnbBPfvE3RWEfX9n6JLnS3fynSl2gTywu6hrlmYCoh9
fzYJbIvqu/XNogy0RixF+vM2cZKbx4TzlKejjoKGVKDV3OFceZS6CNBO9LmqrzQkaJB0xBnunT7f
YKBq2g7Qik63QKWFGdEaKNVeckvijZV39Df7ua/wZnC42y8R2hQI66A3RmLw4NTCTjnM/mFH4IMG
pD/6LLaEOI5gspJPoKZMoT3caTezcWL6oQbEea3LeuGXszwCFrVGg0G+1m65PVMkYVhQ4tmYoAie
c+hjkzc3n7T0ZoWnkBBjWgbG9cTcZxBLwN9YiOe9+W/Vs7gbSD4TzwLztg5nbractYLEXpeuDXUi
GiSvl7ZkpIisyHK/bjw2rHcOio8p/onhT14aelIaOPfWSZ3xjnvTLdo3EyUo+LTfqDEKENC28r9f
CzSd94/7b1R+FMgaV0Ch07SZBbDzf3uPy2wo1KC5UDA5ZMxRlatCKRVo2l+brTTCtd7VXCGYjWhc
7JOrlutMRQjtqyD7anqWEZJM1s/Y3VAqDOUq4to4io5cwPGbx+AghpFCRXWIr2yAPN+p0MOSHUIg
+WMFPMw1Tt+vX5AXrdHrFWkfCTBi1M9/yz52MXBGtfDAaoxhY549zPRnK3PyAq6PbqtX5eNxwSoH
LEZrD8YXeBCuociYQO1lfeYcWynLWG3hIfcspW2Wna4prCCq93FaqcA/n6GDRryS/PY4DKkvNw8u
XJ+wbVu0bftKtZHVuJORnmQ8sdQwxIGtgM9ixM8rSxuZJpNjJ0GWzYYgHI6SK3QBlxc43MCvUkSy
u63L1nfdfW3ng+jDUdbMMUnyb5xmGWeRR4lCHfcqXKbLuNo43lAWQ+gzsrEevLkCrkiKv6YtUdGc
KOnRS7joqNINqlK1W/uBH+4ms+fe8yRErDZhfB6GD53ZwICt6gpwMYdITfIw1P5sE5wKPO0besjk
ZQVo/MYhvPwpyt3lVCJJQvD+tILqxg2Ngtd0bMvknZCmOImPeP2k4mACi0CHPt8wZ1bcIOgSg5g2
beBxJFMe+KV3OkY7Ogum8A0gB2DGmZCbZwJ2duhh0v8VcK6EtZzYYXRO6RsipytDfcoamgpH51N9
ocrEHo9rzWnJ0Hwt0Xy4Ip71vvo0xBdRRfaqqb3+TwXaIMGJXz0dtutdWVu8C4rWpElW5q4eiYY0
KJoQ2meeKOkrdm+xKvE8CL9vqqWPFb89EpE9zmBKUB95k3tj7lESc8+FpIaCMBbUL1oQ/tmB6qZ5
5QMcrpYE4s0o1rl0jVm6Ypp8b49KX1zBTGC28VwzuZQ/htjhwfP78xsMlA7cxvNZkPM/etY09iFH
Bl+CidD/GXIGOeYxrqP9VlVkImPBx8hwNhS3X18BET1K+vkXWYoUECJMrBizNrqJPjkQRvfOYHJ7
gBTBQfEgCaucdoBscyHkmWKP3J3cGYTLwiKUDzs0rR8yNQkTanea0Gas6e8nS1zuHOWwaPj7q9f2
ByXYSnNrghOKM580uY6m4/211kz7FmJY+QCZXs/4AWehTHKP5tdxvsDB/CNc8oIw+zHmEeHXAF48
Oy06cnNtNZkENxjvnZD45TuptHn5P6tkKbxf79Hzsqq9Kx7GklBLJgzX5eO1KIh3/uHDpMvFUZeP
FLlIjsAvIP86dLigXoHY4xbyKP8XGLDdJrbwIFBlgG5bNtWE/R3h9PwXnPS0rsLojrODiuFlxjQa
W0VuDN/8dT0TnsTxHNx7MJ6l5qVYgPKO5PZVKeH44KdxitZBecw0xmJ7jn1folBqfro4Aj4ABIkm
HIw/bJSN1fO5v036CgL+uqs+LhjFMHdk2ZXDbEvL/QdSdWpEkkeJwVUco0elfpOS1s+qrUYrnX4B
q6F6465FCDjk4RRDts7sH0CJArCCpJdd/91YNL35jdhi+rmkXOgMqa8cX0phXRe2Jb0niYurssvZ
d7hmIx2YpcxiHrpHg1AFNj8Q7B6JvvPAOZE6PPgE306RfhSJlAy8RJ2OgTG4MufgaG/B+S2jcmgd
Uek14Djqchvd4ifJa5jekkLLy4VJ9/iDiFZK3CzL2dbhKtdxZcUD3MK+li1UUXOlKfBffO7DMygw
pPERuStlWvBDlkdNJurBLK0Oft6DzcTVDFG8f6pFui5svkM0QoIrR4QIzNT6DJyQAZDyenfVX9Qt
Zfa/GpqLE1mZunGWxvSnsksBQBSnHTpbtD+fz2EJgb9JCtljEQ/yK79uNVB+rHD80Fmynb6oOiVR
brnnS2lPj8s7KU+FRXy0pTOvEz/zvSZCf7lvxrFwVaWjsf08SrDYPyGlP5BvOmYe1oODho55KeQQ
olA2DtKyWqPnxr5HBL702waiyPnr3c5XRYVI+ReVTDq8sj+WYGCSaLOmVuOOgFmwfXyZeqGGvQJN
kK/40z8IGEZyR22tEQtsnqW0wrsvcG/WIZaRxPJsIC7AyvwfIfjq4aCJeZ1dnnxR9VKycaRPN+nq
t/FdKWFtXu0RcrKL9XjReuDNzXkZcfSdWH5hjR6yrtJ4T6vJ1eQBOPsI71z7h5DXAQk2wYCWI+Lu
3DfYqeldVhyBAcmQTLV0V/SKt2lKccPCyK/ITDOM6EO/YVl98GCrG80fdus3MRlBU0fkel1NTTV5
yHf5Mh8GGK8TYb4M0s/brfIT9ffguCFzug1wblFgaEB/YvaF0CYfRHfzrs6eLV+N9SSdQxSZJV/p
oKejQi5QuXMjJek+I6HdrwO5V5lHLU70Fs85ZP/oUdy4UCYQhAjcLvS+CXQWmrJSRksmTvlLBdYB
C341E95BrfxMDpb8SecbNhtROLnhmj4YMR3xPawh5WcaKCkn9cRdnT5D9NBq/R2mRmylD70fRVuq
9/83HFdzi60J4XQOMEQ3wE2kb0xJMvO+yUJUPQB8vGL4gyIGgw9vcnCND5wkQv6qaLFX/bpDRavM
ANnxo7x6iZ4hIzFJEXNTEm2jQLbc9aHrQAGpidiS05qmHvFUzrzV7hrsTqBqHhPT1xQ6LY0RP6MI
R6tx9Su7995O588lzv5+MzcUm8z0IearCkJsedMXrOA16GPvr4AoEzPHg+O4opP09CYwWFuAziEQ
r0vwzb81KNFo6fx6GrG3HJgH7yfMDD2dBGZnxs7MLGMDKd9SLmHE8MYrRgJEKrihxUW2KZq7ognD
8nd/OlItlvneVAitbJFZMplowMvY/QzVsJX2bPqUV74MzZv/3hzrCPX58mtz66Z5QKBD4Hl9Vmr2
ExuIbZ38UO8LkxUs9Iz53EKuh50UiSj8himAWkxJrBZuQYRLFm5I5qkBBZMZg85HDNsDInlLQKbU
lucqVZlYCrvzcqOJQh947UsfkENLeGVNCtR+AUDu6wrYhX9T/X2VGunf/cqi5Pl0TC4rWo5a412j
NXrM6KvtimOC0dGAD9yDs70tbrQb7KegFYiDYbkI67Q4f1UWpFkpiN0XfoeDQl5pBASbFhNFr2Cr
2IvqO3L0u/tI2PXgQp2tC74miZQHz/Xa+YbqV0ftefNXfrFAnSUo/ccO5hVpggKU3aAwHuo6jaUk
d9bvO1tBhJM5p1wgg5YRoKws7W7BT76DEmLE6ElqppxZLnPlO8dtlwlfDrvmZs+Rcsnszx2aiKyi
xrVI7iYKbYis4L+nnl9r4JNS+6jIb3AN9ugnNdqG8H9vR305mAN38OivGza917mzsUSMUcc/uCi7
Tt2tYA2ojpxLUHAZFRrfr2oCENx8Ep0Y/G/JHZ+Dk+Hxo0oJ+7bwZtCmHAUfvIkdydt7eNsrVm6l
A7h9VTiJM3Eo67JXG2tdvi7j6e5wS358/tCFxlwjiIHIzftwiBtD4uPovpuPMscxIZ5kWhXkaAkz
O3GFPjs72gBqeu0DlpLTrHU7xjGUmKvZpBdupxfLPmmw2EwjtZCYYRmVyREu5f7tROwCDjkrH15r
eDN2d/n+glmYcsi/05avoyt6cIE1LYE3Dguuix0Ki+MhnrJeSlTQ9OrR0sqyJBtDmY53SdH8wI0L
KH84lGp/c6oJZ4MXTGeAofjjcCQ+Cjbmz1HbLfp2RG7Flty1fk27rZv7Rm0tAUCk9IwJPoZLatDR
vgxYgPhlyIctHWmuHQVQ1bBOyZ7Z8D3Ncibxd0t1uLLpQbh400kJ8r1nbgor6hicrRrHYBDb978K
+SZzccT79Lq7neMPJiHj65ulbr4LOALfQsMEeo619TMpp5q9o9sfAAgn6nzBaXmfTXU9r5t9hav8
yp46XRdfzxidbkHnwHnxjj6hSSIFKS3Ya955oLpXfFNtOUfKIvcr2qm7zXBiNE3zZQvY7xAD9161
7NVF3z/biNkGSfQ9bX7WHI6OkvhEvkp8ZB0/nMr2StltJyixi0h2+k5GdhXudY6XZ639m2EchQ1o
30s1A+LpJeaCmJHhE1oXwdcWPx8xnehNvmbm2hPiRk1aG9DVQlYR1JdbTyvAJRQpWliRU1VMy3iW
7pHgUoLuRc+mPJiQJsaR7XrGWTv3V6NGzOmt2ZZmCaPEjCSq/sI3CLjIVwIlN6kVUxYm6T9Mw8ok
lbAk+fkwafFTrND1qNL3Mzdu61B6MjehrKCEkZ1ZfVCkWYOJ86t/ssGx8NFxp0uvQxqHJQifbgUB
qcxg6he5iaaeG1hRv7AOaj7FGl6bbQH5eg0XVUN8DcLTlBH2L7JiIfVCCg3L+3iYLwRsF54mKejF
hkgjAroJFVgV/X3ym5Dume5H33ZnHO85BsgjqonhqlaiDFHF9KJlRhh2g/PGAJ97Gl3y0jzlQLiG
pkDnMaxOV5ekAx0OS+QeeeMLvj+wX0+Ehn6f47aPpvi0A8g1vSYp5Obk1z+3SIg2UpWrfVIdcHpZ
7SwNSoJsY8l6t8mUrQGWyJcYwciRS65VmI8bdv3R6u1kPR+aBIO5Ob+deuqmbabA0ZXVoSKFyMqz
1gM5Nhd3OQSQvIJ8AlwqCPWcaRyj4r9CJGxbBB8L4DcuEamOEJ7kBoq8VuB16ooc+vxbtHIoekdJ
oEabh1/RXjYWEfi5n81874xXv8/S2FKu8Id07YliGIyNEVBu8h0j4KR4klis6TSkwqMvacL9NJg0
0hBBGwhWpv6HH3XSBEDCBy/BCmYCFewtugtiJbi1QrDmnCN78a78pqB4F8G7rTJrehXQLdSJeW5y
UVV801/sWuZU6o4kP/pkqIXxz8BUEIP4pjKXVSi8BUCUFnfJhuNK4pozEfb89rye0LNhKwn+Wh4D
Qumd23j+OMZEf6x/OnTDPmM5xfx6LYf+rfaAOo1SFTqYi7AGaiilM9CubiWmr7ioyVZ80wA1UcFs
eOWVMEuq/zcahfdFyaomJq3ix0bUkSdqYKsffslrlUu8o3KivxQdeGntYTcbUotRamFNQUwudD/q
ZeJ8WeeoFBf1BPhYfZVZJhjjYKBfpQHHV5TlfGq1hhvWQ0idYYhqSauD/AAlLr2dX7gaEX9pg2O6
J4T/yQJ+M+p/c5IQ8Lzgp7E57+6Uj5hjAI7d1FAlR54Vzbufq+kaen8c4cdnvVf5oLBoP9UPEvab
TffU1/rAkhMnDMFSi4q2dWb7gV7hXJkv/66xvzKXGND+8ZKF32JyW2Waq3An1QPPjaoDQwQvcK2M
e0rHYmiZtmGOCyHo5NzR0YfTVjFcLskNUOhdkQEFM7TmGozafUpH3SETGX+mKbTcJzKAKaZlxIcH
yu7IpuirIFdq47uSGeJr+hw3R9yXT4ANsjpJGdP/p4bW1EwPO+fEFka9zkbBjuudP713IZX2+7Kr
O9/wWQC7Hk09gqNZVG3r9SeBKs/nNhe4id56v0lpFztn+pB7SEBBsL+5dQ1pNXiOWW6VegnxnOPQ
ZB5Sx3FFuaK3nbVbBG/5A86R65OxK876wCKnyRpL3XyDtotlsLWYP9Cq5ElBlClsdRCvjx3mmk/H
zYfP0Zv0xYDqNbPmIoNyx7y2O+hNJDJecztaDt5iBw31K1MD34igjrT4LGSSz7yDqyzIcH2vUXa8
TY3XS2D6Tp5UWDbrhLtsCuH4OxL0MXmYKq5f05huiqiN+gsbzeRUO8ncgX4KM+wk+KQ7CXRyk3Jr
tw/NDf1++CA8IAZx+4hAL+QPEyh8im7QBc7PuHhHXzESQ4GPQ26e2X0Fj6OrNfhFP9d5MaxsajdA
gLECAye3U2w9LaW+zcmRt1btfYHr5+u7oppA1tZoXkWnM1awjaCQ3TjybUllu0zEfv/eDymyY95y
MOpmBLaM7P12cI3c4jXnrsQf4rrUmZRZE4zsP6uvIK0+fN4ITgHbZxHljQWh59uXaY4x/vluTM6r
EpZItunEEyqgFxCCBJPvwiPDO2hjW8QSL7HyYrw5SsVUoEQlwoqbYsxEtJDZSOghikrq2jxLi2df
T7jCxOEWH9jD4TWgaP8BQTjP1RZ7tV10xBoSCMkNyE4BBiwGxgTy/Gg+GS7KQc16cXESggzbyIPz
M6kIKrPdHBTbhoOdACgog961XxNGDWiIK8CwXCDCkbgDzGDiWgCJWFBQfta4ox4DEOnjR/Mq3W5Z
+7RSXy5bDOGqvmIVVfvzLUbd0grRpeAognlUGzSupjBucInXf7j6UYCJCcXBP4FEjpK8GhIVEE9M
o/TIxuP/rWzfdzuJJM9e+XbPVMyfmY5oGrqbxaF40D00raPUju3Fn3lUKVOgNoERhROAkBRMVgFq
fBir7fYpHWooWymd5dxSgbixTUVcHnT1KLQO7VbMVYMTqUk84jh71p2Eyyn2IfEkt+4WxFPCHoeT
UyKtEeWMxq2L0lJJOW0SfLC1bcYgE88CYvAHW3NVQ9ZaI6haaTrR0Mov0b1gB3gRun0RHy4AT+4H
LS2n8uNt4v5+ix/FhPTN3YDE+MDQybay1F3yqoZcI/+B90oraIf/3eqB/zO3rQIZQJPV0+retUFI
yR47JJf4a3eillc3We/WygcUm+W0TCvuy3gFSjQbPJHFqU090zM4KwJ32HnT5MBJIA1MCj6Vh7S8
I6CQi/3pDoJS8SGZ/ZmgJG45mx5vbxKJojaQgQ898wh/2UTioPXUqc6F9X5EYAVHuNHOFnpdpjJ8
GIhz2Vja83is3TpNjD90pIegSMRixMtEDaZLKuzm/tpQ1liwTHV7AWh73qyj0CA33K0wX45GyH9U
7iDODvntalBc5cRQL/BWYJ+XGC7Ui4Fgp3801lXwSOIDYQLESN3OlTi1pmHrroZ+jI4BQ3/lctj9
inHoueLNNtVSSLDD//m31oHiHDoN4jPaswW/ghAjbANUPVBkI74xUxRTRDuXOoBhGovJ5NNK0LwZ
f2cx/RJVRmS7mlhX0B98XkKJU9ecDxo2s0xkOL4alKVrPwzLCIjxpQXxx9XgZ+PIXIL5Y2h5/QKX
YsciWASxJAoU4UBWtGefbBM1r6VYFM5xVvN4Ty/Pn6TusuXPNyylXdQ98wZ7u5p95XWv0oovGz7D
JSJAwv691xfBTUXv8dIlpjb3VvCQFBqAe7SLacrwkgrXmOHg8JPKzMMX+Jm6DIXRn5XmQwsw+Egv
9646O0CYqLJGhyLUsPYHLol0wGg32CrlLRHwL63sr+pxz2+H0JHaJILXmb69IKNstJtaxxeedO/d
yZh2GRz9AqnC7Sr7raE/4ox2+4M7T78/GTIQ0FolrieMFW1BZICzniOsl8kVbwuCgEZcfJg+L1kW
ExUI8m6G2ukNN1g0eMq1mbYtUSVV8Maxs37r/8KUtg5E8/WaF1CswtdjLYCDfrYfZPTJny2M+ORq
hXT51+FFDsHJkT5LRJTkjfWDQWF6V0v+xTl+YKHCTFkGHegw5zEOY8RIgxF2GMfzo1lDp0/y2TLK
/LmutR4SS78mbhKH+0CFupY9iGXNJBx98O6pQn3kmJyL03vyVGXqi0vy/NEbEE4r2SbM2/ZI/6SE
XRxv+WMVvnCwWEk6C0rPV0N46cRKCX8Q3ozU70QaBORdMa1B4Ex3WLCrkYF92vB2sK2q2+oR+eMa
IR2+f4jykbT64B+fps6MjB28XV0Be/w3GArh/uotyAqlaJXm6DkZApdRhSZwQiXbdNVR0X5S0bSh
Y4S2iZt0pu9b5WUKNPIgesjg+XhPQyIvetND8f22hpSuui/MbrGmNu5DMLC/K5d5YNIxJZv1tCax
iQWWePvk1mhOj2LOkOHHWvA7KIZ8Cb/mp+d0aHiP9hsy6WVgLDA+YL4+mGM+leiRWWez0uKdLJsF
o8yMXYdS2BushTyNfNyl89sSPjFx6ous3yh0bA3rtlpUcnf84jErVWSEga2a7s+Oknl96VpQGojW
vEvdN5DErifp0b2HuzaLTKN304FbYY1NWJF6tfAu6xO2slRx1+u8lCojFlS1OHpDwYo8DNNdLSzq
UITAn0kEuqsae5GaWnQ07dGt7p2bh6ei05xz9WR7C/5TZ9dt0Pbo5P+Bh9qfnfqLIIJtkEqOXPIl
m908uf8Un+mc5hsVHNTHQ0GN6REP7HuET+M+XpLI5XcB2/qsTUauvlSOjLtN2QZl+7r7U4IBVva4
1QpvOa11iLM/5FC0d4tCC5AREOqcTmWyqdD0zsz5drc2qlpJG6YLgspOUe+mjwvArXTdhqT9AtGS
1G3q6fT+hywxH7o0NFe+LaOqIZVjlK9Op2MAGWRu1LBAeKmseM3Ad5fTitrnYCnS261ICgxxUf7U
xnLK/wrWXO3x04lKTFP74+Vf93jeiSdtYslWh4MSY8tOLhfoy6OcANguIAk2ryZ1BK5YifWzrxII
d42KUHGiowKqF8ElYBnToAOQJD+SXGubMQ013Uo5J38y1Mg2+YjDsfAv15g1en7P4zOmzctjx/oc
A9vvlXR55kqrwpm8jt2Xzk/AKofC79HBkAfE6jeuERVjw6So3AkpcyAsoHnFlp8JR8rrCPk3GJ5r
UnIqJv+6PSkZlX8/+HSan19l4edS+SKhmbduCFQt1h47Fv8lEGBiAbs93AO/8FUTRZMnMKiliW3t
JLc3IOZwjQb+RjYaZVmBHdu+YWkEPANI9eTFtABMk2clPgJwPMxT0H9ed8FbLzjT9Jkbs2tO8OxG
rl09fED1hjZ9Hd/hUExAcjQdDBYTZoUy8a0G5JI/xbiy4YKErT4376fGxgQ1B1tuvkScyVPN43n/
8AkFKZBkLBXa748XqE6h5/+/Fa/gi9Lq1LIuuumbcnxOvFDLgKFKPXmHzrnFezNee7GckpHPHIJ9
peZrWnnIiegxEktFuf+a3mFblN0LQeLDm0Nzlsx76S1KrxBKtY9jgCusKOUOEM1lys/sP96eWueM
Zpgy5JHgrF+PmMZUxOlgWOKJNPxVDFSrb5oMpGTyr4wbRH5yg/221q44Cxy6x9zcahSfkA19Cmp/
S30oSAzY6OvPz1Lns5A/ROpvDxMULCwNNY4h559GxCk1RRO3ygnZmNzVCCS+3niKJ5iEPJZJHyfW
eQ4qwel4Jdwauox9WiellPlWKfnfl+i4sXM4nHuSyAkWQYnYfIbNDvWkI+UcN4YEUpWoOG63edXA
kPvA2HKypV06EkmWcEWS0bYvRFnoKgApYZp7fxNz0UPGDJuJbt9KMTTlXxrd6F8c2dBdfIqsh4xH
DQti/FwiHh27ZOax/Lh1+FpcRL7PzAgAfpm/uetM9eRt8SG2SfayVlAz9Ld1OKY8jmCWrzn3l6Bu
8XHlIDmBV8woUYcFMOLxLN2fxLWz+ZOS+mHPxEjVfG9Rn35hD7VuCOkCtKW+qcFBdY924CPT56d5
vo0i0tPWcSbC1hoirsrYipJPn6IcLuKKaN+QwSJCGs/m+rDGbC0GnmY/Q/8hiCJV5lr3XdPS4nKE
P2i33LFGTDfwFI7cYOiB+8H69oSGzLZcefqLZPEP/VQd0lONlxdiziYyjnRoKP+PmkU7abUmSDOq
ZyZiwxNpW5LyuQRu+gvKkQjx75n4QCDhnOygpSwZrIczLyB/Jo3ajCw2zrDkPIeoVQouGwZbIfO3
Yetf2yjghVClQwiJ/VC5ZkUWh+upd4OmFEuhdn9mfu7TTNYGCdpsClNsLOllhL26n7h8Vo47zQhp
jS9+5CaudtDiJyGoCNY1dakJgBzsc73a0DNZAFnybzUGHmTc9w1P66aSDu5xsghA5bwQbYl51pRI
AhpEMnwdry+JAmyn0AGjrk6wjH51kMXNWfwas9REoZmjKJ+X63AGrjj6o2YIrSzgXDrX290gGfht
nrbSM5lpyG4WbueKNeXcb9JFJSq3aOGkL1CYRh7IbS8gM5IPJhdJxYDmFZwwnaMpPKz50xE7FIci
ueQqybrIDHMWa0xUsW4UsqqFCCRYMOst3hleEJeFtBQRFGju/Of0HGXTJgQeVSuQ5gxGf3E7QUKp
tX4IbH1HY10/q1dADk2I1lW6colnpG9/DAEpVdgIuG9+Msblpjj7Fjt0Wn9K8oE7CoEqkC0g394V
1xAvBP6i1UsR+U0HyY7t6nvsyiY6sB7MQ1qvUbgMqxAofF7g8Y7fFhZ5oOHok20gB84iXmbnT2p/
OHNu5cp2HNg02dOqZkkwsH6tJCIRDFSYpyokiHDJIy58DEWx27PGllnyrtZxMMXqbhdN02RLiLJA
NIzU9H79Ys0p3kZ4el178ZM+iGRzysSfVyLFjRPkkG0+RdUfNPHw/2GZJcrhBVIj5/K5E57XtnTu
V/pSQ7NUM9pEda1DNDRUJfveorauBbSyREsiLOmD6GkfDx3CP6n+iXqoPGKQ1NaCxMCf9NfBkFi3
JsDyS+L6KQwhnC1Ntme/lgCP+r38iaT60SOKXaNZx3NQ4JBboA9JGnCfilM5q1Qxl5R7DDgWmnht
l78/4byd96E9/KNN86Ik5VcPLu06F4JLs3SJuUJp5zakRjA7XXoe/AkzwOQcyx2o9WNmaqjRcChe
oRqBbYOJiZkA9l/xz/nt4vMoK4V8PsUpP1SuPPIO2Bb1XMbnBEDiAeERCsJ2mltChsWqxZBMFsNK
Nlinx78wWHyiyjhw+yzv1zyAv1C4fJTUmgP+e8lLQvZdqtibwsStaUqcTUn7DxF3WJfcEskNAY+I
TgVNbAZAtrdipETav3YNhj7LxUlfy0vwX4cOCvfNphm5a+tBeTxyVIc7hHxnPddMU5aCbLbnRUT4
CVRlrfyc8dnuTVb0K4dvO55gwAOFfiMlUCWj+zUdYKK8Viq2/7rtwhKZN3qPGOMqvIiEcahSLiqn
NINJJs+q8rdBtrVyXskMK9vEcEwLuxYXs3cz30okmfLZAjUMCACsOuZaCig2E0Q2yrWa4flJp4om
swtLR4ov+7GddMkbeshJ77iagYqNoKwcmXHEzjkHeIDBC/4PxzuRhIzyzc6HiJXgxMgRxq28eZO0
UAbMOx6wRUQ1RnMIuT8zhl2OjLtbK7HIvPSpKZb30HOLQJhDX8CXIj/Xr69hNxxAxMh07CgMqd7C
49P+HvYuOjmOBF+K4aMBsabEmtJTSPl5EJMuSWKF7vIGlNTNb6TY/X8i3kqK3ZaN7Y3GE9yRsEdX
IDcAbomQTr/3nCpQUn9rFfH9Gxbw1TWedxHc7T/pAr984ImSgoTOXOGbZHaY4dIUPkc8C4luqW7d
5NRVx6DWaSkr67I15kf4asGccRIFNiesmLRwna4TNVoWFwZd9VlY/AVSUealI4ruiFnsz4QOidjA
kRzv6pcpxGSRpzuLIZkqfsGQBvjsRtwB0S8RmedrB5gF91zSotRzItwMl+y8fgTNb69GTiDzKbg8
e72i/cZK4wZmVIDkgF275T3hqxdWyvD6LJOHgNdO5hneXKYkyB8e0acum78YbrwU9ftroQ63u61S
Q/rY3JxD9gcjRBgGOaFsLZpAu8gbcrfF+obHT3AghNIu2t6MSbCETbtrkD6JpHOkLzFmLavUNZHi
aQwBkFvfLRI365151PmSLUZAGkZJo5VgW2qDEcRHoc/ZGB+lLLE7hPVPO1eqvxJBkirFDsb2JE/E
aOeFvl5QrDlUcW4bftFULNANURubjjYxBtKm596Z5TuM4ZMJAdFYadiCItPLm28SowIIYGz6VvI1
y9IVvdJCMd7LyPekTRFZ5sdMluuTM41xaonHVKKFD7EcGQBPeThotCumu3ZOkl9puNh5vlCZo3Aa
5GQjaoYNLQTZlfKp8pxdUdUOWOeDytbV2HHj0Qd4Ivtt53CJPPezrEyQn49bKWjwOvGMUpGsnh1T
ZibT7LkxJhNVZHcRSE1k/A7XFVmpRvIGDsTCAZkaPJSYDG9W+nkn3BVpime3w4+o/9ZFLV+SBqKN
CiQj/aknPyYg3TcYt83yEJzb1LTFfxg0Vr828wStf9rdLZWDi7ZR/GISxAcMBLzHOM1NZTth/U9Z
8noEofH3yGwhCjsZhPRTXmOACyl3189fIdW/WslzjAd+JOVzTO4j70Lgz46mN0jMwOmRG6cB98B/
BkmI6eaRTMbZ9d+dPS2KErS5fDwB4Hjr6Av1zLqdLOXIkLGa9bQV+CrEfGVPyXlyKDytvHvOHgBf
dPBx810oQCDIkwUuNdM+b+CjZDkcQIdqRqIhFbT7wKkGg8x445A9Utoyj0ihwaZ2f/W8phUa0mnA
4zD8xdh2UJBsfPBE571lWGDWQS1VEtGiI7JuJ8pLTVqoYQwjwlLOYlu2l4yWQEAUgXI3PBBBIn0t
ijSMxIV5QdLrfttITQF8vlHz4P0Hi7lpGaP/yjhP6CC8N8czqPOyNxJPXv4dQKwzNyPKuut035bI
/i9xluuOQXoO02LtrKnvE/6NxGZhDFpbw9XOJ85oLy/ZbL6dVXKNXfLYspAt24Q6bQXAEQMH94Wu
gLIa2NnidbQn4wvwRu4a6jslmR2aq9OKsu3W1+XLXBKICMfEzGgGzOH/kOX1Cjzol+dXSgWIN110
znPxbPMunamnBQ3zeS5FiJdsZ5I2QRCURtoSKkWOGXMRmwPiKisacYHKcVgYRPQ5VPKHjYEysEvX
d96ChVLDet6UsFQA7WSw+rgh1UoITGp0NdRAJgwuWCSv6Qr+Vsz6QKM6CwyqZqmkWsfyt8VZVsgn
LHH/4sXyEcoh+2WEPfGgLAI4ArYl0nXOXUcyfE+YMiazcrTZDXDDnnEQhmpGdZFVsgyPsW1rRLDs
3fU2XOtojcDPMoIiXTc/uPsuo4tXRUQz09oyn6opS7t1XmIfifta0z3ySO7PsixiR9LPq5x3ChNQ
toJzkVkF5pOSs3+1zL1LeFq8+vSX27+7xcO9fFGCfwVZz1Iy0MdjBl9qxCJma7Ja+gr+SHuBi0Bm
4ObmF1qfMRROC5+laBZXep3HXEXzfGeRhe78wQorYEHAZaFRVHWdVYSh+NDusuzoU1BVFuBoTDNz
ahaP9DQek73x9+EoAnAqO0B1whSswK6FrCp90QzXtshc8jBSAjxQfID5sMwDMjNfsYe5emRRGTkR
z7vrxPRn/iTsud/TsxnzkUr4Ayv0Kq2hK8mC1z7ygRUyW2vr9TRFHQCHfhkX6z7GmpgXeydFzUfE
FIPZyQnMb4+MDZptubfNbdA6z111+DoKyxjmR42KaF4ypmvY9V2RkWv9CeuBUkPaEZy/vWgAP6Ni
tXpDTb7Fxkj2uzM37ZBBMDVVVvis+aAqZGM/efZNP2Us2qriKZHP80eatKGI9eWPwgKkkSO60/y6
6X51/sEr43QbnadIrUys4OHckEYH0x24HcaS02OnJufS9Qro5Rz8IGEh1Z70LwUvQUFZw3T6rEt9
WCyAvEYR6tL2Lg2iK94lMgFYJNkeOxweaC5M05jC2sOteUy+H83Qwsnz9gnkbxtk64NuhxLRJ23P
TyeUZVqzQDYdvFw8YxWU2X7iAfOQrhW7kCQqi73pH+wADgX+knuVbSxG3hxvMGzJN4eRH5QQJ6wR
hConCNE61ASd5NNlhtlphvnDAwQnjkqJNHG76i8vYRVzborNdyG49tyD0PiigJNH79TGe90Qfats
mMNQLTiB0lEqbOGg+roklwX4UguXUDPGgB4Tfm65zAWe3aNeFF0KImX+ioWQFbIItFGz6aNUt7W/
u/w+WJAYbE98lMNSEqhhgxERrr5on9Fds7Bm0UqxK2RPe69bCQ2t5OWpk+wyZ4ZJzWS4lbpOzp80
fiYnfqPh0HHFo+qoNiP7Lj18kqO7WBhOGpKtbjA4j4kYAln6hXLJ3UsoPNfQGVoQrIjkXPQUdzJ8
0sMQ8JXqRtaH1MQaDbc6hl3wlX3MyHNeH/I/+lDcvL7f1EqScYUk/r6MBZYNLfk0k1MTjEAxlkxT
3uGFxBZykrlpMleOejZVgUiKigFWAu3ZQdG/BD4cCW0BpQXzkCOD72ZR+YqaAs9IGNHlUB/KtPe8
DPFj/TnQZFylSk49dTPWmaehx/KqS0gkBXLWIIebcUa6ioFgpArmAh70e4xON/FGe4m9kgHRpHoZ
lneG5PFz5iA/Knr2j41cv1afs1CDDMTXHMJku05OV4qo1DII7s/GGTpxHaQxviFcjn1XgZRHFWjK
3/YhHYUy/ytgW+g7FxbjhS7QcgnU04UtCB3cjLJeQYTlqgbwLSPtO1MthOm2u6O0rRCUnLZT8fQf
5wua5MesRAaNF1guOYHOcX/AfjsWUa0FCLouvPQA8EIvTcqTxK3SIDAOHFmpyXwCgESjSnOckVRC
KCliVJhSggfQrv1PC2TprS0gCr+ujS1yDDK2pHulLgTxMBmkcCYQR3ts5UJ15rWYfqQ8ZSmkc1vg
z4VnS1dyoKo2rchGADf745aC0hNH7TiOlJo258Nr65vIVnkCxi4oK6HTbcrRxJeiMY6bE6kCWbZu
0+2S+FiLGt57epGl7iYpktBFiWKzGtb1RbOCuVSO0YI99yAXb7xNzXgbOsLm8yn52DXYW0UOfE2G
ovhuaK3ETVZOzgmuMhBPtmbyp5uADZ+c/FqxAdv39VbD1QCtqPMxFUtBh/aioBQQx8G3WwnZCWw0
EJ3+KwkRssEaSZ0MrWxqQ7Nt2w/5LgQT+gsb0zqOVRUYFcsqmLVFRrfWWEVhjdMgZ4e5xMpQgoQQ
9TeguhXcGfxdOb4DGNYfQv//5WLyWdTmxhpj62XMCz/oUH4kh1sXJsg3+OWciG5dNrMDRamT+gyg
h5SVdgdA+/Y32IMy8BPpqrztD5NZ2bvUmofg93R5HlqPxu1LJS/CZHX1Orh1bnGcvnpgl91Rpmqe
/eh5oopA79mO+r06SYX5LKPAxSdLApiDBC/xaZrzN3MNsX7DF0JpqW8KqHk4JC7vWiEcDrwZVFP8
x3boNxz9SsjZNXIqRnhDE6IPU4RXHgd1+2PEceUw5CFA9UIbojgIcmJsgsF7ZeZQv0s43uYcGu7+
NnDFxLwNOwIkfcYAro/iWzIvMZrL0cORXasHtCkcER9KgMIv1vaAnRseQU+LuPJA3kVeHwtcmfr0
sdo8gnAetLoWu8DyllTqs9MFUfVywYX5uZhG0sHCMEeV+/9FK8J61qhu2nRuojDqgFfFxcmyTKuw
lyqnGEloAhyr3J7PO8gxj//jzPxhxUdTm4LG9KnJgl4JTqeYzPZREWRfcbAXr55oHUri3Xm32ZJ5
5xaA7R4MDRJAm4aKQatI9/P3vuzqw97MUwmuFisEzJOnl8W/M743yWWedK0O1mOsNlG2VOXAZC/q
ereQa7z5FbGT9sPZjQYleRNT/yoRxy7FjUylBq4NjjtQmwwPnKwlTBrGetfG1YCNEQcN/RcPoTFL
RZ7O0/WB/p6Nbgnzp6jj6XU7YHXWC94/f1H4EiNoG1oT1ZBKwoV3FielXAGSoIRYlRqFizdrtu/Z
ha5ZV/In5INd6JrkPzGrlc7BAUJvDnl63byOQ93iOW3GNKFA0Xgb0uTm4UtUc+J8QWgB9146MEF0
G7POBxrZqsE5Im3PJlyVpldWjNflvbhJUG1z3k//eIh7PoiFiZ1hCvzrRZxRsyhS1A/Muxz7IecE
RV067HTUamVD7N/74BKcay9fjObesGl+e+hAOsQ8EbYwghn4iWt7dmaFiZXQpykkCUAPxsxEGd5e
9Il3v84mH2epM2YOS3ww3bXlN3tZcwGztShi+8lrxrrcH+y5CZiQJlEp3V3YpYMcVFkJvbVAxpim
J0D7eyA32fBPPhzssE3vCeGgZ9WDXkdsMT9LXvxSPKQirMmNiSkApFUN19SyBj+jia35VqT9SjKb
+WWpcWoUfJrJjOdQ+nVWY8+XOj/FJw+4SKo+XB5iki3dXMDDVDHKKu7Yu0U3NrjMF9NhxFxgmxRV
KCaGnPS5H3DtIaAEAzcinp3DVevMAqvXIlQ8SGGTmmDRko9DnUVwwQTlIQyEUpRvd+E/I26p91z4
1CuAD/C/dl3qqr/2L2pdFauaNvVQZNtR0xn/9yC3PrSsvmJyxS1ViPP8rfO9jd2G+6uxj3+wvqng
itPNKXYsH/NATBwpKI1dVl+MjBwRvSn5p6lGHXQYF22pFF5dbcP0gs73sPA2B1Xn7BjGiyzzp/5Z
HTuP5xeOAAZrqW7AxbGEmB7lmWmi2CVaCsBrCiF9XstJEYing1Se5La77ijHtr0/b/CTBn9pFivy
dFEiX3a1uHT1cd7+PkT4cRCM4gLXcAR5c65EwTBq3ewAlhZp3zQQ/CfRJiMiSRWlGt0A46odPFnh
cgPWjbBwCqHQ/HnblMlrTNmWxBUDGhSnK7eHGfHMOuJmk6gPAeQjofB2puutjSb3EJDcqd8MfKl/
pMtveB8sc7EikjG9SowF7w08/b53D9RLnV/V7bbMg51KRavOTj/LErxBnoPBBoI0F0wWmrn0dNzZ
dTZT5KVf+4rv2JRqYzYEHOZSxUFjV7YPHbqu7DpJIj7eXj5a9VJE+p2AZvd2a6TluY8YtVJaMRiV
O28tn+r/4qlsp0wNcjoCfyOg2vNs/WTGPmAh5M3ZfNVnpBSKgkSiiuwrAjEWjEPmal3Sj5/LkbEx
QbRxKq7cGbp4FOyp+qdyMvczIrSxznW/0VcsGtC68oXXfBF8RDtcCMkKtBQAQqay27cHaqX6V7zK
+Ima3MIt9HCm4br8OnPHYvsrVGCqmaZk7/J0csKZaMVfbUKYkEVlotnOirDd/LJPBnH6KY9KrpxT
z3t0BwcjtqQFBnW/THFaZ4LHRToulpeymqWQjwtfkfprOAxC6afnLu/OuxET1IVY6aRjp0UFvWTC
MXlU4iB0exeOuX+xm+zQkQv4n6Mers0p3JrZ5IvtES7BRolz0Mq3N+MUQP5XqQHE8fTqQWeSeUOh
LwohvkMCI7HvwiBKDTDzEgX2YADkREO5n6Jexegve7hZUZJsay7zpKa3daBFoF0nDAqUBkL9TvKx
79QmfLgB57kJq5NSUJ5MkY1hbZNiOxPOiPUx4XNvCCLt0DW4smhDCFUs5eDDfzpND/lBK81RxCao
Q6H9oUhGuMplv4ieF01lijSTLccxX1zuBVhN8a71e+QXqg/NUb6D09CCUZ9VZkCeBg9M5POKARQH
JcWqjDkJzpC1TEedLyptb/ZCMnBB5IOSdJstjUTSD6QTOS+UeXk9R5so80ITqzarhQ/tD2AMtkGQ
QmZPLnA8hXeHbakcrTm6h1BQxhwqf7ek3Kt7mC2fEp2Bt7+y02fu+tjztJuHjOS1d+gxNOG/6Tls
lSadAs+y/HbPGNjZgGd049wS0lfAPWZgzE1fwrbPFgblziMHZIBf7At1xlJ+BX0+fSZC5cpPW520
o/Ceg6XIw/XYJxI/O3pBy7uLtE02qV1bmSUCUJQzKPJ3J2leroIkdcazzqlPbxc9HSjdiumTanb7
ecFgNA8JwfJjc00UyLcMp83kJHGGz0rfTHXctTR+jdC+0g55XWmpDiAdOQYS9TicsU67PtGw4Vq6
j0FLOvLr17/kfLjxitZJOIOptMeYDswHe/5hWXSN+niRQOelHkgpK0tbqeHQ6vXDEtwCGCu2pXzj
Sg/o2upVgX8WfumUbbWJwSyXFOrQky5ceUnWDtulNfeZFtZfQamPrBPw5N0NH5CSjk1JqeXd2Ttc
dIUy24rhdnXvi2TxI500krPbFPXNZUQ0jcrC3gZRZmo8KiNpN727QBWtZudkjj9xzv5KJN9+oYvi
9bATGqD0DElSQ2BRSQ5bbZuUyRBKj7sx0cN5TC2thhhsW47PlgaLpsyrFhZIoVxQLC1ddouLPWN2
la+Bozq1sRJLUCaW1qJol6qeGDPS8DD3Y5vjC9hNaRsAgNlRc/zD31UAwKF7X0lijCbbH3MDK/Rh
9mXlklEf4t4qnP9FkGWZogYhsLu7jkWT26Yo2Hg5m+rUp5seMsU4l+0gknTd8aQV1QSC90QXddyq
ZBmIdVLupZiuOC8KgV3jsrC3CHfZDiOhPY89GrRnetSZBgxNHDFT3y5qAN8HnZEpKAWdJ6o1Fj4s
egVxzzZ5t+hgrePDaUZBwuXSE1XZ3ruSRG+l+vnm6AqrbzE8LAM/0yNo/W6A+NT8cU1nH/wp/2vP
yECDY99fCKyf2XK9+TbDuO4EODvWYy6at3daHE8abxeigMuqCDBgMbptFz8V8Yz2M7zMyOs6MsnO
EesliCTVYmhf/mWC3xbIV+iaXqp5PTqDog6A6FXLA/tX8NOT5ngh8vrF1x+7FD7seGd7wHPQXxqm
baOo1Ed76wAfeaRInxhAXmRV4+ZHIjvLBorcuPgS6sTvm68zFURoXoUiw8KjICOQCJt3Zw+UPML7
IQzTBJIr/RX3zmIwQbvbV/N2mfRa4w1BWyv5tKYShjswoGYyChmhzVdVOYDtc+yY3FclWbyrfG5k
XTNssoc+2FsKZWTp2OEFW1WDBRTQHLqraYPOtvRpVPXertnkVeiIFKz9MZ0tgXowp+33LVkEA2zp
dm2ntQ+E+mcBX1Ikqndn/qfO0xKAyiePdnHN22McNzKi/eInuo76ISu9Cb5Q9IHMjW+0mGRvTLYu
uireAybdwkjFSyzHuQXvYJjSulMyR50MZLmmjrRUtUssugY+mUrxXWllCB77g3nBOmztkAoth/r/
IHLdQ1ooQrR6+AsWLrGbt0HoJLf9k8Oyn26+X6d4jbglHIanhFWWnSX113h9k1vBkvnQk9nnyI2P
pj4GsEEFbtjtql92gnmyer7vlkLBPX39uX2jTsGs1p5Orc1A/Rgs3PlXh9C1Gvhkj1BvPETf/6nV
sgjGb9GyEah0ezIOamG4b8BbtKMdG0dufS9OALxQ5E+R64g+a2+mD0dW79cRyvdpjdXjs5kohfjD
Yb0WxLlhgopOKM5FFzb1PqzADbWLyCghNccOyQsfypqPjx9fxb9PcLLrUkzY9r+C+ssQxGc5wzdt
pIjFYcESkY3CvgJaUvzFaCgqZBlaWpcCWmNz0DA6j8OSk8SXS75LPP/RIxUERADlT5XDQAXDtYDd
oyXUhI/bNMF/Jda1axL95NyLwuCBm9nA4Lu+zDB50k8mvLKBZY4qQDpsAiCwsxnZjO4Tfd0fcnfc
/trn/tpxhMNMfkS1hmDIyqfQvUIbT13+Lkt7yuxIuz+PaAXa1ec0WewWZuNPvjdQ+zpAFfBTkDiM
5AEbYG8mRWXkfFe3OshzSrJ4h1Sh6GVPNqevbjxPBlltnTE3KasAKVRaPNADpUZxUyLtzHXAtCE1
dO9DFj6H7f5RCp7qV8I/BH30URCIfaYJ1rzRkAshYml4fPhjZlwZAhcDAfYXuUDhw4opX1tXPi/E
Qocejgj1N18bfsUibOjd0VUXscAT5XYtAoiEQUye1Si+C9AKLL3rl6LWR4e4ZK09XwvoOMnVqdbV
f386zcF5gKjPJ8npLmEAvXZfS3AR7xBkJ9cwX4djxqpwg3zILAdRnscTW/51x4cfh+80DxdOencZ
ZM3zmHzNnjlS8w+u0RBxsp/j3et6dwW/W7WtWvkcR2Q4SGagXjpherwTpecg7+4uleEfu7Ki3y59
CEpqhjiODrgUq+kr2D6mco/RLrf39UNELqApuciiq458PdhKi8lg54gpKEMuX5kfy7V5wALOwdl1
L/2/l720Yo1E5byaqUa1FzqTP0jVyg/pvKVe2TwdFmsRol96sOsAAk39Q30meOFE/bwR59A9AGp8
6kJz7VWbDhxrpZle091HbT1dF79fXNmiyrcBz/kIWubYZJP7o7I1L3eV+JHlEOdEGXW5SHeC+bvC
rxWuBafl2uP4SUstxi3xJyE1OJUGDNP8PxWNuvTIbJPQAqIiESrPz+V/kxubLyuwm1UIYg26xc2d
JsG+4UjdlofF+iUZSLTYwZISuC8kQ238dTKMGw6ZzfnYooPGRa14zinl0xJH9P3fMptqYetlKijY
O+PeqXa1D90I01TlOzcKQUYU1JdnIsSs3nCvJ7YHrbTu/aKzu0PWOb/5A8OOOYnoNkxT0EE7NsUx
73ReEwyRj8RGrNF71zifs85P3yg83Ip3aV8h4oUI9/3BmLUo66hZP2DePmtcu8+rTLMmP49LhLN+
9yb4UPGYdTbgwAnb4XX8a/g4q9hTfx8H1CEG8CIox/bZeMQnwONdoZsiDFNiGwsZTEIKok7Ztz8e
GKZse1RTCEQHV7A1rO4zgKm3ckkE7p/PdEiL6oYnmOOjQ25reoJBHnE7WuCbkmDEdS744596ikrV
KwN704bMtrBv/UWy8T7fUA6cwNIiYmnqtHjUHZpt/UJBd8mf1eDlZ7X17I6CgdnMUP6CDYt64eB7
1zutycjk26mM3CaII+ytDaKrI0vOVfCj3YOMVmij0KbrI7SdwpnbIB7+HlaBjNTJxciQkfNUvX4J
lRLIatipag5D1VVR4xJE6Ua7fHkmC1UUxEhoh4B2a9hXLs56Hh3S2pvh3eRdumDTGX+AytR9UEKZ
Zw1wDquIkNfEOsoHiA70uDP7xw5fyE1MSigsd6SbP34nyojc0dv2mjK8YJFlkv1z1vym9Qz14pkb
UxBw9IyDP7pFudMnX0QsPian9NffgRrNWCTsrIW+iuuse89ZiCEWQe03D0YEyM/w/LWGGIzxKA4f
2o5FnS8irF9Iu/VXMC8R3I4YBhI7chFd/+PgfCJkw4BbHb0bszQjtL2wWPGYWMJkyC89IAgfAb3R
b3HrxHghUIkeaP6l74cyborv3UptolOLnm16N5bQfIv2j/1hSwQXLQwuAw/tek/HbM0KgRI3BOuo
95AzoG1168yBCInXUD+WFivvs59X4pRgbr2JKZzAmjDe63Mp4ItMgejK49z6lTzYKsFW8vUamUXz
jQjJ++6bvSIAPj9WuYBn47zdt0QX6jnVs9r/miBa9JU7yPWAL+nq8gIzYcOy1r3pA6lmN7TiZO3Q
gsml4Jb//+L1zSeey0Ilz8xWQw5mDhBdGnUj9dqoQoLBZ38Jeb2d12kvs7HLYsFUZWOUUr8w2Ah/
AahMNJJYNAkiBHjGJuiQ1c6upM6sjlOD+i3xSQhcGyUA+ydTv6RwiuifdT7NDXoy0IlV8U8yBeos
n4TJk7I7pMMxALXRouuVm+2jf6eTjgCtx7Cl5rknulQYcaPB4V1t1RN6L0Xtf1TXKDm09Cqb8FVz
jQexLGuwJJOBHGF5t1CtfJFwcnVgV2Lu7/wYJz8IMz86T1VkcZSrDPtOqwM8ILp6rGBuloDPI5IG
aQ8a94UxR3XoCVul8629dd4vV9Vn5iqkxGu6yRZlhwGG3tpIfisOBdnu2xwJLEV1Z+xOgTsSRot5
/q9p3QOnZFzeo1Ma2ALbGNniebWCN0PQ82qIKH13oEecZOyqg5L/NOtvyqjkPwemEJnO5srLuZ7M
4JyXfpXKKS6iBPpgs7dKFzkWePeNMLy5DQjkaua9k4usIU6qswKrROqBeJg+Jd5Zi51NBBNNY3y+
+TyJopK2M49gK5LxyzeKAWoKJmmQnmi+86SvR5kIM9FCd24HyC/2gW13NVvxa4AbNb430DHErOYJ
V/0d6yqKs3tC+1ggkZYq4tbPupPEzURy/56DtLA/jneEHsNyeBF/LbKsroK4CM4utC0ySUcNmHik
Q8j7NNkfNgYsBmk5s201FLxrMbFCV6XOfj9tB8bgTNBuGjRoWpp7V+SVZ0lu/ztbP8/EaCUCmxXA
afDWOpOcU7ZX8+BuCIFx4OV7OHuYP7H7/x1k0r3DLkdqJqkL7vxbD2R02vBpHOsswsoOc8YgmTfo
OD/ZkCJOcXDhBEXyGUQuc473A9WGoqDl3+PK/Z9uFeHE4MuS6dNolRSW7c7LmMdEnZKHj4b5d968
mP4fiyYo4bue+kALEPg9UHdOpntvagq6ziL7ij8DVdovOIqZjm+m/uz8TWCLp5GLJYXgRFj6PZ1K
2wjHnSXZD6H502d+Arcx3MKaAviC9HO8yziI25jHnKr6AH61SVTnv3SrCZlEfCTbKDhPSkXGyH+y
r/aoBJzIQmO3YCbIaTemZKqb7TOK3Z9QreeDYs1mN6bvXbhy0ox3SSDPnEq+iCvIPMZFu3gHLa2P
/TdfllR1u8hgxRp+P8heE47Cq2ttlVAtyrC0CZfs95VJjl0U0bQrsBCouWTo9qDV8FByX1dpRdZH
uiLkYZadjkqxnlxlLEqaiZde6GP4TKwYBPqwHF4A5nin5qe+fsUG/+MXJFpNHP2ARuhSiGPPUM+1
18LRig8KqsofLwEcO/p6ceoLRea05KrHAxiG3d5/6CulxVXsxktMR4Mm1gr9GjvvROwHTXc/cvno
gs6txpbCNnBXlDbwNr1TEpKEiypiJRrIV44kSZkdBPwWXOz1kbNdL3tRICeJB1Ic6oHWDmN2XpmD
9kt6kcD5BkHJpOlcwPOzegTGjiWh/g5PfMKfWHU2dpBMXsAKW2lXbqNPmbS5GXEd9iXdBG3n/qn4
7uewgvqG4z20HtOqgGBXl6Zibp7/VV6gUhYalQTBB0CfA2LHAvUArJcQtnBSCwbiKuwjnFHoeewQ
zNwBI7lcDOijQub4Nf4deaqnDuTemdn2FyXR2dv8BR67sLJIezei01xUFqQKX+tcg/Wj5tElsAaM
kWC2XW+aNSWr3h/gtq9poCNeAWzUhhWQE4hOdmTidRiuuw1H+ggHi6vv/4iBvpqYYUxIVfRcAcZT
eM3xhHH55PgA88bCfPAzxwc5BEpgCf0qqivDqWkmeuG4tc2AgYhfBP6vsBY35HLIzeQMxO61YYRc
7nwE+Y13cyNz8mWj2bQl7ZnXpPuAc8jydTEjQVfrCDoCmtZLjocuCy8IABAaNsgml2k6HsDI1dgY
Baq1IHwHhg8vKBub0vNeeO5uFmqhfKxv3OAV9lA3XsrECtm3ZrFIPne2fNJyaBzm6ghJFMibA04T
tlhJTdPugVziwkIPKYb5g/MDq9/YSvNxQYJ9UASe953emsRnZcoq9EiOkejkZM83OKh3rtxjbl4G
Nn6M7dxUmNxaekZRwYCwqrhB+PZV1qyuVb9ZZ6zrhH5sMTf+Z/1Y+H6vZ1ybKkgLTPMCjyankyY5
87g22uo0yRHv5jYXDTwlRMkJtLWXuUrLbl/f/sqjnCZpgtZrPmCiglXfwlVgeT1hMcSRYzt3yqg/
dfw+V1T1CjUHrFAZk4du2J1YT9N+WpvlLIw0fkHEX3joY84EmJJM6e5dy4SkmVJeNI+02o7uHvuu
Io9tDoUo9tDDZ/R9lDFNePy2Q1LsORuXEdRoCkLFZMh+AVFy2t6JqgGE/kknvLgxbBlNI1zKF2Hr
jreM8glvmT4RiQEtcGTf+FLKBoanasc1v8apzOAJe0pgrWcX7ZavuerevNbOpt3yHEVxURTkcTiu
TL4Wbsze4Sp9fPrW7o9hIrjdZGaivJGxJUOiBAGSlBamB7doSXr4yOLwp8X6y55z3YIczhbSO9fF
rimRt6vczDBfk5E04LVmiIphQ+zFlFpCy+FFLBbGHIdgJaMZM6VSMPVPzvVhiK/bwduwNEgn+W7G
1y90IYVpiMMx4w3VbOiWGtuWXbcInqDqz2vbttsN5jvqNftcNrN3m3K3i21LEPA6X/TuArBPYVrM
tUWDtYrOjc5z3Hvo7v1EsJEZ7Os9fXrhGwR5Tx9yLO5Ppq6V/qOuGe4dqsuZukepp4u31GoUQy4O
Qzk6jg590U8b0S7h9FIlwCM837tBmJLL6EBey3Tpl3enpNlVdUVq3z11p/eKExeu7gpvQHiDd+vH
nW104HafU1Ai/UFDtr/XGPh+AMUq5s/8jMskzWF64R3IG4zj1/GgZT02VNo5YH8p7h3NJNS8aWVV
a37dtjPmSF8bREpcwjcLDMmWo6weNx9mPihDUDoB7FLmqolk9fZVnDW6CkPqtAtZ+5Z8nNl0XRwJ
IwGMQh47iCf9ho75I8/p0Gc8cX+rgxo21txMWvqVKFghk98rU4jkRspbX8eAzuGzs4+JWJyBtBB9
I2n6Wp3nKLXW42IVlIoRoz+FEPQiB6eIR8+3x9z5129q1Rdb4D4gDcx5Bq/uLJCzoA6XHaED+MXb
2pTO4DAWmn66AqAPm60/CXPDs7jjTfe8KEA+yjq95Ao7iKR8+cAN4SIKGq4krVrBlAqt9mwO0jzb
gL1mh+kMAE1oZWGr90mZ2j9LzT63XfA3cj14dFoFFDUOM2Ag+0yM1d4pPru3T3/IhO7wqjVRk0FR
CHUuRpXp4Y63KX9u8rj3XFjK8wV5FuU2fhnb3BvbsCz8r0NJQ9toy8KOiLOOMV5IP0xfkgM1cKz0
NJX3z7sZeb0mKNThEMN/EG0LgWZXzjzCIV8BhZP9Y18kD9zZSWRy/Z2abWa7qr+ZB1C1ROeLEKYb
pboVAi/FjHpsreznQ2klbyVHDBc5/Wmzdi92sXdyxRa3YrlKR594O4+aQOp/MoMVjp4uRcGVqv+5
xRYRX+TzSRKgICm22Q2LJWPKv4ahfjiCCqmzjuorMlxaZA68ofP0Y6hDYl3GI7H+sYKQjE+gJ/Vv
hOM6BZvPtjjCjdYOBNgh8rpp60LTY58zd5IR9BIPv5A0UuExtN1rG25uwN0yK1JqZpcumsxAImoJ
rArbrhN1wwItw6XCaXBX/mOUl87PaaHnmiwHnZ3Ydk2jZfiX4rhdoDMlRtrEYG9zCRe+kqK4wpnq
6GDqwlNs2wheuAykgYoXezI2jYVn8TdPtJ2pkIBRkawQAVd1h5Hy/5lHWGTy2SBs/IaJvuM8SVcW
RgZ+ibC+Vs0qfeoASaAB+UlpNx11XAzLzKwcisdK8gj/hlMDLCwA/17pQfrD/QmNjn/esNmwyk64
QxRp/2g/5gTtyxXXbHg6tPRM9VbGMurueoJ9/+S9Eu2oi2juzOalA6khZ3Eqdz4+wV97RnvqTv/8
4/FfR/gAwxXvzAOEMMUgMgRuycpHC1fVDsnZIQQJciZ2CWzRgvQJ1CMxTjbKKx8B1eQkHMqdo2KG
mIw0QJNRjChmU8AVkd8Gv8N9ygZU3XnuES1BG424k8h7s9F7F6gQtDjYteMqzsvRV90h4k9N76tN
qeyu/9Fhdy7wkN1Dd2gLwL803CVlx/bRD5mbaCYqDoW1ezV1q9SWpov6+94X1oNZhh3hs/4u9045
+7CrKq78FYJbPyH6K1wkj95r1v4SzNM6gfCcL5eqLwPfksoZvPMzZ5shfmAqj7bbAh4kVXrtKe5h
92XR4iJOoikhUV+3qZUNKqtl0PLB1plGz6XHUiLq/nAYOxTDXRi1DCCirilEKAjiUnRe78nfHM/m
FgQwQ6dwrSIj6PHlBZFWnp5qYhDDpgm1HKCq3wTwlKZcE5hC5lpwptAE7GYzB8sAvjwS+/1/v9P6
r751pzpFiTPauAaUn1m7Rd7+4SmGoriXO36jG0YdtieSrJuRFWzMqwH5t02yZ4dc4y2gAHi5HfiC
6HHbcQJrvqP60YfpNZ/TAlFU2jwirbPbR0CIbpAXMN9C5o+ENjHJHYEKl2+X0zfNNTIGVc520aMK
lE9gUU4fH6cZJYnpnnF+M1aRn5ApUbj7KmJgdh/01vKVbxMu1xRJb2XeyIsPpqL8jGxOl1GqfV+O
axkRzpNkL+ud0stJffGrgt7GxUCwLmUrlP8Wzu1BKeQNDFq5Tmj1yy/5WK5Un4Qyg+atwqgJbF4c
iIHIVYi7vmnstcHxaFmuv51o8TfbB1VplbMF93JvkQ9pQUrPpQykTrzJhfpSEnMoWHBjRlS/tgKw
CeJPg/0BmLwek2lZ23pkJ/Xjg0rVZV90iSXc91Spy5JGZXiZy9/+mCSM23lCJgRQ4aSfjzgu6RUs
x+ALBZDMiSwzZer+LOMNSebx1OzFwTCekuxY6G+bKlhOUhjt6XgAvviZX9PatWrfjwwpv+R9C1Mg
9DMxsZdHrto9644KldDKnxVKMXxyprSIYXa5irX6zaoDByXEJM62eElIp3lz2pIVxG7ij9Odi6gt
JAHCWUpYwB2YQ3/m7a3AWjIbu8UTmshxTNCUSc9dWZ9opdO0abJ4PmMwIgBW3TAFoAZhbG3KLcu5
yGORfyRFMU3URbdfIzTQRAWLYfTJZHBRv/8YlNR87iS+dBXauhl1swvSEK0hD/KBqH2e0zr1q+eS
h2WvxzyEBXr+0IfePY2kjcpoWC1o6k9wFUuuNEJyeWN+zrum/jIqVJ+FaDD2dhzwfrKJxjIBJLfQ
nYwofqYLXxNILUaUwjcjSNlMIQ7ZtgXnuN3td+twsBq/GFUXbLWvxBj4g28XyqTPB+0g22cV2/Gw
wU2Ooe9iu/KR/UAu0fzQjAYbpPL5mX+Dj7NtCjryp2AXmSbiBWe5CmHjNMjEYaRuqc8zdk5sim3P
EHd4sr31DW1nFkUTBkRb3scM2bgWmr5PP4RxBx5y3hrChuWDhlU4GL+9b19sgO6SPKTRaPSq61R5
fu6fd9VbW576w3/77npy08oDfOf2QYoaHFmWjc5QDSBDf/SrSWWNUIEoNYO+yQGCFZY4r/AvfJ8q
vUkTI0V/nJlRa4eovtAmMdY7HbM5eHrFe7zqpqmtS1it3IEfH3UgJ6FiIm1vHmKxD6t2nGzsSX0r
+puCHbeih8Q3X0tmA7razB2PSjRzzZicLTzfo/1o5HuvukGya6Ysc8RySMpKI6PTfAJRnH+57nu4
VBGuDmvhA1eqXm+B1l6bejrxrq7XwaTRUsxb9ogWNgPY4ZBUQ7bb2QhB47p4HzO2dX/5tbhP8Dzi
u5wLgwZMfOka4REfsvfydV2DFTlvcDupA0L74PSqkBeM/yvbjbfbTjaZzM77Vq/UBIW7J0oR3A5b
63tjZQjO85TAwnI/MyoBAxufzsJ+tvhNNuTmbMQfDuLxkq3ZbDb47Gs1YJCIN6FH2wmRehX9YUZg
WmN376xQRzpINuz4FV6HxMEGxLfBuWh0U+ZYNPMsQRoMWOsodF19Uf+KgiQH8g0jcZd2ijNUnPv8
JmJNtuVkAm94Ey28GrhhbI5jjDdVb5iCmpU1VKB3ssLDxxwx0u1Nw7t6guPgGI4NIEKMHqBp7x0+
h/CtPRASo2RoCdW8aHZzf+TktGgm27MvjDIEBAJitnfDu3JvNs/7bOqkAhgUPs23tdR0UW6VIeEb
Zeea7plsrR599iL6c/ENWoHPCyoW3wC23i3GYt6IU/n7pAfqPeaMNoUYhnHnyXJRvChwI7IybbVs
FPxV0cnhXUKdXklUPEn0b7D/itHVljZEzZpTtf5P5+AqtiOWoGr5B5a2ZHjPWl17kmtC4uFPsIa8
vyH4UeZcM0kLnRWyle12cgmLXgzb3NzWJ9BMhAMgX6KD63TZ8Np31RXvh1D1cUtlULB/mQvNd31f
jy6RwXni+cFMXTZoxB94A7aj/PabNzSwyIYQTqxmxdQKfqi9DZi3qiYXX6+vDOvF7e2Te510pyo7
ynq8TIfgqmfokH//Q0mUdZRC5d6AMpRep0WNcwYa6kDvAnpp1pkxxkv+spXMnwVUMTXc1yV7AywX
KH5bHtqTBhFbGWQOXlcfGGTnfGf+xdfsK6OuEZMqXvWJ4Af7W/v2LCFwRSzD/jBeNLJH9kDK9xw5
OiyU2tLfUr6/drKMEkVE05U4CtAtEnYDPcPOqd8Az0JlFZjYiPH8z674iBF1vEh/YR2A0dlVI+o0
rfIDCClBd8MEZPFH6Y4nvEnbl79SrkkkHG4s7AZmHdswBcNF1RoMRxRPQHFo4mPTei93ZTL/Fn+i
xDJrShVd36Fj7bqmvLqkjl1d2IZzkHwEtGQUjgclWH5jWXydrQD2oA0Pq7HnD5TsDZiUSjdQJT01
OEjnspnuG7nje1b28dE8EpfU680GWaSmAnHa0bya81nYD7TWrIcJ4ra7oNqWBkW+ndePh/lC+Ufv
AX/uPSUAGYVxFpVXBpdkP/cbCvIlDRfIuYbpRKYhGGwwyWU0AcUAug8nQL3GeIugbaV1PBJxKuAg
kI3cxWMvqq0PfMbJIlE3PBUn8cSvCceXjwtqG53wb5ucEvyPKDfDjSRmX4MmZc1bRXkbkiRmDlbZ
k4RPDH+q/l28sAJ04HmoejyG5HGFAQd1SqKnwku/wwKMYoeuAPQsZouerHynV1szCg0P+7eqxjAw
D8e2Sak/msa9lz7C2Usne73ZqcFqT1Xh/zlzpHiQL1cCb9NnJMJpyn6P7pG3N6Jp7CrZkEJ509QJ
nnNBQOyk8TVjvkxDTDBxyDB2XmfQZeAUwnY3CGx1BNRDXlGpqzG89/9O888n4llbLhKt7U4Dy3o7
cP1ymSS9s820iqMkbVq9mXXJthItcvC4qqVx1BhLncxn2KP875hVFr2SdUmow7N+dN5Ndlo8Yong
jaHGc51gURCNmOpMn43lzxgdeCNUZQ2vmlc6LoskHv2EE1zfpGoVdlgioMR0zFepAHEYufTLuKgn
UeGqVM8fLogl1ITgC70mF2JijuwjawmeDe5Aun35N8BWxxrzBVOYVm5rXYOWUPrgQ3n54qfas9IY
WqTkS1mVU60+kM0/eDigOfLWK7ODOgiuJWkIFGsBVzZUuflgB87gQ7+6Dxhs4SZUqu52HJjFYyaB
tabcjImmLQheSU0QvCvRxVSP0JqoIEtJ/MsqAaKxq4tB19asmAaPco+e9PlZMvX93G/luYkjWAlg
Yzu7N9OVww4a78QH2S4ekLHaNBDNgBLzeFbzaTw8+bdfQYTX3o02MJXtAHI4Y6VQ2OSZ5jvZt6Wi
xYd/53uuvv2Bo4H2h7Pylm1yJdY5aTHmIzSXu2VHMPw6BH5XHBdTVeBDEKzOoWYn7hxKHBm5FRee
xq6ZNDzCco58ht8VaW3eOsC40H9ZK+2U72hE9X7jS2xnyaDCWjtdRyqlIQpY7dJJcbN+LKgHMeZl
E0SSUHfDITraGFgudY7TmbVcvdbwB2JAr5iS0KIvtiZDsH+32Iu9vYvLV13UaIysv2Tx0EHEgeXg
QLVP7FrHEMxUgfWjBdOnYOsNnGk7wqN03q1+GXuO98lEfnVCEojGHfHunXdKw4/ZCV64gOZlLhHu
7sikkoHSprJERMo3BX2xPu3Vy6QmHsBIPfipcrRxs8b7ff5qWL0NW4222N6KHVcePEdJNxAtpJj/
hkRkbKWiSCRPxEA04PG2TQLU2JdEM5fyr55Dqv784A4zsM1+GSOSHyAtInTsN+D6SgfUN6P0WXfs
q1qwVJ7gkhHwSy6urYYl+JxNMc0N0ZKlAoERC1phQxsGj/70WWLkKnOhHNh9PaatksJz+buO2Vr6
Bswe7PNr3q4QrKxbXpSJoFWY7e/mUdCQPS8sJQkUPlpQxzTLZQgjg16kJjQ8NGSjnHsFVQSxTnKv
63s+DiBiaY0GYwveOVgoIsI/lwUTgPnKyTHA4X2USSJcSCL7x8SOCp69d163IxDs7XGsnyXZr8ca
7UyMlgTENUnlkRAWbn7BvvLJXdG0v72JqTONaGqhbjVuTDAB1uz59KwLTMCknhyKVE/Qoh24u3ie
FSMSyUQ5APUw0f2Hbk7bU2on+EMBBQq0f8o3YhW5CnqEp5gySsqTslS5t43br+KWzqmVN4IvJeV+
Ov0Lc2TSSLkH8+dKvswRFHa8XVTNaTKU32waS/Ckolkl7t1dpL1nEs6iMNVEDAtMSsovvFPhv7z/
ZMC9l7NrII8GB8Yd+1uzmzoagwjbWxjSDNdNtX8qBWBAp848+mqZ+175nT8cw489gmo1Kfr3n3C1
pZGzQ2xx5IeMqpi7awfL88+5MlThFYeIumMaZyxTcX9mT0aNQI05bP2mJgGKeo183bzd0wWUNiNx
tayINGYCZ8WCDr89AvrmXETvPEGgnwjIP2LLZkxZhWJE1YQns7EGYEhQso4FeKnM6fs8Y0U66L7g
XsnuLmwlSoCcpWgj4AbXVzwlx8ieOJljC+jdNl20oBzOoD57g87VfYD3vOFOEljr4o1t3Le34ESV
vTUF3t3Ow4cwiS52q/BVg5KPB4ogft77/hKxsjWXfCb54ECOiWE3cbjcxRn4x/XYRGnS/mSo4HK5
8quO6L6thllC6XOpKznBCVGq6hwTxRCJrAgJWuh2nJyVY7krrgR9/zOytgKtnWwfL5lNPhHCzNpR
rOAsvO/sYzB2Lol2EndgKMlbXjfOHbXjiFgOqeY9YJZ9kJuZ99SC7ihkFe1e6uZYnMeDlUf3gXGH
MPrPNhA8tXa5jBx8uIep/fRN121YmLpo29NKLYgW5ctRNeUQjTKKlXibA4XnHyjqcCkXkHqbqkNZ
Y+LXjZdsV59LVMwXxWh6AO/9thiRdFngQrpD+s1usH0qsO82CdDB68aFdKO1kmeL8XmWZYh3Ux+M
gDoOpjSRv+GUlzkF1mKSxKhEmWfUUcILvIoxJn3OSTCQsdRTa8v3kgsB5kF3l+DveZ5ut97prWo+
/Tyw57ss5Hm/Qb+8GfaBeLfMVk9Bth21kvfpwhTN7J/oSotwRVvvnWKFKqONEapi+zWQeOWioN0J
bYt1qFL+GNfh2W5bDuiDN/cMf5tjXvxKFCT3WoEMEbwMmRiTeNGotDavTx4mUemExpFQiTEJkcGi
O21/zD8inh+bZiS/5Qej8QG/M2E7PullAqbyYRQZ0UZcKKokEIyTWwrii7yktf9byRz9DZAvyfc3
24T+E+aopOUXOX481HJM9O6X+mbAcdWkEQ7nW9AULXbm/7ZDxEhzPDvTOtpg8+9Js1pdXcgoeTqK
ltHNq3V10W/BdHt19OTddl+xqU3wgvnljm6wytZ1kqls5EzX6zq2kPSiP9U0mHscw47qwUPfQR0B
XX5D1C0+6ivawoDTC0iPjhxlMyeYuNe4gQmzgNZ8Anr0yEIX/zy2pGbQnA/5CllQIGXWoQ9bYqd2
bMZNW1InLRl8K3N/gzUj8dSzdD0vrSfP2fPGvvMI3zYD+mPfbHhX5MDksEv5afx8bHVEYNrZ+Pqy
+nlaNAPyujyjYRzkO5S90Wi9M/Pyjd4PBRwSq6Nmpu8MPigdLJDkyunGF6Y7QkFj3iE7VjIKvkkT
DaMMqpqMtsaFBW96WdgTFmgnO8605CcgUDlQL/Wtwt8fQ+h/dlz1mme/K97935kgqVSQtd41fS6x
npx7TInrNSaarwpgxq25fTgAUydHNGhOGLGBwQ9krjLBCyOrKQcMIuurxWlZND2LMTvrR8iYQMid
VHmWPXFQSIZgndJzMS8Qa3byrnTou/oIbgRmOx9rGtKcEQ8AFwERnbeIlja8Lw78UdhGIwaJutaB
YtfmOpEXfw956ZjdWAtui3r+jK2+Z3Yd7QBp3erGh3t15gjSRnZ+c8RgMJ4TQUZmaNbCJSoXx7m2
K7upa7DxtJyVPFSrrJXSwPcAOXaVKTEajMiDMPBsA+JJyVYhjaJUoXRYoeq4+Ap3SU1Li+PpW8Sd
oDYM8jC0i7yduJ5yT4ttMCBRxJ3IxeWNq7wqa/AKfVoJ5WGIGIHRto9B3x3TfwwxaERQfBMG0cue
xPewSUGxQQNDCAy765XoHJ18uVlAAVhanZ6dIkMJpm2ogcL9UpwlhVxJiEpCuht7JsYxxm6MAsap
c/01WLdNbFUYL9b8PWAp9bOSt1DoO+hzw0t9Gw+yPSnbq+nNOmMH2fcl3Nmbnc/5GGImru75W6Za
3MTgQAjPpQkGsjbwqBHZ3+6yRUEQgQw0F51wgCRRVptsZXb9TnzKUwQtZW65Upbw40/Xndi95Oli
7Pd+Owit/Hym1yAQQut7XC8VX19YQ0LP5WWem2wMvmAxuuSSRdoagpKFEFwomEG3Tg8TKUuY+WR3
Q6uV3pNOKZ+HcG3xN3P/JSLh5CcCtSEdZIynTPh4Kz6maJzaCwVgRytEluhZzi9RyajigtWk6gNB
AMg9qwIjeD6fLG1T+ZGLMunafBSnNIWrtQ8NyI3Ek1GxQFAfHccQiEpTGx8vk2D9nV6n16OqJ2s6
+D3hO69e0JA0rJiT5gXU6sHVM3M9b7xcnlNoLTB8BiDW0RaKM2rDoj9jCuHR4JDIoxine2dxVQEh
fXxepOu7VD25MNSCa5avEbga6LNmkAWC7Px+6yJQixoH2JCB+raMp9E0WhFkTd+O3Kq0zR4RzR1X
eZKyfhr2YP8R6aD9n+AONcsI1m3Z9d283D4nePd9QSxQvB/O9Xid7f6DexS6SV8/KLYkEjI8cIuR
LM57yJHtwoLeMG7XqA1LjW3s59mATNI7K2PEs5a/RoCZIry19msWe2LK3MYbSMJzJIK3XhQNZNTg
J6cEWFo+CaSmBK8LBhzgmiIwI6A93Uyc12gBQLopf6AYIypZD9RMXkccMi2EPwVq76ABM8VXFaSk
3LR8wUwkmpZlqf98iBv/3eF32+42iRfvMmktcWctDRHcXfvxkfjAFCekWwVTok7nuf4MSJFVyVU2
Wh/Gi5OYhP3FbzgGDd+29quxq4HooMrW/vAu0AvW0sivCwVxWJkvRofECuPYFwWJ8KyYmXo0Bxgf
qsqymjlFpjNplIGHUd36REDniXl1SULwRKOchCYqgn9OZgVdcIDNfsihLprAaDshgcjBVbIrd7h0
RRifv6WdWo8SKgeKAeqr6IHaNWaB1BTGdlwuUHcnAbElmfYa2f+PcLCNTIMdSTtK9KFK/kXkTOu7
1+deSpGmLFpfOO1uw5PM2dgeV+wmGZ8lz7AHHCGobiSZ0uu7wP6wlsi2+DTPZ+8K1rPZvrpM8Ayn
QgTmMRIplYbE0atO7fS6IgxTt6doBQ3KbAgLhHG9X7dnLTOHqLtTBq2A/VREXlzmtdh4v6Tyxs26
sWB2UcCA7o9MzcOovNPm+WLLasSUO+KEIUfH2it8pX3LL02zazfqcGkmkxGaARjWrpHxgP7x0yOp
m0+c9N0LYgd9C5Jm3go65QvxANt11zh3sJbBX5DkQfAvRbM1H94D/6LxJsyndgCUnXt8U0RZiS1B
4nhz90tzmkqStXNjCtc7zImmalcze25uloKYmvzPdRmmu2tsIGbodiraWywHuei8Qkh7oDrSWwQT
YXd8WwIXhak/LuGbLs7vfcJWgh4jUZ/9x9w6HlIt7m4nPFxAjLkTx6SpEjwg9EwaXgSLsxRRx3Fl
v5+YeeoBl7DJFy/aZ+sfnMATAJNET/AO/yDoqDcrE1y97OLuzhsfvg9f0G91yw2J+4SuQHAZeMxJ
pyaWuQz+VlPnX8S75NeNYeLk2Fg/Ne+bs1d/Ufcv/GK9ij5Y+giJZyt8NQhICSJpqEptfe7bdiFC
LzkQk6cqr9C0F6nkVylHAbFO82Rq4WiTUpCM1rx3Hp++KPB09aYs8ubKh/JoWrhj+8hkksP9drSB
0ALLP/4WxcAoL+ifQcIVHitftbmzquFtFCL2shYb2ymclQ9egy9HpWwFGAKXWSq941hME/e1aRAT
LHyDoq6WnacBETbLUH2WalnJB7kOsYkkUq/6/qvgMzOiyLgTpHsUniij5MH5PC6lqZdhgMo+qPgX
WyRb40br3dR3nLRLWM9L1TcD0TbFncihU0eAUSNV3UTfag6o8oSwPwdayPVjUmHT3d4njSHm1Q3Y
ZYYTrz65dP9FZTBwDKfXiRCG69LxoVuKSvYUnBpnZWdAZG6W7okubQYLS7E4WkR9tEtize8fR9x/
Xf3HbWk8ehrMHVyecz6Dh0VtTvcvQhJ38JcG7rJmaXMI/B+u7lO3hq4sfFL+YB7k3GyVIQ8ak49i
DhNsT6foZQIyNjssMnUSH2mlg6VNA3pXFPwlHatiVewE5OjOh7PzruIlAATA8GufquSAezHInP5K
rmd4mQ7l0zeebj1EsHm6N3jHOK1e8lyRWicFNBC+DZHFgQ6e/UgaWtoulm45fgHdBoC2HGGQxG9Y
mrnIcVyPEGhAbkGhArR370BxjxoZohgVrvmwYatVnVfpbm4AOCXA1vAWBPugA0xsg1ru8vj25hWg
VU+GW7IISPAhaxwP0qkefsYVPfZytoOX3pCBcUjQ56sDlkAhZqo5wDRmEoMQ3d5eerZXjjZWZwkm
28MYqKI4NxkqiFZUgPzrJtby7T4N+G70qJ0FynCA9c5xXAyncJd0UOZICCcAB601vUZguCQBdSbl
s9l2ku+CECTy5wPSxBtgVZ7CKLPo0OiUIalGcjUZAJOKuvbIyRxP+wf25hwP5ohmzguaU0mcXEpT
I3IKB4XwG4+/hL1GlPR4tmikYyp4e5T1YcBfDH6ceMTMAk9JfCf0Msd57v8HyZXSHblreJ40wglb
1ppmr3jRLpFXdaTDC5OK5xOctrhci6T2BLSImXQw/O7xkrpRr05Jj0CDPi1QFZ1ryI2r4hHUHI88
XP0NIoAMDke+CcQvJr40uuxz8eCr7QFvqN8XIRg6Q53oZqCckj/UqCufJbs7qxEn2VCMU73otFkB
idWCD2Sh0pUcPRQy/kHno8Ca1O50WtaPw0w2AsEo+F5aCHK+DfFw/wIp2pJtAueQrluj9yVxwzrU
psUie3Imq3xdw9FveADAXn9odcpFf5G/Slph80qtlZQO0DXx3zhIp7lncjQUi2z/6WbniqGWW0rM
kyFkhQNyyK3j+Z7lyB43s25GCzmhl3Me6oNollC20xAPYNTZwQ4+j8VXY3Z7pcjIFfGOTbivT6hO
GaTJP3y9PbAxX+w6pam4pHkYbW7cljQ7EyCFPRkGB35/KG4ujjiwI1xXI8AtJXCMZBBDbPRro0jb
ajrckOTMwS6zZromUH6ZKWS9HA5zS0JoqThQfr7vCfmk/Buy1/vikqi/BGCjb6qgM9w7B0uV59Fp
uGCgEAEkx8WbKVtZCHgy5Pzt5utuu6+ELueeeK30r9XVWp0Zj3OUGGqRbHshFTqlCF9WQDXQT4D8
2U68LtLrv28S0HkBeQPj50ddG8jaHzF7eOoLXtPZNivf5O6bM0yBlAoAsDlzgYuf4seucrcbFvd3
dC5VYiGqYzwzmqDJXt46zFH31OcS/oe/ArP9JOX8kBXQG85i7yuda7Zl4ChcCdqA47vNHCzZ9Ix0
OiGIBC/t7HDmac5LHEcl4guLBlE1cRMofRulfMAZP+a4yHZYseSK50tWQK1pAu0frwYQLkWrR4vt
CbGs49VyoX8YDxF4Mq1nbSTVe4hv5hrSp61DPxmYZA8izsRShdvAr2gytk18BN1E15qDeTw2aa5P
KH5MVrGPlXOTYIbKOlSmb3njsfHUDHN//nW0ooOYgsj85H1RGBJMMHQsmCG9odTQsJ3G4VnCyye8
ym7SpcgKOykIQDi6rYnsg7Mm6DkuqP9TPZHhkaCImVhGChjs86Y/fXjcD3au0NyV+poLnON/RKhf
YYNRWmxTq5VshFe6fVuDdZcmeW76z/uTFLCleHCqQY6NZavvGSK97OHvNVDuaMR7T3lvEiF9GjyV
wrvRTN5QVc5mPz6zf5CCJX5i7WlAIxWYx9rNM6O4v1zeLfHhK2TdHQdEdPJkCPKiKbOVUFon2MqY
oXpUw2Cz9QXrml+h4JNmiRbzSqbLM5BJWMLjkYtsyU+2TbaDRVlcE9m+PQ8IFtx8gXYADUWrJhgZ
W9UYX9quaLVznmrOlPUiubhuEcG5xn0RwOUqBznKW8lhcvGgYo75JoyodGlwP+ns57aXLH7hw9vo
phE+H+rzGC5bn3e0L1/mFNufVv/oXqALm1dnP6JfAjjpv1o8TS3eKdGqPtzphhpqDYs+rF5/DexZ
JxewnHqmm8iUrcebByJ9/5nx/hw6pO1QAY5r6zKGt6JV6Wegb0VHBALS3T1drNZyW3qoETcTLCeg
xtBCb+iQsMLB6w5a+jZ4Zydnji9ghavNj9qKUonDmi3JPJUoWjE0MnbS9G9ffXjrg0s6jHCW0TDP
ZJfGk9TN7TVEIbuV/482Mw4zPa1oa2eJwFvuT31nmDiEVhwBbUivNEsqWQx3dhiYyIV/qtxUnlWS
4/wVXn42wAicIz+xY9pfaygxNSmUYjx3yG4zSa2GtcyKPvVE9CD/Ivt8TqyazU31kobpDelBrve+
DT9p1Jb5pVFdTTx6zU4HvfjIl6iPO66qdqajLwUcingL3UW+UcvWvdL9n5oWDudpTe2ymJSQ6JRm
LxjaPvWTgmRyDl7vISjoPc9fq07f6ekYOEo1HZC9xkLmNSutQNbGI33BQjfGH0Ie8bUxt5QvPtWR
QpKHvlDSdqRMyxk6tRYJPVCKwBRzqpsZeGQucEHDNRiW4L8STiPVeqh6BMRCMZbMQdW63mR7Azi1
OqLf+e2P7k3nHy5SOTaV3TqXfO14mWLsTf20/CWGJ+lUIUnp7nxZQXGwp/V/1ajwn+TeqsdVgEwo
8X4+YDY+IZVMswYOU9uPxY8hohwe30EM3lj+gKkJKmHuDgzmXUAxIhDUua1/sAWmxCNLFA9ua07i
Q+1s+7LubOJvr6gLGHSI54f7vxxOAUG8X9ZnGQvSidEbPCWMf75LNmFMTExxUsJovWb0oYFYwGnK
zq2CQIL98lFbJrlLqcFSJHESdyoEsYtez7xa460CmEZOQXNktCvfitM5cG2ydAAVX5OMLqMUzTSH
CKsOViNPjbL8zesmILOBddXQay6wVqC43F3A24Yfc9v6IXpa0c5WfsZ2/XePrMgeTAbvdZderZFC
A2hN42ek6JSsu3WAkZl1p7nsA+NjIW30l9at1AtsTTS5+H6Y51UA0YxOcfdo6mx3IIxp4l1a64FL
eX5YdIWEM0o+tn8MrhN6h6JATmaM9sXoMQJO8kCIgDXaF4Y=
`protect end_protected
