`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mBAyWnpffJBg6RsIxSVtXfOFT8e927Z5oGbLv8d6aqsoj7QMTyR3TW1oZ2Z5Z9vo/8KKNjXIPuEQ
PwR9zYQrHA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Eyxc97bRAwwk36zty6+1JVsjPcjrG1p7IB8m7Z6yQ2opAGoqqEypLgHR21O5mWoYoxCMQwdKe2Me
VzFtOfKNJZWjjMvgkEaxqRc/fQDkPGqfF6Qr56mvvjCXKEDnf3bd9mGi9SlsS7XtcakhDsY/YAiz
rKEIzHszUToflDNDclU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ApMKGgTER/U2YlkdleFC5GzRbRJ2og9tp8PONPNtufQ3LX0P2JDZbH4PMSISBUs5bnEnwqYuzBi1
Oa4zBxRSlEIAB4pjToBdJ/ANsBPDvukqI/9b1ih00aQArADWRItL/E+l2C7KQMdn+UrmUc00Pw0o
hQCOUf0IuAWa0ytW2yQuDNa5h5Q8LQvuC9pt3+DN9xn1XWCloDozF9qcbFFtOa6H4ob6w8J4b9BC
Hf4xuxnwBUZPQz+4IfuBb+dvc/LEvjau2gJ+80b3Ggx+RF5FNL3GNe2UR486BTPgZztsDAFYnQOo
YuzAfPV5DEkDGSP2Gki1EayY8QjUdgtrAjtkYA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EhoI5pRd6Gu2HtCMZCL0J+UArQfJyP9Fy444ySPF2qjz+fyLqXFcp/622Iznd35CkMfMMtCTmeMC
CEEP+qp5bidxmUbQp6IVRiqh1FrPBjFJUCqm/G58SD0it8fzGTNrkliIOuS0Kwsbk9rjMqN0BrUm
9zrzZPtvRXumkBFeTDs=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iZgCXagSnV1Gs82hZLRRKPcJ1z0y5DkEfBbsdMUPXi3TJKDqjiBshMvFCka27PEXc2JVwd4O7PCL
x3KxBnqpj5Lphu3r9D/bS6kA4XNKJXB3ZJqZIySZc54xbi4nJa1f65BakB2Q4gLNuWDzjoXbHA8x
tr4Nj/yx7K+1zII319hNZqA2mfife8bPF1Ln2OYx3XwP7TLMnBzGutzqxUaJ0XUV8uyylDnzHBFC
Nk7IrdgoJiHSmFQ2AV4BGjUxpCthZ2ByJcemLGvM8sjcG0FIeYujh0ab76q34ZELayfb/CYwR3ZY
B58bu/g1K5e6prwQH4uZjmh6KKtQJRyGwmHw8A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 28320)
`protect data_block
ZwJqTBXJzgkqiN9jkgyQWHo8cXCWIVdB8a3I4MOLoYgountD6DoeTDAmgChtCcqjf1y8YxCrpEu8
G2E7Y46rmpQe1JeMGC5jCtmzCMau2N+6nAJCWIsC0CtFT/gE6wkDhhr8c16Y0WQvQGls3YrhQCa0
8yiR8ZN0tDmzENIsKldX0SIa5reRhTcI+xHhWSOSrcegRtGGE9InpgFTlcQCDRz597muucApQuAy
BtJViTgbOjGGOOEO1gnzdmIF+SJDz/tO64A+aQRRJPrzaWWbb5SbFuTLHuISLbPPtCvwbHW41sY3
2k8hNQ38pdDNbmaXR9TyRwqBtzlMFikLOccnG0S5qMZyMlEVCcEM0AEy9HB1CCDmGxLTQD9Xxuf+
ic/pt7w+mAAHHNOxAFaN+qS2fTow2hHgqkRORd1o6rskYuCKf1eIPE3dcAmMdizCIPXwhnXKtCZ0
n3V8UZLJR5YyRI7dTd6gl7wPS0LYeNC1RhDiY/CbEcR0vZ2SUSLOWKwZqn6/38ojhFB3vY/Xlhhi
IlydJ0vv3oX0ySK1WIneyDfqmhKdlje1CU2mpUhFQnwLz5ntF6j+ZG7vSrTXEP/wRWtxmohzgz9D
85HJycvoGiuZ5ubTppCrNG9h36aNRXqPwKYs+obyNKNtsEvJgOdFNifjZ/fu+TLXgskb+mFJW6JW
99Cayjcse0DoHSWhEpsqZx6Vn4vPoUkAJcZWXUJDtALfehLHUBXlENvJm6SjGhVDWJa0OgGFtaIt
X+8l8RJGMGVqwayM2HXB5w12KaB/mqf3foxNmZF6DDcfLKI9gAa6FP33osSM7mfqgzDSihrmAG/Y
977H87Mh6wRVeBKJSXFGyVDRMNffQRYNB+MlKdiMevyjol01Z6huR68qTOGKln6W+t8MxDQJfSvl
HVDDB0YJtxd8qHCstzvhKdiBR6pSlO8Mf8kdvR6g8s9fg471+ftQSVH1ZU1mRy9oo6mmEapN+IWJ
nOAwf09OATasosHUESwLWl0zhXFSMv9B7sEx7ITJVIKGyHaDKjG0wEIpKmSnY5DRBlksDgK+SY+w
f3ZkjC6Vt4I7h5md1nnykntxc7OjhrROFSedZ4feElG+/0G1/G0n+F2YcbFIQHuL+TWJ3qkhgU8B
SiAqMr/aRfNa9jtu+/9dEYL5rpkTl0e2XEDpJ983f5EbAUpdgQ/mKOWeqScv66AyjYoF2+Y1w9jR
tvxdZn2rgN6FyFTPp6Gku+jZvjiSFe39jPiDELm7wf1ymQse1TsayU2h2c0o5wgICLwMnY0E/ogh
bm91xEM5d+mnqihOEgLQHuHFLGj66eAbFw81aiWgwzkUFRux56AEDF0ae3fbdVh/Z7TMtsUapEPf
dHEKmZpfuCbp50NflCpomqXTHGFfVVQdU94z9q02+Kac4svEA//3QH9pwiX7qQRABfLCJwuHo8Vy
ca6EcFpW6HjLBqH8xIgepas/CQqVjQgUVlxSMPEKRaJG7Ox/hszAQmSFABOuSnglykrvyBbeVGPI
6eNF2Jy4Z96GMVSOR1y5TeHH9Gq9fq0JhSBPMHfu0FDM2AJ0wpO/V2wzL6I8/TjDN9VeGSX2FIgU
Dl9J+HXt4OvwWlDQtdpuWFdSfX15YVCQGtvyAz8hT27XOCmyix4pbBFATSYmjjA6t4PaVZp8FUpg
biUw+/hG+vtUN4J/wsuQYXy6FJoK8wWPGzNt2pYKxnMcEuscUfd5FuzjEp/k1ozVLxQmdvW56m1a
zEWUOfbQ9AuIlFGxefbcri02CfJsd+dZK1L9ocZbL9TneuoebsMAGdUZ5lVIj9pA83z9C3Q6ArpI
rudyXblPOrLBR65gu/mXT5yA7L0xaGmcHvJj9IT+kq7o4yzxPUAqIK/2JQylO6FcAUrOYguraeOn
+4ijVs3WI0zku10Am/sV1KKZSfJNTAhS3418Cn37rqLuqnQNR2HBhJFRq6of8xhrP/MtktxRmPGu
XQPr/B0jZkn9w6iLi1zLbYFaHMk8YN47XWhP0dRS+JxRBwHZuJQ1icPuEgYwS1G0amhClLjbtm05
uI0tetTzbBy4GY13AJwV+LqIv0rP16boz8tk7uJPaPWbFqo5t8vTX3VuFScEUYoIszWPPP8sBEOG
t/1oeEtQMygq78xF6JsEBa+oVk6fBYsmBNoDPnhYe7oinOP/8w7PBJpRsyKh9lyQ1mHsk23/7npA
B6O1L4oa7Wbf8qiMm9orqFZqNRmio5wKzmQy7VQhXUDOfkPUX8bemCPETk6c0yytz2L77WQTjJet
/IQaSnh/8DoLyaxywQZ4YzrMcZ+sR+hMD6Dzgt1xAT3gfi6NBjrqdG/sndUqNk9XwMWbyxR0p0Rl
skKGrl1lOXCu7nzqiXFRvzcWMLBZaaXhRetyLrqPa+rrzzRM8andP7bSAQUqRN2YF68YJKSouGTu
7BAfQwYQJsDD62IcGIBhqmGrm656qqisx5NdDY86AmPupVUWPDeKq2pkNHjZRiBTLSahjqALqs+e
be8LOitCAvKmvUFJWG8fJhd/lQ2Zy0ojetJYqaPvnyvAHoD2Ih+UIeJjrl1bNIKOouS8VVs9Ch52
pmItskkEueFssECvOH5DrS/LcWOGWqIhmaaUPtrlOcYIFu8OSfChjNUfovMIiWWHaLh5wWC/t/1h
K/JabXYPCvpixpxaTGu+Hd3/ZvpzAYNuc24GBptAICiU0m9s13v78lWo7ACzs/oBu/w/5Xw1wki5
wXkvBEzy+GJNacyfsg4iw3KxL1XfiIhSloC8tWRcwgMik2Wn4keCx7c3qAGuknKpcX7i7UobdIsv
DHTCHznunebb0MQLhgEu2sZYhZJB4zHf1aYTi/8KbvJtypJtXNcakWWRFg2m4lpKaGECMDZTxPCN
QlVPggo5iWJj8HQx2rSVj1BF63GzL73a6LUdhWkpSH0UnSbxaNbEaL/T4AjVKa/XVgas7Shjje0/
6QT++BdeAJZqLeEQv4d4AE0XjBmehXaazEW9Mnvg0QDgG5ToC7F2OSynHXKRybRjS1An5wFUCPdW
jp4PKCPWOMccCoqDbVCN5ncSa+wdhBXG+0Ohpvq0ZqgzZUs1cSAQ2w5TqqA8Y2rdL1xs1Wx6Hr7H
uuwcMNZHnMZOl5bAFPyffVWGOiLO5bMwR7STRgBA8Ew9Iv6cl8czws96p2s8GTMgzYjVEcNxwpaJ
S3pd9Ojunmv88QVIchM0elhZbr7A9bbL3ljRgzZ72+FoGOM6kwZrMNO6IhVqtpu8toEcdIXJficI
aRcKspbJGBjS+zAQkw6OSsZ533jzLBrpQeWjE4ZO+62MItg6RKy4FEbW4vMx+IgpZjflbFxAk97k
T975olKT7KWziXAVizWdSxwHF4eGj49SDnMRSIozYz5+GXENjFNEMKiFgK3L41IMPheKru4BU482
alCJv/Xsw8R5Lq6upuAo8PQmSNNxaFP9o0NI20YLt9ax7dZ/9bq/A+GK05A/BJeVM28uEMSsvDEi
XXL/uTqA2A84/FD+7BqeAglQTkqx1prbB38ZCj6DrxTFvwZDcMRqfa+jKcTvN6wAj/AOUU3qEfMY
NCcScl8qPK3JyTrqEhiJetcEhbSzY8dueoiQvkFVxKYri9iaNPyRF0d/dh5LyL0wDH4OFPitONzw
NsXDXuHK81ogz9ESKP9dAplpaHgiczYTR6uVNXKYXOKWxT7jtxO9UK55fhBp863xEgLeHrJ6lJDo
jxGy4gfPhyUgLHkpLwOHSbmAPjw9V6EZCgMQNRyNEj1ElBmDKnJYEyNkS1xgEfRYlGJLa40l9Ahb
MjHuAMK08kN6uYAfCCVdachfkmTRkiuN/yiXt9kBsvxlZFrS0nUJnY2qCpOjc2xE2UQX8A7bfiO6
tMVer7tW6f5M/cA1gWnH13tvGt4euMvZ/Js6+7sH8r8K/XHJkTdPPIlzLfR4TrlOHfBZihiY9S81
Dja572kwx1DaIBODctJmLGdlq+WZVLTY91Gf78O6IRyq4WqmIjiazZ/dyEvw8obGz7YcaM5JADHJ
ElkqMO058uMxKMtxV/ibQ+4tzOnpaB5WHEIy4EyPKP0NMjDxfNK67W8dzwdyyGvqW5FcoVFTG+23
LXv0p1Wc7lwpTT+IHyrK4mUGGCSXv/rLd8QsbryrnmS68O9Ft8a5M4GmoXLs6dYvY8JgzUVALasq
nVrKjttta0Pm0rstsHSC9GfLQwySsNSfjtqLGiOUdiOIO+gCc1tnd0AP+8fRukD5hw2rMLL109t3
yqU6wPu73OZcZclymGmDblSLBabz3KuRMNG70pox0nKzQWenf4QBGY/PC2O2FUQPuUL50jWU6+Vx
28y7cNMTL2idXDoG3BVRFp05ca8MhgeRWrc6sexwcNUhDAp8yJr40uLdIwiLQ0HlL57fUP4W9NSG
nIVB8HJJZvhImsQi5jvl1Cq2DmccRenvAEOpddd2NQNtWl2fWsNtmWh/orZmO+LydJVLC4Wz9Cgf
XxFCLIkDGXLtVFZ8FJZx/UYRmIlj1wpofBwBQ2ygyngHaYkU68pg7pte4OdIJ26fpU36idyK3N+j
2ceteFGKiMPM6RLsLz7D/KZAYiP3HN92Yib/ZTY0KgMNfRKhtgBMYA2AelHhnnBAZilg100Kydpo
ohvFJgBRzz0QER2Yc8InrqyFviFYVeAfVfzjyA96VIkbdB/Wu0e/WwWbg8b3H9HR/qLS5bnWtPX8
856qb8KXhxD8rwyDi3EeKgFzf1FTZbE3WaOzkJo9TMRZLsGSIKCW0TqzRh9qpoMgLImjmadEq9bM
9NqElwwcxDVf5f7e43jOgCG0YodHSYxfKI0UfBdjv5YxGHxfMPtTE4zbUbjKEBDL5PxnRf1sMFHg
aiSOYoQZZsL1tQcLC55xWV7xoz2zur8Xz9lOpdQS31RwELA5gFEeM74DgwjKGF8B4jlKSWgsNk+I
f0fMcpW8yqXCxTKE3l2mM1C5ELD9KumyzS6oWAwjyzEaU0bX+imoTPeKqCyx0yMulH1QkG8Dv8Ww
ykmRUTGMFwakh0qSl+cTS9ZZzFCibduwZftNBPyoE+qiWxg0VYLEZdnw9EhRwFKcObHV7d/EBze2
MH/NfoRFf8A3QhiesrBnX/lmUH+p6pt0wTBQMmrDnkz7J714uUdv06E8rxP12n3DU/fCAE9nxIGx
z4OY8UP/YAjrvjT5y1jrLY7YTktavql8gAmHcc5Ca9IpamkJYGaX+4/8/8xG2HwNwtjY0Myfo8lm
NQhB39TrkWGify2I0AL6y9mJESJh/zwGLT4r/lRWTMvwW8YLYuSzUWFw03mgVk2fAjHYmvKclAyC
UUC0o6xWje9ZYE6ER6psR1vIFX/WlHjUHST/cHyt6IalyTwRgc2qxi+mIueVLNfrVigvKZiBF04k
lgzj9IQLChwWiMxVQFW6vrSMTrVLi6NJSjHNBgkQYWcyubb+47KPDQ7GnY2VxQmd9tV23a7ed7qV
9zT+iAs+NRLabmjAUTdAsEukQQVOXnqvqg3lC1HPkpJO15iUHkGlmLj4lauE5+U/Ez4AWmqdsAs4
yVwDVz+RLaUCV4hFOIRai1e9MJ4SgQ5yBLJMAgFzR5U+VRYPn8s0/j942Bj9BIwVQL47KsLI7HUe
mi3mL7otqWXTsBWjPum6TDWKb2+Rtz7nB2ghK2aqcIu1NV+DMipaUgigH8phVFx6Xln7Ami/SvbE
gdISZOdZiIeSYAFuBwjGyML6JAjxeZLfaRshsvrG5XlY+1q0OhiQO8mN+oY0VP72M0myPbUSm56k
AoaIpcB2TFMnmI3414kshsVQnyQqOqo1efSZXT1g0Uwe0wYET9mYgSDMNXKO1nHC+WhWt3NLiGnG
JSpT8fs8Te7lASkAJaFiml3DjgRGHG5wvzQjIX+CnSNv91dggW0i01zwMsO30eOrS8Oi4CMcmz3I
xte1kzohEaZUh6DwW4fD1a9gmFNcxX0SyNvVLRilBV2OshDGGZaMWaAQFRzRkPSE5Kk++kQNLA8j
OFptlgRJNslryONJ8jWwggO2IdY7iZsDQC4WaspgIOku53FyBfx0ggNJO8jHR1jHwi+IYehKq1sD
wtG3WRdRYLZRC1Q7mAFGxqpz1YU5WEF24U6LSBjy7xc64yTP6Y9+hwhJeoc5QtQMQa/45j0si1o2
5RbkkOKzyeqHp7sl+ehaATw9h/Cx8OKWUtdiz+vGgzL0ndNBuTl0lUf7KCh6wOJqmOxU2LrULcW0
WuMaB79qy3wY79Y04LWtMSdmV98WD8QQDx65POIpinZ/Rgu7KhW4sAchtvVMVbEyubPy8DffMvU2
7kGIul0nNAL1EMS8XJxTzbOFqMtLXuiQ4+mDIQzIxyt2JBrumLS2z2jdpoHjSp6C7X/ghQvkM3im
0L8PMHdR75BYV4396dpX2Qc94KvTsnuAAiVjyFO/Vxgu7Pq7b7bP2UfqqWctWqo4UD4UWhud9ZvQ
Z28VYxHTd2+q1hjyoBg2hOmsDiWx42mLwpvADioKf17l4EnqPkUPQaSoCmKDdtSVKhKfdkxrEiaV
gHEU6XZYdT86vvzfsS9H7FC6yaxbWTGLKG7HlpLEWnMAZDVobQ23jUFewVD147prbinOwhq/ICxz
NAZYgh+fI8FbP7ZzJtuw3EeocEzWWACgkbor2qXo2BP2Nk5Eg5PtSUPZD3b4cWkLKqS6PzjSpm9I
38k2rmY3kO0iMmFfatgisi7eVjfZ/kMavplqQc+uEVbCciBaGi5rTm/uvH5b69lzdziNn57+IZT8
lpIuMfSyuPSoknapbbfQXXhcvVfXHay7P7JDHmS5Cqdfu3R/oOHMRMwJc9KXEagHviJoooWNAHuh
wZyzsB4MShSqyTrs1DhkpH3pdPmVK/+2cspWNIsF/vCOC8AUifBzuADQ2tuuFLL2wcHtAxTrjFOL
f6lUE95em3QLgc3QBMaL7DfoIN40E4Mo9OpQVOQDg9usnvuRkQLjA83nw8ZcvqE35aoejnTr4syB
RrnB127nnEFhCqgUb9gLpRfp0oVtNWrrGAHSzQKNEUsWRTIU/Rmm8oN5Nu2qluEEbeaHe/yofFN+
nP4YISoQunkfVU4BSCEHKgF+b3KQRRDjE7uK9SYwbet1NVD/N7VRnsadvwOQOYSrRr3lWv3Y4kV0
TianBLi0vOvoWgYfMd2wPjkIkB7fLWJUVPg3eEylYTviLATHyZnuaRygb1UF2r65buhu/SIOx7/w
hRZZILMOqitlNjkTMKnVD2XfzD41W+qoaGQ8/ueInyh/+RYNS+Jjgb2//mzgmhgOH17x6AzpXPIx
xvzH+PciZ579kA4M0+IOp/kZdNKqt7Qc9U6bXUBcrqepr44+CNJTKnxd2CxoVTXVUF9ODc02APvI
YR/C0ct32ONiQuXnz6JQgIp9Fj1F9GNaYRrRmv+VNFRv2FZmNiSKtxX6O43y6LEE9GkVr0OIsjs9
ByjvA6pTCSfuxabXof13uGnYlla55K4Fq47m0vkfSwdXsufSSi1amuVQjwmjhAzkURbiiRIUdXQ6
ZtR8u9nAcfHPUe4OD8VPz6CQOic1LBe12N+EVPNVYqdwbOduIAW3zVAmCArh4Tg2QnvtE/IM9FpU
pP1D4TmKv2PBLoy3fZ9DkJiRON3q5pp1u7BGoa0hJnOF8AAV88+dCIAGF2KHLtjhImrhqFsB0k20
IkcbquPr7yUsdRELy3/EmgCXEwRBVnC+qol96Bwkorx2d8CvCQUt4q8Emrd24Qam3x9lsABq8keh
yUaqYzMhoNhApdTZTK70gsAYAB7CSusqJ3uBOf0/SSYrVzLi+JdS/a7DqZsT0EA1OL8eyaWezNz7
XyKdw05VFwKa5dp2fb8tJhNyeGWy+pJSEcxpibug+5bWqcEvR81IlCNnSiNHEEZKMTt1onnsuZvk
t5h+AHOrEJohR1+9G2rAYvBkgpGWXDAFjVX9hvXv63146qMbb9MOCDufLu9a/4QAL/HXgHBgA8R2
XiZ9QmnIp9ihyhoQnJynRFRbvP+Qyn4gtfzEeTt6m/GGHcQDytLB9gPLuUG91i2QmQ9vhweHFQQI
w1PNKkLs8Wzf4/P1nPYwi4t6Seob5xz6u7jG/TUChJPT8cL2G0xhD5Z62Hc2reGFPy+GjXELXy1J
WGPc/zu9NLVjpyfaQP90MhtJ7UinoSRrlsTZUm4fLT/rftdQTz2DcxAtGgSouEEPs28MTUewOARF
WkIsKYQTCXEQSONHgx3uNR/vvncDhaJ99K80tLVHrGQu/gTRggBLpI6Vx5XaWizauC0NWHWBK9uY
u7aEChE5i3Xr7j8g5Tospjt0dzzF/1P9L16lc/aE8us9GJecfUd/s7sllpn0Sy6wdi4AwMHR1f+H
pmEfJYlm4ObNLvfGC93OcD92EeIzybNfcpy2vH5gEVNhOlfFwB0G2pRc8iH/LEKYhX99EadiPq8h
sWyl+aZPgdr9mLN0W6qIMQJzYdR4hieWRsM3TUdDWaTTvJYphgBW/NPtFpaHyEOKg9Sl0+zHeuKz
rFYWi/qHWfzQ4DfqycaL5r+mWYyEeFj80xII9t2QldWJUssZNr+uULcxUqGaFqxImTZZhlsUBXCU
gv4c6NSQckb1KqMpoYylB9ed241gKI5MpecQ4wQY5L5nqaXLhmL98mz/MRWVLLOWnvy13YL64x66
AhDxePn7vR92oUGQm4w80HhuyuXW9s7S2c7OgzdGtg4myz0FzYfT1R1QXOxRHgOgDxOYRph6QvCt
AZYfQGp+CiqNkEsEEwmPPcQcV9w0RjkkMLxPJdlYQKASrpOfhO7D9Ma3GRgQ7aOLCBOy7gihkR6E
E4wkVJqo9BdIDCI+7ItD4EitjfyZy6iO4KITYardCJlYUgMtDt53CuxNoc7/pR9tu3W8bVKyMwXu
POM6UNriv6Ep4nGp8bo5d4IQLa3s971Ri/QN9WyNYAMxGPuQQcd0lzoJBFipB8IhKDy3xpHfOfna
tfgSB722c+WmfpWp6q4juuCylsU+rjNxWwhRWZmZxBpYujk34SgYJC5UKvA3cVE/KV1ssBU6/9qV
XKxZw0bzVDCwxX9Vzr+9fenhIveoVSS+6g6Pvg2vvodYpuTDlzDkXaMrQdIkCj1R2g1WpmcLQRel
Be60Qiv8I+eNMs7/U4L6qzS7gI1osyk8c/a61Y5GM3o+hOT3qgmx4Nzp9fmMNWi4pZA2ynkzrYFj
Lrb1Oei20lORihgoxHFbWcNDuldGeLe3LDOCLZsCy6udeKb8vWyH3U0Pr+8uDqbaB+JJJGsdoBC0
Vk3kFW1sUm2x3rgoAYDzPpFJTsMCFKV5rnXwoT2W5kHa8G7LArcwhLe8l9r/USiaZY9ulnbAJ1wa
nORjymE+i2ruEgmf47rB+z6qPzjHVUmFMwdspbt00dJ5dW4NWMmO8R0BaM3pIMVJhEAj50CMS5d9
cYJgLGz7HSu+qBdcNeBJu3mxYHuQvNznCs/Zk4939K2BDCKyPp8aWFt2MkCNROMqAd5pjQSdKWJR
HZybuB448eBc7qmEKJ5MX1lb/Up6PWOpLtL509I07d4EHb5k8KVoWSobqkEWDMDePSVQYJE8VwGA
EBt3d2QOwxOHysm/0r6aYfcKsTydoJptfPkCrygdxQWwSmnxjAUxMYHV1r4gjPtgvPtbpDCOFMG7
jJSNok7SKYuXapj4w+FrJ9KQi4OIYSEMp1Y2w4fjlM6bChowZqya4wuhnAwje2fa5Ky6fZ+th833
Z4fJrPfaLLQX1DAv1zFjW3Q9pRREKpGhZy2olFpbJUiIGxN50VbMoyxRPlV8PR2nrI6ak9BBkyX6
vSPfvNAAUxNM3rSTCppYsrfunzemcSbMt0i0Obes+xgGMCKCRPW/KeqqLcU5DeUNNSUsN6iAfKtZ
dk7zaZuqHEHsS6hE0poz3gdVgAX1Gq578ZdG2dchh8F0pyXkANAhZG5KGx8I1tX2ibHPyK9GaDh4
i9DLmESM8j2fStl+dMn2vLmPOLFVe4qxA+nJmwRHYtn2U811K/MaE6sj9krak83J6BOns9B7xDcN
UW4GEc89E3bAbp3TmWBHblq2H+z9oeIQbxT6MhHULsAXraYC8NPefXchsXcJGhFe0ASr5SlyqRIR
jHgvVclyoJpHT/nQ23oOr13E6Te37+Xp75UcbPxdY6lxXm/8/Ik4kcO/kaAI8yWJShK93Z24kpg4
YqsPNavPoLZ3zd0GmoMbGk4FbtDC4Ib9bTHqfo6J6v5XzBgqAME80QTtIHMr2e2ukzgiSsuOJjVV
2xRbvNM/+WgmNb6Ahv+lXHBGqJ0uV2mMf8A8Bhe5pBdeHGdLs6U0WwpijE2HIXZw9ViaCYJRogzi
c+VJyRj0dZqiSAHq3Xeuhma14cUuvxxfer1VHlL8/z6o6XJ19l0IYKa86WME4dzEaq5x0iwN1JTq
rBek//O1eVdVNYZjBJ8TZxnljdg3Ga3hqqp8f2rVKn8vlN+GOEd65lu5bT/TRGZSzpYaNNMC7+DW
Vywqe9epOg6TS9uknokosMFG2Qt30iTicFrID4zggEDRtBB4M7ooDTJDjqCh4BoQzliXAqCrRZSA
x2ygYbKygd8qKsbHOd8Zr21Qyucjs2asd+QucBkhegV6rv+1ADtZQv+Oe9j2GgaNNIIPyROsjQY5
azYBaw6bDykk/voJWEMLWqSYlDZlt78GgSIPWS8kzCrxxB01rXasN4n6rn3zYqfW/9GnRbX/mvyb
+/f1rA/4Ui/1i6TatH4RebpUZZrBzMGP0oxBq/aqVEyeRS/Z4BVEYS7rLLFeeObdUQxnzi87b22s
DDQgO0pKiVNT2X7ee51IZ2upmOwrkqW7I8aqG8pHupvztEOt8LmTqexn6txCeGXH/JJ3JPMa+ZIB
6YMuVInujQtzV4CTMabNyVnv2ofU3KbC3NUZGnBUSbW6tuqv2tpMeKCRnrZGseYnZgtFnmAMF8ZF
lM/2KDf9PF8JQe3cHc0CcT6Tp9htVP92MZRHEp0w1y4HI1YI5n2IN9Q6Bqx9e9l8T1WfoXG8IGB7
47RH0DxG946O+/YG2HhN2HPh7x9vYRXzG92bo3F0PH/qHKOsWYY9D9lHV0DfsWV7eM3YfjA0m+1i
jixed/AMQ3xU/zbo4saYQL5Ps1s+GP7cZTlZ8w8vmafMBSRWaAtXDLGeQcyjW302C/vw05coq6bI
wGIfHm57e0xcGPv6uSRS1SW2jreJrskvtLPMWoRbRGVG/Byei0xOnSuIcWxZRV4VwEX2MjgX2nGl
AI8ii/VXMx3zNNYZYrlmRguEG6bMib6t5RhQUeTVrz3i6GKfMzg1jmQ95G36xWvhIpUEZVst+m3M
czTZEJVoK30YmUPlePwm+vU8vz79p5k/Ge5jS1zjoWEmgRSTmGcYpa3r/s24G8XafMuwHhP5yC/t
yaKzoaHhuYuGBEoREM0yxmkxkOfyro9oTAFgz2JHIOPc+QdcKkcNknI+zgOTVQV2Nw8ATjLGfV5Q
frH0P9GBpngmw7eD3QCZ/QadXyvWdi66oIW0B1h/S0lv57xFB7Vcn4Btg16g/40WAPJ2/lsQzRao
psxVaJZml3ybkW0XpIiuLMwL9pxpvmFlH1oAz/qvfzMwAXl7LSPVvXBmk80npAKXfS3ZQWur4BJt
8LHCjedW/h9L6OzhgzOOl2DIs1tNH0qgPdMUrtEQ/HkBi7g3HTdNheOcmTEnbX1Ybvri5cV+7iBr
sUGaSHYV8FE/44BQeYUkh0OeI+2Csg4xbsSL68CJI3WaU+lutgXP+YwURcIT2ukHPP0ojs4f6EUL
YpEPj9rAUSrxmFP7bhUIkxS89rFP+qCmwIuhxpMvDPTPMPBs8/Ww4jz3YwALJATai6nxw3+wGu2z
gTxrS/esehvD6twrXk5MeWEpx/55G1Y7A++ZihylnkImVdLYh5ovqPicIqqnA0pwy1hYBOrGvBt5
SbovxJ0cmmF6M78txTstbMp/Zi0sti+F117B1fHvt7/eCYz8htry/qHtTH6HpdPnIbqoBs4Ge/V7
aSxJ8H2COmmtm41X0aNZxc5v/CXSE+iLZtg/alzo7GQDaDObRmHA4gdhNyeihcVwAJdLzcLu1szu
rbzEPs3tKMr0eF5h8zAc2l3nmAspbrnDiJYFRTxLUX6JtZFNDYFGsO9kPRK0TmDYUDoE+NZq1mpv
101uKkp1kggjJw7eV5MBFKI/SHTd8T18/Wkh7Q+CxvImgokak8dZlHV74wCm7LJCxx+j6Pv/kzQx
CuBpJJHHR1cWujzmb3GwfjPM5T+KbkRjvVG3Zul0dj5yoZ9K5KqYr3TozxVjJx89nnUTvku65WDr
O9xUWSjoe7wBJOdHEoS6BL0Q3qsockFkK5MwBqdOjfi6hFKPEeL2JLnk7lDfUqF2hk5A3RKCATQ+
PmR2JozDA7fg9EkgdmThlOvy7Q0Z9OaE5c6OvDjZ7AKBUHt52r9Y00n6eq6CmVU/hUFeNpB7N9UZ
U70G+R+x9K71XUpKVQu62Ha0BkPVSmhJNKv9GFudceCorEJfLdIbSeTgsCb6ytNNF1zNxtbzQSp+
V+b15wEI4fqyD5V8QZNy2VsnNFT6OAAYHeDS1ReO0rYI4E/Xu/x0fb1xG5Do5IKfcDp4BiVkmrSr
b8Yqv6wAyhJ0WS6mu0k1IqGCcP8lPyiNyufq3gUnveHMIHY6tfMmPma3b32IrgAKArOf35On2jW9
s2J7RDAs3mZHSZ+/ZZ94kTYFj/9bXAskWTo9TjZh9AFKiXj55/vy0gYiPlUtYRHYG99wRSNC6bx4
RU3eqhrQ/2nau30pZZUZvJZyoMjWIhimrBuCTXPAl+MpLg+V/uOUWYF0bqNW/1jWiIlpNlgG5RTC
x5kzYHMqAGxuisrWqCIitlOVKIzlYKdKUJ/AjFihPe+p/9687eb4HT/CcWsCGlRYL8+gLTZ7ZiXn
UouqSKnMJoaQ277UhN9MHqiEWLqL+wfn4+1HM7qbwSjYCqo5TDekb2c30Q6TZVGFJ+jRsUEHsqq8
Exlbt8LjEjvSaPxYa9a5lVQjbFEAGx24nKgXANJigPnZJZSj/LayFUsc5xBMGIeaS7s7Gbi3pSUf
a9yKao9Pjx0tcgiv+GzdcF2ioqJVdTKR1BgVfKRRZW0UBc+x7S0kCufo/jjEb/1Y8Bt9QC16xRXU
nJf44YhrmUIcud4n6TaDD0jS2RjoFkFTd8Gk1v38l/FiiSJWWkoO9kUmBqoLm/nNndt9aWQSPjj8
Ee6oIIX+lVC4o22rAl50yaJ+Yiwu2jHYkJS5aK0syGSAgjwENme7jK8EXQOnmQzzoqaa+0fdhCKU
w2bAVzYIBy8OTiEkgpCDqH1ruYsKQbrnBzcXPKS5mUwESYtwm9mEITDlJiUmcIY9ubFTXlYF+yTC
/tYp1iHwBLshm2RIA6B7v7pMVeBITTRHYjFsWHy4CS6Bx707R1ONd0tSZUprZ7ZFNtUoMOWE8Jjq
Ag7ZnXJ/c+kJYhL5veMDRM44UVbCA6y1iGn/3K++AV8A5RTn1T/5JVr8l0TYYmLapW8DeAENiqxU
2/traNmz098yem6nvZ6gzxJlDuk9D86EUJ3BShZ+fR/rI1lvvbiRABdb7o9DttQ77GgZyBsGpGZG
tE5zLcN9WwbCwddjnpBD+kar9VTXM3WvXP1wXUKaKr3yYk03FNUJVxr7U5HYX2QEmd+WNZhev3cL
vb4hcmfWdCTfEEim1TyvbyClMuFK2BmBpz9PH0fzBmZ6Gk7FnhAPDxEF3RTJ7Rrf2iad3zRLLfcq
FKoSaLSFSjS7TErA79SwkwT/tmur4PGA7H63n1Zbn7uPyzSXFRJIHjsFbh3AaLAr6ZQYFRkiN7ZP
hJPC4Qn0RIJIXINZrJTTRUgkdBnAeUB0JWjyRpJhSwBKSnij3IjHHqkH3IFEBXJpgarv1P8NCp/W
9mx+B5TCPJNWUev6Fs8I63OStEAM17PRp/yS/FCrRTbZN0jlFgpX7e31L6+UaDA60Inl/fBVL+tj
WV5P//pkjvX+FX8HsQwzmbE73a9qupEjCQXYxL9mGXGXZ5KMyNEzUTF8Y18fKYZ410vfvgFOZ7an
Nf7NQtbgn0bFyZQL+65I2krLTWRuchO97H0Htau5Gi93fynL0dk7rWNFFicrrCmu9rLSf785bcNc
QjOY99QQVc3mVx0IleXKYl7VwUb1UmvBmshzukFLtdRkPsnT0vcxI8ucnU9fbo2i95SvUfAaspkR
vLk7k6ynW0u6oQhID8i8AariggH4jGd59AuKscJcEfryI3dUxg3ymlurop/h/UrZ1vdmG7pVL8BW
aTJ3Io74Aa7/aEjeSq6kaf7Owye7yuBpkfksItdXvtfSqsUQaXK+t/TdCMm9bvTZJ2g7k8LbHzOh
mj3tPVX5UK7QSRCn8c/Ob2/d54uoys/VXL0uQcaKno4CbQf7RkpIspBPp8Hb7QR1FODCvKu3P8Qy
tNVyaCsZXg2orzc4Dwq6hYGZhmOb59jY/0Dqjcjnlz2zCAQXXSeaPwlhp7rdGaVvE2ukdacbfxXo
vpMddJc39cukww3iyM+5o6CtYDW8cpE64xXhQmyTrOijCWUgv3JCCEAnH73nQr2YTAj8H2uR5I4v
hHdbtpXRoQKx7LMegzaI/H0EwgxfJoOXveBPiBOJhv2PlC++YglTWUBM/+XHh9GZZaiK1dEmlnZo
z9OXjLWlRQGjDztH5vawSoOgF767HEymc2yKs3RkJKimoXw6P3o63iXgs81PGqrtwHTbFupCtEIG
mJYf4E1QhZvgKivU2SrTZR3Orwq4pOqmfQvCgPKHeorHTW/TQeIUp3Bvwf0nRw/P8dlJjcIbhclv
ICEXfpv04/sdUd8OVzaeG8jWZm+NaQ/oeTUxR1NNzd9DkOg2WL67j9/SU1+8x/MoyOpxvnfjb6wa
Rv+ZDa4qPg5HzjROv+b+iN0etjJbCOIhyepElkV+4joWHyWGQV7+Bm4rMc0xQ/Z3is/PlcGJy82g
CIxKau3C/vbXsv37MXPedLXQEUUbED7doQOzfUa98C8wfA4IRb1OhGc7AATPCmhXhqQBCSJ0aIjW
+d/bx1zsTTxRQa9KChey9N8KB/XECnPjO3jtTNfmYq+A9oHWxO2d6MGH+LMpKEKiaCcJuk53Y28J
d2kZv6Pd0dNoSRqc0J6TF50SCZlklWFhTu8imaQ93hqI6vWY7Vz9MRY36pk+77nqZQSoK9TdsSOq
cJMIKoBWX6DELDfPALe8+34+LiBNsvdNxgLoJD5XGz2PzvVEIjkWAECSKiqk01xcrV6qKWZ+dyte
TYYO6+lTLpM6E+yRG4XJSnGXew7mM96keNPQq5MqnI7CS0U0xcNtSK3WHrL/3GEk9bvGnX8mKqDD
DSBd52LhJtXPLX9CnIlBGXn1yavVO4oD84Qv97idvq9DX6zA328KceNfrCUrEtiSuUe5o3iatN/z
OtLuZ8Q2bbxS1kYz/FdFDT6Hu/noSF7pzHhYod5wPGcSHf9aejZoMQz0182U063VG5H2Wi7/AbGF
dzgvTcC5DW/jbssCOqjbEbNY+Cnl43x1l8htjYEj8FG3SmPMGDfeKIr7KwRap+2NnpCxqJr9M2a9
yIIXnJYf0+z+mOP6y6WXXHt/+QhgCvzVMKW3G1QTDkfUlpX6kMoh7uGSzrZcTRwD/y8JwoLF0jqE
4K57iuNUPypPNCSorNQtvtEUqRKiup4HOYRKzSULtcgmHOWhVVJdl7D4hYqERh9YZWaASQ7GDJfi
Kwdy/QcwW3Yb3zr7o7oNLCnuLQWazkpBAbSSaNiNfXodFdvqK3rCUACVt/6Q0I0CIBTSDYqgqLzW
d3G8b6pGNQEI6E5pBcgU12LjSt4f8S8wyGCe4S808YwPdzbIyMsj7xvDG6qdguW0N07B0VQoJKbC
ILDKodYxKokWaiXOtqq+VgwFryN6WikGdYnwGTjMgxyXGfDLGGMjAzwL0Na40GMAaq/NoYKFSjdS
mYZioGOYUdfW6bZReLKMVYMCBTXEKVAu9/t2Be+PyreHPwVF3rnV5bKGy4KkQL/H5dkMSJexda8z
iIc0IHnJ0R3OnQyF5VLl/IfiVcLqhH3c3uns5PMCMW8oS8x0hrSCFOrm3nP0tfFPPmJry6C2d74u
5uQIh2q7f9Xx5So9kUXAgeTXg/8mL9CuHJrutzT2lGB9Pyy7hhcTJYmbk7fIo7RtDPtgyO+nA3n0
dRZQcpCAUI2gGn3Ym9HnfkeEGJkAeRQV+Om8rfi7v+9dbTRVoOGvCXvWLClUIdP+ZoW7BcD5/6J8
APN/qSxwWvEBPkCXG2SVNAXfWBpTlfQvdjNvZmFXuct5ZHH7Lh/i02HGVM7aNrA87qm2VIcryNgv
9Yb2QwRihyu6zCUouMZg7SL7D6W65dulfiZnPIS7Sant13dmugZ43zensOZYi67lUdZlwhmWu27T
ZzHm3SzQJwwtoXLfx93hhLGjzCIuvZwLgdSKVBLrXbzNBoXxdnApFl5FLZ/o6v6rUjBvF58K+bBW
t7idIXcdhwC/tfZe8a6EUwenstk9iOt+EahivdFlQCKrX0Wqs21KWVvWc+ZEPFxoZv2hLKdtyx8e
DRefkpshp+9PeBlyXDZJnLgcp4M/hkl/337cQ0G93g6kp5DKn6DRXoD+3qyD3RbxkENu06OjXeHj
sgaQBrYJkP4VbNuJPx9IVOP+0NhQfJs+qHfAUFQmYi3VpKBtP8wmwyt4TYAJqDQR1BEBIJmN9SsL
0I/GjcmoY80KQ2mGPNPkJT8CJ313nENrQgGOBgxQ8784JQSURoyK/YrwzU16i8Q26t3zFixdEl1T
4iEhG2Z56FeGBoMqVBPBXj6f21eUbOIZw0inygM0M02MP8IlOwMyxJFBytlMar1agFVuRAwc5OGX
40HZ4mJbG/AB3d53bjuc6NQp2fQ2H45gJ6DzxkrlZXti5kbG1GKZIXUMNpD0jzeYzcRcJXjAAxBZ
CxqUD2TzYMPO1qwHJw9/zo1KvJvaP+GcxdkXRPoNT/LPU7i2j/hbqn8kmlvSXhHgkF3M+Ao5w3Ab
DUMJuGgpSnizUk/FVGUWAeRHAMo9C93O752VS1fEbxmQFC4EQshVknkUs5DF4F30L+rbijjC4Zz2
3kaDkaPCuQHzjVupEsV8I3h7zvRzbiELQC3vbsr0OzLWpJaidAMxtR43fAZGGhayq0QCcY8+KKiR
nFCsQrNF1K0BGQh7A9hmCuYfxv2h6Wr+9adwOZZwsHv+2yVTHKLkoVBL+X8FRPbUxSKOeeNTw5mB
Cpm7PX5uR3CXvyPqi4wg6suX6RKRi17UddMRiyFVQaGzlGiTzC5OEChOMxscLWYgTEUVc2jhBoDn
WSmGsYI+dJIE6OyhofCbOqMlIPDSraU6QPI+Mqwkg+KsVNmJHQ2sZOLdeSLRLR2cqFL2vHZCVCTW
VEUendS1Kwfep3iI8eZk2vEmUhtyEoMX/gIeNWufHLV2+0sLF5j+/PYlgQ72lxxpIii518ZfS8hS
T3uTIQM6J/1uaByVrF0e/gwYel7SfT533hD+cUlVKpCUq7aI7/e7jQpteUuskq6vqwLXU7TeqcH2
eYMaIeJ6E1nq9ZI5HASjqO0xEdKV0BZvW3nTw2RoHc3iQu2zrXa4Fh0GlK8lgbX2MqnLgqzT99cf
+Wml/f3yPqcp31uRcp3ydI0HYQtqUmxBS6zhOQXuWeIWtLFrTqEL39JYubbLG7jB07OxthpC9i3W
k/omShyVoX8c+suvK9WIv9OBil37/oN3RnFvS4INisPKB8KG7r5oCotPPYMx5ltLlSvIeQOKc6XF
I+3ISaBk1PyJTecJiaqwv5ySAJ/OyyXn7lfA+7Hn6jPW5XEcma/DYC6BOwGIIg4tzrNLjGgRZPCB
/tC3ek+DXw2XgxhSusNrFRCH1A2ugOnvruI/8XBaGvgJR/I7JqCtwl38PqYyavLTIrzM+1vnPxiE
VuzXHVxqIGpsCpam9R+UXIcUTHWQWwYWO8M5ORrCyfngf7dFI04W557ewT5a39fnGZQ91hGuuBaJ
FQcrzL6qSXdp+/RtXzorLKCie1h9k0hldTCZCgWip1G5VMDBMjVZCwn7JlqfzNZy1q05jOvx8ZuD
ipIqcLmCFsj7i9IESA+SgWcAoz/1EIBx90895WlGb39SHuiyXtgvBoo9r+zC2wL4guNDP7ygxxh+
6nugVNZH+18a13y7gtvqRnZpm+ch86mcWomQbQ8GtV3qMDJzFAMFSTuXzihpfl7+2S3XifE6rIPH
nqzWzpu6BXg/3UQTdm466T58Sdkxv3sKWNLXMSWKNM+MFGKMrPM64zEAAdP8OAg4KqQYZxtB69X2
LehUZoClgxyND05U1kfREr54FIwC8WBCln66/foY4yE9syr0b+DMOMRgTasqrAqVazzzhVjqHT6+
CIKSJ/uRxk83Sd0p6K5MIAB0Agiep5oND/UF6pwKQRjlX4WS5ogbAqUeODJQdKrnoSN2CtBJ/kif
kiuCnNRcKUapxrj9kBVphViNLBrVljRd5gGuKP8vEX4iOiBN4Jp6MZs3qQ2GM4UeuPEDKd4kFUlY
pCgImepVAWNXz++hW1txjROF85RssPJkKv9mS/K54ww6SCENHn9njHWe4obpnLBFjK1j90/ewqBS
6EOd0SEkqn3R6KZyGwr0fxltsT8SQUCGaeHog2yKW7PTYunUnbg+OQR+yvYVBFkMFuDmz3/8sjDZ
TtuXv8dJ5H8skTDtr8lDMFPj4eYaGkvqVH2dTMzO1utv1vWqte00mfsQfAftnoS9uEZXGqtq3B0L
KeIXMllD+VRPH9lUnwtnBXGvdp4f9hGy8YNsIslWjw1bpgmLESYDDbwqC5PB1szcG1KOlPCbTbFc
quHDHlgJSjUMK8er4wiH4qigStsZ8YvhZT7+YP2YKLc7nXu0AjSKuXkjYzA7f7pwO8z+SUoBEa+5
89v5xGOsK5FoO7vl4Cj6gImD3VZMFl1RN62uHpz0EL5IUmxzBf12u8wXIA//vkvoSRyPJrMWXGW6
FkVsGPpvOT9Ep0QBJtRyyCTOo5wp+8Om9Bga3CbbHryhMSb2Zkxfpe/vYegiWyUeX9RWoHx9WaCm
tacaZYLccgBOpzX2gqyKm09FLCvUHD8Q21GF9QRdsF+D6KjQBFuU727gzu/YrJ8quurM3t56fogr
zjXpF368S5gnc/7WGInCNlWhWytXQNP44xDSWe8x4+atDBGCx+p0l1vZC3kBg5Ov59EGp+LYcf59
GpfH4o9ygNmzNLiKRBjDkC07H1qGXOkj+8zfzGs0RlPn+PnfNrHeaFAXroNL7Qyj25kDVk+n6aCP
GLpqHazsWAsgH5wO/rU0d0kwkWgOsC0GunoRyIeLRLtt7qfkJHMLoLan0XBHISLqw7nABLtcCWEU
CadlVi3HSHvy2n+RPTzwgwhUYUv1eyiKVcoq4vk+0J7LA3UTPwLkPWXxI8XvI/9djhRfi0Lw11L0
w7oK2K3YukjuWjhVHOjGsXpth8hp6eSsP1XLDhhDIkFJiX81/OW/pyT7YkoxRSxLjoqTGUjz8rTh
fInoF/w9HuJkHjuB7LTJ8cfl2N+F/di4fEwhzQ7miPspE9lHJ6JTZEmcF6ZlCGqiNQRQ9uoMvNnN
IQRLHhh9BFwipU22xxi6Mi5bAr40gUU5Cis7L2UKHwauTBISZtlyYbYZ/AWkICJASlrXuiIElh1P
m8pwL1BLMEVWf3T97WuFw5voLXFS/rAatQ9zb4TsG30o7WEQ4h0s0/Gyh6OzS4MmeMffpMbYUz5s
1b1/KOgMZhZbEiM3N03GZouR58lTQ4FphA4pfBsEWAnHBVJ/gTxNGX49aeyTv2FbEQnA3ktSiAB7
vo2WXj+f8WCizP34cMz5MWQeQnso8Tjg1FU/39K46c2qW2sZY+/xOm03tLcv2y39TAUi+iLCa8L2
bQzeOvd4YYgwCkJtxzJFBSouU5AI4CDhmlUZweFhkOrLxVqsGFCARgcrmSyIXzHJ1+V2q9F3qohD
0zmaBcTeppYKz+LrB1gCu+fwUDQfM2wck35UBeywmY2can/qi1KAod0MoZEkclzq6fUlbHAPRT1Z
P4HL4sADyYOjjwgv9UKuQ3zcLaSUSJcoc8/cOhIFnD8FshBUqQhWkkHHzJPnUxF5SM9lNBHqBsN7
MhL2qo2/0SlESXR12cV3RqZK72swtibTPpxCvyYgCgSHOOoDX/PHDbjih7uAFlRNebIdbBkXSt4L
Queawe5Dsl0oQUVy9s4x4UM8OqJ1rC+gRWIP8K9gFnatsK6oCb0g0oeXPRpVkJFZY637hmoWEajz
bkYMfPWGCuMr/mAju9q74+jWYgjVZyafdUQFoT8D+/c6h2kb9jiE0Gz7cJYfVXgkeNIWNgBuvnyY
SFgqBEwd0ZEatA+JN42/j/KRYxYHjdFxaQwies30/u2nb4nyP8tqQhicv3tI4XXpNh4fTWDTKvQP
SkZRCLNHt+iqaM20AtPn7XjKbl8hJoKbjzFvaV/q19ACigNQ5ge48vcI0rwAoUzkB6oqsuLk/ppm
D3y2j4KCTRXOdjUQqVfN22+GpCh73t/lYBv+THgF/d42vTnGSeweGyF8Bco9HpjXlsUg7cy1TQqf
m6YhoHu/RTWFCyL26rU7sETXagGX2kAyIka4G84jijj5LWUdndkEpTc7GoT9AEkq5rl1CHso0b6u
bRUmNMFvUsO5JxgP9wum0iXONtjACi3BGEA1aGAYqzQNSUq6TzQN6247D/iRHWWa27I5jNf4G16y
MwzaWD//7zxvYzDjVXfflNcSJLwHarGyYLeouw45SADk1LHSvGnO5Mn+4KUoIHSyzeH0Nv+kijJI
x4fo+yng9W/EcVX3/KD4i1ogsf5gwW9nvDoVFyWkIUmc+VW4W46smzkgP9bYqF8MfkRduQJvUKu8
/WDBr9Tlw1AgDzirxmEESN4ZZ8gr34tT80vWaGFwg1USW7Gkpu1jqgvJ3oGqIm/HiLZDBr6pyBkl
jXo323TTqNjJVH4pgV37X8wtj5fb9L1aY6Avu2GzNUHcBPeD8XMfaj8/g1TCQ6Y+Cxuu+bwhbB/X
tDIT3pmqSoJAHbYpqhg/3i3f9+C63eXPMw1UBoZ+ojnMuxd4SbapUBAAnt3yUS9MHWr7QvtFEdJw
K3SRyjMWeR9fPevsYeeE8fIC5Y0aa5H1fofkRwvfErgfNQHEJKDAQ1D7FnDlsCxcBgnyC7E4wp4t
AfV/DQNw8V2LIBbjNU4ZAxToC1wg9eR4VVR5tNmLUwwB8E8v9izZZ163nj2h72g8NtZ4zRMASMVm
bo5PK1tq4W42r9tt2F0ijoNctrUTBGvTxoEja7qOpKGzIt3aOpjW2YT30cVOVo7im4fA0OVe3FCe
ddVmOiM0CkCZzSgCEYZXMZVYgpNoWVmnR0s0m54ktBpZdn8wP3nX5lpCkRt76sDeUopW867ZzRhS
1Wrb6o2okdzco/7GG91VX7mgmWwXvzGrNnr8PlD9i2ei7haUIlXs2jTHyXwtcWFDCK9Wo9KT7X76
Q5VlQ9w9sjVpRJGc09GArAdV8aS+mx4M7hvC2hHcwMDlAmwhu78dgDXE4xONvxRwRk0jumJMjh71
4y+JQ7VgtGZY8y4wqCXt/RQpHjCs39Fcp4XmvlzY0yZaYRiAyerGZx8/M/cyCe65OaxCvYMFVvqL
aQbMkAtj22PnzGhEFGhmVxpN06fiFoNgIkAybPn6Bw4Uk1Goro+LBszaCvf7yvEhrvSm9fGZV4tP
rWbDfuV8YMIRp+oiVW4MqoSy+uS4iDYeiQBFg8s/gfYyU53rzw0Ub9NSDCjEurKpKPpv+WAFQi8t
/YssTT8IJ62DKtUGk0cOaeFsUUQeCTYepzONnOf8MYqSJHCH90uRNd2EJDw6vfbyKLxCSebXMPLM
0gZSxlJo6eHe81gTtFqSpu+8T7bIXVfe+XqriaraaJbtkHj8HOWAyBeSQMA5hrw9Dr5SwTK5cb/E
eqUijApuTj7/0B8h9OvXiU18o2uFgJEUGvB0Y54NTEG6f7oCyNF1xc5TZmn5uuiwmD4rHou+C75p
I01Rp4s8QyewKNxtuQsjjFy7++gDh2YwS0rF2MMJnN0L0VSM3F2m5wERqrDuC3bIoAy27dSWECmb
2NFdl7yRTQ7mdKK4WD/jaG/z9zO6M8y4DYoERW4CJM9fzjSkGu2/KgXX63JEElrBhL+9423qVonS
ze1WXoHQeP8oFY1WAVqdcLMlGsWtZ8ORt5+o/667zoVOpaBSZB8nSWoAYI9SowkrOQgoPLsO+cy8
mjRLNbtVWFLLn2Zp+9SIv1rg0WwjBYG4PUDkxhKtUfER0di8rNsliMl8alrVtSuiVCnJOvo4yOKg
wZzw8jhzcmgOfaRahe63jr+MDP6JKlqiHMzlO0stnJdjsr47IApHkSWto6C736BqUDKduC/nwUKr
J4HIkxqkGoJR1+ZPNEixMqSo5DwJXBK6Lob6nYUANTe5Byn8YNTwrBcWAEcAedpUp0h6yK2nK9SP
CZcGXtv/72QoS+SO/eBupFYFRs7xzCffO3iw5QRHuvLADlAbvpx0pH5e1o64HX6jBktv05ZPp9fG
ldqK3O8if3WTx3/0o0PGwJW2ZWQmU0Y/tp0En9FBva6xDDV0nzT4yKWwKwTOOK2RjKmV4YDBZoSI
IQOurTNEGSfAFGkPBfOt93e+EkoLZW4pd6ZtiIDCLdV1edlcN8hCE5ZcESPvW4KIwcsFu2JckEwG
YvGp0hgfZGdkYDY+18DmWLUFqeUDD0U5spguuh4pHaj8uOwdouUGfD2fxWZW0YCm7zYKbiXAR5l4
HZ738LT2e1fIZoAnLqYyNZJW/2pN3KDOZJkPuBmBdbGJbhWGZL5/ZiRv0uQN0ORIR71m2MAWH26c
gXb2wKTgK9pMPHCHRQjTnOhy+LE/Gx4Q6c4qFWQc/US2iLYBsmjHmyee5rmL9Gp+uk+PQqOMAT65
U7EEn+X6oduo9pJQc7ptACH+hoZHcoPF5w8m14NDd3TB8F1LoUsUvaeBDagGzhrqHeKaGX1Gt+Iz
Mid6Caq4YM1uaK8AwzJlavk13C4ll+wNI1Pc1MTfWulInajuSP9YDeHLrZiIp7UIadIqKMcCGWLi
L3uzHPZzSExo5T0hmawxwMYZ7KZAP72BU1kUd1bxM2KLrgaUBVSx8DiaeS5NCIKebk4E8kuAm+As
mgPLBD4jJGipUJLte6QYTo3n0e7BZcP6VBGV/1wvhkmCVzXQ2EmVRM32/5clkive5PB4ffbHIGbW
+Zum1sUoFDM4mZbVRnzMSew4V6SnyLkJNzOcT3iPGpU+xn64/eIybgdEyFztu+liZEXi/YrxxaXF
GZSrGJ1jf0533tqxd8u3Br8HxPsXt89qXBFVqoAbzBNw9RGXADGHy1IdoEwl5kOlRYlesBHiZb/W
eMwM1HvT+qQChxkVQhr4BR3KWRaynsOHdvosdShE8cvvQIUd2gl1shmOA44LUgaTaiagIboaNPOi
by1kGjggUIermvl7lmVigSnxUxIJkSArEXG402X/gIjVwaynCBkFO5cP0Xt89Fh9yiZSbZ3b2hSP
srwGR5hNG7MJZQAByKQLVKwwHNxxBNCHsjk8p2LQm9KiDmlAJfxcaLv5VVlMrRxdhUZRANdqjPj1
au2cV9sMKRjFaYxTo6AfGnvVLjm3QmMlS/XAEy1F8SIW2FC6qIGipyAyvlNtZ6pifkFJneAAo6L0
9RuklKJZuDAXsiBvbp4QHmGbHMfroMlcabfpXQfvY2TwoYjzCzsLDChxY7Ap0hd/BwCQ2NuBOJqU
glcD/VnJ1UOzHHeuJu+dcERadxqW47HDXl0pYjjXQT5/bEioreg+1SnP0Zod+XudGpSbr4gvFmOJ
dJwkv19yBVvdBNCGi4Lywd12mjAsy8ZkZQiWfbfYvmtwJfC1rGTyYACd5f2Ht2b9FG1zqoI3pCsP
BbEKebQ9SyhmgGPwsm3sap+W/PrOKk0MKgBCrwd/Qp6uzFYFZnjJSZKUBnk0bD6Nr8N4pjxGD/Ad
jJvyNLJq/UHkYRh74JSa32rZGDTTJOeYyuIUqxy1al3Tqrh25Fz+KCInEQzJv7yb4W799+HKTnu4
NJViZ1UQchvGoRPsGAnVnbpaSMvTYopOmr42iQYFTQmQMUHYr5T1cft7+e2wJeJm6PB/aJ8xWj1a
ixnQg8dLmly6NI1HgMJVcB2iLKmo2PDaEZ1K27xZlhkzDZ3iJRC5t4wkV9lv28Rx5APpKFN5qSNo
GNOJ92mOB2c+jR7q5iOMZlmyvywTWWdByJVf2z9V34ojV0GqjZC7EU5iECeEVuxXpVjW1Pz/8Yxd
3AWudWmen9g8vuxFAIFMzeh5+L4B9lC9acBes6rQNGXnPOmrNbSoXD3h9AkVZrYUQJSBQ3/OxNCd
IVBMtxpyDC3btgMX4PtSVezTCo615lyHq/dR5rO413IeRDCUaUQacVyZNDgBqCPW15G/kO4Di5I9
71Ao45QO6zsvLpeqM4p+yJsdGhs1LzyN9QrPqg4LHpV7AmeoSGHoa8rB2FcxItI1xwcmYdv/vL3p
QFwDnxsV7yCiJYpvlF0Gf4zKCw1v6G2ZHFqK4JybEy7uTn/wpl252Rp2SURArDOALa9QtfBCoYop
DE2UG8oWs0Xak03R7+OaHXSrQzNvze1MrKdJmE3Ym2BCZfmPgGoAA5iSWn4Y9JZ5thTduHPwpyl/
43RAtY1iZwllCTGf9UxyjAHN+oOdaVe7MzXPi7GQUO3eNLM5HkXkI7zpqoggB+EGrYqNFTr7QXHO
JalkZe87rs1bMvNPVXnoKXwO3fOf3EHC0+kxMVskvEH2ST0Ok7OC+/nB7YNu5ChATciazRehPi06
GoAP0NYPldquPb/QlM65+Of5zha6sYuFsOYDfod57kQrVowGmjMLEel2yHmLciei/NkS2wvKWVXM
Y8uUbeogM5R7y86N/RMtrFz+FODBA+687O/EaPVIN4CMIB8ZQ184PoMqoW0spYBrwqCsbgiq/ZlH
QygYZmunkZvWxLHzlGeE0wP8/sZrNRbXhoA3EKFxXD0PkoffPWA1zj6MK+oGe4QSbijfA3x7jgEV
N7U2kdwzdda8NeFU7FicmW3lk/GpgFppzWMPV0yfKZzzztEFnneX+3Y6MgHJ/Xv0hVBUJMbIBF4w
Yo37sSFGK9EPPa9c6+JoqeImaeft7PvMQ7+mPB1dwjxt2U86ACd3AHzA6ueOehi2bu1sUGmAmecs
ls6Bipq8PPYEPuOwUibxfsV/m9NWgyNBXLCKE2Qza0RhYaqqhqnUts7Uphv2e3Vbm3X/FHdOzG02
wLrLaPrughCzBDKRYqKMzTAZ6TkiJGnvfNKL0Phlf7J3BOQhngPzmm5cKMGptRqMKc7AA7zMp0gL
wUpdgdkDZJNZg18O5qZ1XIAJF+cNKUALRU+S+zqjDR4eMCTk9ZOtorpXE+UYerGGyWsd3UnuGL2Z
y+MY9l+qtGGNPillBt7qDVFyvV4GJ+OmTE8Hnb59MYnwqUHmnndqdIueb2bDZIZp38GOfAlJC423
5A2SOTGXM3GvKk+bIEVkpsDwePMjeWKgp1D+KF4sE7L7szx133noQciOiVC/o+/3vPPe14MkX/r0
Nb6JG7o7zL8eSuku7X9SpsUFXrNURSSz/kSvmOzGIUpxn+YgTNKWCt/pp7WaHeueWMTfqWWnXbeD
IhCcZi88xe3tzhTEZgD6gOA4FxtM0WIPH//Vcw+RX72T6+b1Fz9XGgVrLbRdWQ3Jv9++FpKldmzQ
UmBihvLb4qv9uJUCWzfWPyH9LoGNAzDKRrtk2JvYHABsc+NIFKQDrKDOd3p5eGyDzdryp99GVcz9
POKfyIkvBeDkAhigmFUd5nJOwLKcqG0cs3rYBfHllVx0Lu9D4v2a0X7LTXK6f4/a8K+/5A2+AcWH
O2w7afDCm8AK1tDy4WXsV/WIQ1tpFOl3AJDMJm5LOhwdqbGHgbD61+Fzc3rxgnYxwM/8hLwhfKS7
dyA+siFZ16l16w9V1uazdSOOsmS/MK90/ob1UQ0nnlU9JjgjzXAIQoPdCv9jV1rQezYYjyyx0k0x
ApkCEyFZbD0MUw14P5y9qV9JqeU6bC3RSCpIsiIOgZEPaJPByn0aX7lN2sdIoBx4dENSTsLCFPUb
AZXp7xXoCVVJqBV9x8AGbLyh6vvlfwCWorran0MECXu3NJR2k71nMkqDQFExQtpq6RW9I/5gmgRP
CHsX2VvhNiNxSUMSeQnOHKzln7U/8bSy5hwxYDfC6ejtMT4QsCDzj+o2hgiiZ6MHLy2eCEOwUM/m
FMfBr/B86Afd80WTXTodC4UnVNkDa1fFhzWcQ6/GGtW06mli7xNQmC2+Te0uROeOWuxvbt9rKoVZ
9YEAPVoxEdqufDlxdQOlKTGc/P1Jnz7o9XDsnog1jg0F0sLk/pkkTpONGcFbKDXqcpuap00MTQag
S7lDF99KnlilL+pjZ3BHkvf61SVITNgpos6KAtXTfgxIfm1M2sEQe5bKZ1eOeC4L+Go9lUfn8zSR
j30V6FXCcOjMCwsa6BSmHDKaXjDXugjjFAIZ0jMhRDfRrvdUz7w8fhqGuhHGRM3T+QN0iMUI5DIR
iszYbrpnaNH6pLZCfrg/S0+6UB+15JKxhKre5JXI4r5jawWARHfT58EIWKvkC51AElkv/+jq6dOO
aK/edD4YWMmrOGDN4zuBMq4R6GJbzkBK6NbOsD+auvcMOCx+XMXqnwnk8Vurik7BamZ+wtfSmt0x
df2fVXOvmpMOPnofe2K1eZsWWls0R3wxZIQw1iMbqB5y4rMD/H2x+uayH/MY2BtXGNoPpkit34mI
aeMNoHhv8vRkZetzlvZxjPk84ZTlBvs1ROVu/BBTYHOm0IhvuGzoVzGTTq9bDPvw/BfRNdACvKLY
0A2EJoE1jk22GN3B2+w1Z66jAqKNiP+B7O/7V82h+imYGX3RfDGlA2fYozis/P/DJrYnyIDEoOv+
4zPbzWRBUPXAr501XSuUrbxF7Mbfu31BBdJuRxBJtMfSRfSbReHV9olpRti0v5ZId26Xk9GhOin3
fL7aLcUr8JtLcvOTzfzfe5iym3GsL1umElXXIC/wgb+arfyfK4Wd4No3sc/JR2KyvXmqHrNmDlPr
AQ1+wnaXQB+w9vmpe8WXs6Y7dUuXKS80MmxkewJY75TynM4k8DHea9QCl7e+PXJwzGdr21vMRkUP
4jT++tjua4S7xBd8D3ZXPyIVpj7hUrbkSwKMUPsV35laYt5pVSnvKwEigevksW0vasTxw1LWH95D
xLnFlZeq7M5eoaY5xlpwwMUGJcp8ups7qGCQ+hXucGC9KOy59IAG1RcnJHW0dhdYLT3WKghi/sQL
iL9uUAH1+pIy3KOW38G9i826gvl2+qbLR/68Yoxlxk5WmtVuV1aHyK0xj9aXRj8L5nAArpacas3y
dKORxKDL9Z1adBOvzvOYM5FQOpqJLNghM9VZH29o0ZE6aQ8UqKBKqMLin27h2V18Ucj23GmljVir
ZqC7fAXYTv/XJdvGEWjSlIJ0ao3ymgr9hFScV+6xCkrGGBH2OgYXP+vgiJVRcwakRNRBx+bNbHXb
dKgLpm49WsOK0+SnppggbmkJiP2N/31CxqeZ4qgmOuA5tky/mPtK/4QnF8Rq4eENuEJoInlo+zdc
bp3G+SyV7mxIZ7Ezg5kdWLdBqhrX2/7dEiojIACqIHQhO7QVZ8O9JHkGVIZLLD9Xa11+0rik+Wai
a+TQOl7jrl1YdYQvJC6vAN20WiVIcsnXjDefCiUSRUilCIvoWMWADu5swYRqSJEZpQzs9ADq2qu4
rjI/Ydfo9z3gLnHNivAZYolP4LnXsRdwkplMXnVbtTRbU7fvuizelOKcZlp3iZWScXUbGOJBABxH
FvY5jErEfADUQHbcr10TZ+wf8Sct62KmUaDH3KH+3rWAVz7rVQ4lXI05Isr1dJlWHf2uJBjx7hRF
K164Cdet7K6e6JhMxKx0A1hPR2uY2CaDvqGJ2nQ/Lkq2dBRtyd5fDjaEYgh3l0lMtcq65YhXpehq
831Eiq5LNL733XoQNqyZGnk86yap8f1Y8J8RWC/ie5r7/ZGxvfmuHRqBtjre1erMXA5y7L9RM8RW
LGYFsSvu0cbfpRhDz/teuYA3rUbDv2F8aS/udnwntFw0NFy47Hx6PSDFxwdvUaHFPR0HZCDCr5jy
QqMjwuC7NTRyXZZYhlpcS9c/w9LBs6QLQYnzPNFU8M1x8tnnaTtPXH5dzNkkOfG8Bwy1cfIvyrFS
hdn0dLt8Qy++i6maS61KjMZvc0QtLmD5vCpOkaxoWMCghW51tbCzljNuPuzdthW9O4oNMkz01U9H
BMaNZTtjUDhDmJh9f0LE8/KUop8Pt6Awv2UBnix5WYft5YHeI9dyB/s8wY99bxUae29XR0UOzp0p
OV8t0OCY+oIeRirQv2wQ/yrKYhQDeXy8WhG47D6Sub9jmpKvnjPRpDSg94BhPoBCTGmcDlS/mBRp
EbpV08mxjcxXb7XrpO5uYwq6Cm6eSsO4A8lN53evl/Aof41Zo6SZFu9ASqM+4pN+oaAp1oF/zB6+
nrbJeX5XrI5ncJRvkiZwnoherRgfhMc7YCCy4p1m+fHX4oAN9xljZwecmSLIM57vwj4MkoP3vHVg
aXpvlYA+RpznU+hEf8qku2lNx0euya9jEzJznncQFYlsfjeDrRJK++DKyWYvhcDA1+Op763mo2dc
LAMv3fakPnUv967k+C2SU2P1yLS/oirQUxUYCtp0TBS6kshO5pu7d57Us/GhVXQKxMGV9Ftw8FHg
stg8ywonqAL1vSq99OkqkaHIGWpIB2+KMjumc0nESdRkRkYtfR39F3gb8TL7tKfBdCqdgoYOpYGJ
UW82sPla3OhrHE2XCUYQO5OaGJHiBcsnwSAsRsEGjXiO4Rpa5jMVBN5cSBNDZmqbRwQboB7QUUO/
gKESqD/aGmv3axb45VmQawZMCx4FZCIJ+sIL/f4h+KswClkPMxKHdJCbJDHCB0yrU+tZbMD7BEWF
Bkab2VFsjlXiSGv3VQhfm29USeG6pUq6AQAaoVI64OKws8zd/cOM/z4tZzTN14rrszURkENp/dbz
75CZFvnrInWj4BJ7mrROUB9UEGuoexIIkYobYoYoGa7c5+ZVnUc/oxnPgrQuCmxGYcIJHST2fT+y
NLrUA2gQkPuWlBevPjCPb/vJbW1bv2YJJbvkMzcGHy9lB7mwaTzNBMSsyx0UIEr9yyF4xsWm55ku
JdfxJSY3oyG5WwJfUpcGvas4jYDlP4lhLUX1/NRYfliBV7nfshapukSlmpLde7jqxSKiwASyQgjP
xtK8pexB6rbSw46Qo25XdNyZVGz25XskQgi4ieD3sOzN1bqxpM+KSTbFLbeaNxCk83KYmwc2kg5J
MbpouWiJ+MJ0FM9wfwz11mFbDZsxDvAbK58wB0mvQYyBP/TRCUxOKzSmPSyCBxxGsu81S7WC682/
eqd1T6DWmHYOrla2Az9o3VHFwSFwjAExn7w+mk9unVwvPOldPcOikdT6UhqRcKtyw6pd1OrROAUi
cI9qzPuElPpDOgXG3ejE/+kVxV8yEDsa6tSfz4945Z18+01/8vxl3az435hm3UcaU+TzjyHuAeFd
jY3D1X3fyRJlrVZxetB3Lq2sZzA3TgHcxahJ/MEFTyP1Wb5W52nkTPGK1oGe2rYXbqjX3eiBslBz
Xcj4VqG9x28CuluX7bqY6/iiD58y6Yh7ZNdYIXrjN5UC+BV3q7LBgCr30dJ7pSD+ycXaWeQiZ4N9
PlAAVWMzQA7i6veti4cjklytxY3vaq/lokg6zAu1VsAi1V2rzf+N/fT2KTgPhW4HVHF7HDfiVe2M
KW88uUcELhHNEZekc3qE+L/zXrszP6sYM6rsNyMgLhJ1wydJ/xOZa9NVWAKI6BAblK0jwzqL8Pmk
L4Yb5PPpdJ7ONX3WHWXnub+GjrYElYSfERQofPtQ3f81LM6Z82p+OPgNMWcjctdpVIlCzv7bJGBN
u2pByFGhbu5HH9uUJQK0ebYasGQtwUJ3Hxrfbj4yMt0I7gSavrHKZ4xWCUA/2UFBYPigh3cJSMXg
UYdX60G7Sx8ZpiySuZCl02hiM8zaTBMJc1LZbT3XN+u+f7yAufAtHWTQzbVzqwzOm/d93u+zgurx
61JJa74oJJNvCsAUEIBzR7dxxJFb31uM3rH9eRx24yvlSRhafB+KFQL5BlUD4kkxDwv/v087YfGC
NQbhmzLkSXQTLGaODk/JBWYwy90OQUXIkJzmX+ijY3VRIe3KhMnQTg4Fxe5k1fsh2r6r128/zidE
+qdmRqg1vYnYi+awzgL6bb819Ggnn3w8OdK0SZsAbc07W/gegNQwgIEq21aftHSFqnaV5oZvhwTZ
WOMcpmnMnbxPh2MrB+IqSU2NAhV+ePL9UELVqLImF/z2oBfmJt3zkfjZPYvacw0WgTP+GFOlwqH9
or1cEt5xOpDnvqbhUi5bgSyFF8eJUibsOOcnBx7iRcorw5YwbnJyijqYNkgL8WY1DNgxCfHxR1d3
j+mam/eBO1RtY8An59aEg+G0ZBe1PT6aSA28OjomQyLL34+dU8uJA+vnmtGgJFZNJq9STH4fpeZS
9ZKpA/gRHmzBlu/1Gw+w3yhPDMpGmeiW2W9EYgCPoSsoMXfX3uKJadsy3dDfmIKqhHB0J+DiNrvW
XfZJ5xwVxAZnPP/r+QMoUyDTYvfYZnzAZXBWYjfNBqdc1T0x/TS04Z+Z1iD7ehw3YPff7Jl+qnbm
kZk1kr9DROOY/ONAlorDh1JeW46em6ZQjq9us7B6JJyL+u05i76Yv+YNHsX5AQJBecu1gaQ4g7B+
HtK6T2gQfg7rWFNlf26l+VToT0jtXV84YJsBuiFdFK0T73jr67lG6K59wkLXTvlDsbBQ5uqdj7BY
u2oGcqbOttOx98JLma+ZwGqMsmaGTW285FHlg+ONp0xVm7BBlv3rq+OHMBoedXfla7DvlFuh6MbY
RJRyxX7Mr0qI5Kdu4EmB/vNFucvWvz04h4jBC/nJGXo7BAs6DSV2T/DxAj53SXcuyYqDH6GdDwhX
CGfKCUJ1TU9uHkHfk0rYzxFCuGYD+8mz60xSqWblNN0fHRm0+2VTMaqujLt0/yiGX3XE0Co9ghue
nESds/2rdG4r+zppTc9TQ46yYX8XST+St/NwWiBRwXYVspEnvn85Gkf9XIjxit/S+6NxHPtoJ+9F
NF7UzX/PmnNSkwZSGmPa/uSxZZ5mqZVH9NXro56+TvSvJqa7rFuIt1hamARMOXQsv8jt0uqwtfzJ
/f1o5XY2GOeX/HkCj7FyiimlZw4EwP22I/IaoVDIPQebRX7kEAdiSraAe0v862Iddjw7SPWtTawe
btkl4OK1RsltRVLq9C7BMhJXrTMKVkLQUXCyBMjp4B2wrGQiLEesD0mG5siLMdOlxn4DV6VqiXNy
kXmK6yQqw0adbxYsC65kaP3wH7hryvBwQx/SR4yzYMV3DHPm9ZY9NlgEtslSYd4zatygoxecBNY2
blWp58culxFHE5K7IyfZ4rbHf2ybwDMtfj7pAu9OxiIWMpb0laRwTdIlg/46x1MDA43+54kMNm25
3HUaEbif+ruAbic2jxYc4Hcr9xNdfom8jkhZLKWH1WeMktDgC+k91kt+wx2ogXVMJPtQmzHtLMVV
95wghSQWNkXrSfr8MYUhi4zQHTRPvYYnJONdycAu8MJg53LL6uzoA6kxc7wtwsfN0oeEkLziCcDN
FqgZP8wUldz1e7ra+FBP4Al70FkU8lTusXT7jxAUUum8xy/tR5VqpLA/OItY75LGn/TbUO1sbC5i
RlMJuUyB0oVPw55dvo9K7JYIXoFzL6Ed5Y2RbBWjWnJlQEjSho3uQKcHVTmKmCCfkOk6aKqly7NZ
Me680QWVEH+ooEiuFSNegFY4yQ0yCPecYvkC43pSpmOnA3WagJPvISubpdxb4g79IXu8/61VPl5M
eaTbbXUuX+o/dHtpImJoyH/aWCN2xSZR7qF7JU/6V6Q3on8SU30a/AKzPrIwGTQJVF3PY+RO9Cxg
pVnaAQJZhyPdgkc54CsK2+rJNr2t41rRoHZNC7TEsvwi2yp9JS/t2grMCLJreWLDK8ei7HrimJag
9/GLtEaXiEzc7dtIWC9O4vnVRmTccGT8jos1nzknQaUz66PPmlSymXK5ACEYeJYywnz+U/NrqhZn
89Ya2ihRSLaxQRPszGbeYgyUyx3FtKUpd4q2FtqD2yrUcQWEtdkencA3vW5+9xN5uR8yH6Mo218r
ZnSqcZfNBVnd+bQULM8xTSbQILkXa3p0bQWsmLEutre2TIFd2z9AduPLlDA8taSh1R/TSEL4FoGC
Hco/mcwuSBZ8gOPaLnCAA+vmlOYbB1jjCPPF40iBYvHI/VOYdJg/bC0tcUKR0nxLdAjWZJK96YDm
plluZkKxCJ19mpbOYXHj+pPI6ApQStIftfEuV1+zGceSP3qXTi0IZZq40J50afe/Pc7MWEzB78W/
eWIC1XRYjrw7vZ2uvRpSyBJnzspSrau3LpLZi2eeUjYYgbVRQygKWQbGLe3c/jdnu9JmKIB2pL3q
TRHdBct2gyTOIRRtesr0/K/N8l3sVi5z39EhyK7i2yA6sTQEGbUSBb6XmkmNwASsOyju8HNs4p7F
tG6r5EJdwgrkXwh/1lSLzshKK8NZ1dGT+V5fnMwLmP+kyQgInQFCfaF2Ol6owJqntATBVSuHSkP2
0z/5xum71t2xRjyoq3PaO4REJ80bGDhGhFPoSx5Z4Me79q2+G5wBLBP131HxUiidgIkE6faR5/53
Xo2F0jYvIJHElsf17ZZd+IRAihrT/brR+SxIySgoT8jEGBIAfRvXy06yaYZMNJs3hrnu90fucxhm
KZ6OEyuo6AcKiUtiAXyl9WqiF3Uk8CuQHVocNeYy2UBWCT4qCNzbCbNqMhTBZyx07V3BLks8l/+9
32t7Zh/5fWmHTNctodF2cNZqttyTv02NUopgU6BgaI9OW80Uo0h/ESyFYXYCAJITN2FqFQww21SO
hzOJb5PBG4KTNDekKab6A0UMidW7jBfWn38CaiYTGMRQ10R5a6t6MN5Gak3ZKrhzKqP+BCh9+7i7
xdl7C6Mnd1OpRgpiB9PbQZy+LqaB+IUmjGDA2qEjeGC30JZexelgYq+pDnCvuheyg/Ec5i3hJwBX
KfboD278hxtxuA7DmMsm8ounbF9mBomhUYebBXitvn9kEkhUSrgF9/IPM589Ii68R7C9dSnQWVeR
5Afx6TI36kOdZ3Gz9feoAa9v2wuMeu1MMNKPyMy/L7NPFpz4a7HP9p7N6sEZGegmIX4e363fonoj
NT+2ZfrSkwA/Vp9WYD6loaYBFDcHncdT/XSLpbY0xW75Ux/RHOZrB9xyKgTNBTCW0wdJSkeuf7R5
gLbYWNpC84zh/RiwbAMy2GfewuMmNvHNblPuyvuHO+dPp0JYWUuNZCOYzEAXzSQWtMK6VPSft0Gm
hN07k9PQrMdh1F8PVsFaqgU0y5Mfr2RzHLyZhkBiFLfkg/nnm1JjTSG0P9T3IfSdC/sXfLKx2YGD
aX0zElmoT6IC546fx9yaRkZdBio3Qdu/lnvxoa/z7WH0ervCxX7RgocC1c9i8uvQCi9mNVC3Yzdv
5MuiQoZAUec0jPhAXsn+EnLkAtObNzs5b2a4AlxYbKvkyBFIlQDp4TnN7bw7E/KaOxBi+96NpnNI
jUxfqeazhlYXWa7kRkVNEEoUs0/cax7gHtWKWPRTrRw6ilb2YavPrp36Nx3+lOJwFyW15MNM8PJR
rJqfnE4OTIxRpNAp0iF9Lk7oQiF6z7EuKw2geNmCOYtsEGCNejdR0scgE7hxuA/pQVDZGiWz3axN
Y6aXhYvUK9IXhzpa8QoMs5oEMILNN7iqQjX4TSFHc4tsa7MhS7QWzgzvT2MW5VVyBMYqivoK7afM
kN3ugquNuawgAGvH2rj5WLjuZpHSUCxYF+BoS1yZ42xe2GrNAnDS3x7e/aiwR3cfXnAxGN7nWvLx
ixqTPJwFhCvLechMLQy3FQMLpykOUZRTWFC/wtJzEkmA75t/OGd2x+0xa0rFSK4B+RHn3mFnjY5y
n6xcJ6ja0OuwmsbDhF0PqTIjczgV6LnVCyMPutMFDjjRrMjW3DuI/iX+4cJQgpApYMixIPoCxocY
0igDKfnE5bGO/fchjwp5Tce9L5vq4YR4+c3b+6DF/OHJtxUt74B1SlljY8hxbKah0Tn28UAbbov2
gDfN7m3BnHPSDM9I1mVJ9ZjZHlcMAJoMKivY9qAZmOCqIDiIO882b2oj4Nuc12kybzsCA4qDj9ND
irzvsQT7AhXjZZwJBPh05aDLRpaSPEJCeOiwFC+2GYvgIF1wt5xQb3nTksBw2ySkN3hQJocFSmnd
qieUcfMGyOO8MZ/gSRsZt+KIipXzGHOeYFty74IVfQAr+YZMNlRyuo5zA65Gv0+IwILkJlAHOQjI
6sn5zdaVcPti1NlC1a9kwOWbCyyAw6rLksQK/+CuzlHGZap6nM6c9jBiA7rFo8U0REYalaZCHuzP
dFyis9CoaRSHFVF3Hy9krcwvPfKVg0wc2Qan9cwK2RYDFQOUd7tpMz6nUqAcyNFWEfWtrDZTLPit
PyRA2ntAuzV5b/w84XnH+XefiD8tgNspJMtFe5kocKDBPzFzf4SGMb5Y8zyrLIryC9wH59WVmV/O
g2oJfKauKaNlZm8Cgq37oYAZtQmA81E7yd93vdxSbwysX6oZsK0OAlRZesk7gVysgNwNboXWYnoV
hY+jJnEQ9FFxxkg72+s+k/1pvSD6iIyPammZqDhIoLqliV9dFLLOVsthO8GX1xgnSzapMRbOMwAQ
eg37dNHOZDuk1DvrzXqX89wgc8U19x/8L1sRA6z/thY3SVr7ZFxdkfndIMQujpxEx7s5NJehhIWY
xH5x6bLQjX4SBSJJQyiE0GofPslyisxn+c0XQxuo9slIbkSWpHJXhRs2NdZI3zJCGqltVtUMzPwS
vMsEL4xrsryMY6JdxxPVRetD3MJ4CIfAYmPaxOYQFAZscrPbDLgw8vWdJnVOPhK8DbY6CLd1x9ZH
w9AhrZuRXTw2zWbq11BbUnw67JCU/fndok+ovilQWKkjiVdEqVo0930wka4lwlNgAIwwEMS8HKdg
X8bJbY47VXtyHhiSIJYAvCDpMEpjiUTWBtvXO1qHxRz1XTHN3fLIj+u8TUAO7F4HrxV2cJMVhKI2
RVsLx9S8Fus4hzTBtGdgfDI+55Zj5HOcN/h4nPCgu/ciWgxR8UqB5loNZJaRW0t9l8Ew1ytzB8mX
SfhPAJPlnAJuSeMkkATdN3RSlXSqw7K0FIuA6tDJUMi76nDGxdaqaPnvmfcVjuPMJgu2gzRYzBm4
MRJbw0+O+C0J70JzS0JgRHNYYejC7e1CIx2fvW5hicdBHSbfO1pOMYbL+FmuKItdInDhn+CYv5Ti
r67E8muwtzcQtAxqrdbyhglucXPzQZeew7IlH1CZ3c/M2+4Qudg/hqibl3ZStT3Y0M6HEDTt7g1/
XXprhzjA1mXR3rX/yj8kPhvU1E1KPwPkbGQd8ToTT28bo2L2F7bzG1/Jz1MNDtYrQjM9vADhu666
NliuuAb5b8DgrzTwGpFVuTGRcwh6qeEAxm7Bevr6208+ASBlxdl9jA5WNz7Smax1Y/OOnDpfcN4G
5to/EmPkRdd9e8aqAIS1kmudKE3bUhDOLlHyr7dekPR4W8KlxHR6+9fkJPrYtKAs+uqg13Oa54z5
5tG65khSZC6COxE4imWqv1jxGIabjV/tmIOgt3LbCk33nZUh32tZQFBsgSC257KNI3c85LF/qdpv
lV+D0dQeEMDuANJWYlmh4WCNPmLRrl9uE7tQCgu+Kpedc8JCEqMO7lTmCntvYMhAKrcYoFr9wSqi
iO75IEKXWqLyYfi9ckCe0DIL/E8Kbgsk/LIX7XszRk3xgyt5hDWhq9sIFC8Z6mrmRgDvhVfmINWw
IZmJHi7WM6P4vYvj/h+Se3Jqqpdk72h89EshDdpUY+cubfSTYwN9fj7/9Q9sSZwL0+PX+fneVSKV
pqni4SGoGyqAonxHRQsHp9H7hvt/ZocAyqkH0E5tL32bXpsZYUZ/36Zq1iGQSk8XNlJDkRQ9UZL/
+Li7A9JZ6iBtl56vEH5HHPdGsw5KkyHTEwmsHgtqypjwaJ5bQlk3eX2MbKiGwVa5IfeRH3EM5Qi9
8r+EWeH6sXvgXZiaNZt8IK+8brTtv9Y9NHGzmvNTbor9YSpqfMglsXVZu1Pcc6ynpfgtT3RNtFh/
ALG5GjcGMUZtTIoojDIuyUoK2+V9hoIslBLAP68PIgmCqdcel3AFO1oD0ij9SrNh74dte+ytj6P0
njCb8QhJomRYeymUqkPq6KrqsoGUQJa73iML6k9T46NSMOABIGI9u68/FmY5drL3DNdziYdj7LJy
+RmADqOSPc05nGa3gkTLUE62ZPs64fZIVQ4s7CK24zd+Sd08O1jA67seI/hCOeEdVQluWQbdl5kR
Dv87IYy1xPh6AzUYQudBGXPXyjTuYHoHINwlMGXhJiGeY7QaJ68Ppm0KmVp3MjC2bKTspbwrPjRr
Xnp2gQbSfjZAW/RxP+wgSj24rd60GZyxcr2pFfHlH43eaCKjwxa81p/fsPlbvpPG2bJYxSsfAWcV
3XVJyK7INQUheFh+RpxD37laPMAcehV27/9Ks3LfdN4B3O9QsqSqn1QdaOYVxpIplV68zxD8ahfH
EgbwPI12s//kZoQT1ypzJuOEDMcHJoT8JBCJpc2hkC5BNhNc9zHSzFfsFvuwDIa+6QEuvE/5hkzs
1IocrzP1EIqpHFmVuPQ2h8RJicr+fIPEoTheRRHqdWwZiTTm6bf7nU2M0xKLN60uM+MO132cYzVC
DMoOHMU7cFIHNcN+Ue+aVwWJr/+46PgLjz4QE+53AOtAkgOCwaQDZkTjcmTXam1FddMyxZy6WpTL
dupYVBy3DZOLLb/ViUzm54fEluQT62RhUSHZNWGzaFZmlMzbOO5jAo4KRu0n2LdzAyDd2mGPNXuO
COu7059Vqv7JcuV8wyX6Nvl5yHylUV1awbMTOPKGtfEGQnLVek5ion8NMVsUQloLhEtoJOGoKwQX
cCU9dPhXXNaxKFQCk/hvC+0XvMliRK6Cd1F6kTIr+87vQWglN0KfPSf4hKK2UqMlay+GRdjYdBa3
8xerF4KXYwqNvccG3TnGxkBajVLF69qm+aJ7cC/weEsJwGMrrBMdJXw4YtviTRcwW35qajBWyY1i
kl67hgcwbxp7mkBxr9LWQOrj2xYSO3zSizELeD1eREedxlixhTVBEMVkyloVMxIQZVUZfKMfh6Bu
2gryaePQ0MskK76EsDh1+X2kmAsEcfLAfoRUc4CVWeG7AdqynTpL6k9M2LfXMj4Q+1ckd3JCToTJ
iPTuWrj3dWEthVZE6emHmLFZtFvY4lnkYlDxagbyHt7AVXHUbEK/Ky027yHt5UUt+feUlNwTvv6a
TiQzmpfvseDdffIO+nUJW8M9/dAPiPE/p/pdJdE3c3uJvu+NU7zRISFfvEZHRqBLmBDupm5iVwB/
iN+nYFIMLfXxuhQnEeasp+PWWcC6EwN6lX77+1q4pdj5Sgby2frGV9bVNUAWXAK0gmXb3dwXlJVp
0jdDFLU2iUggqoAWVCUprJpHLpxy5O6D7fRFNZK93XL5pWyShBC8D7DvzDUjW6wN
`protect end_protected
