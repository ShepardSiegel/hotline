`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hq8dqh/p1Mf5V8kov9bDhCgUH7MaFqeSeFKYoGsrgXcrCYiYbGigfjCZer9YQzfBZ4bYouEPQnJ/
stDr8WitgA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dI9tZWNFLe6oSMq1UkJGJJOQm9gAprMtca6JwlmelhEXgeXwFBbTbeNtT5GcxzLj34DtctB8Fn2B
eupoxTvK+d/qbGo05WMVaqbt6J4ZgnFRhI0FF/E+mCL6HPao5pgZMCN68/voFBxwb5NRdbsscFtt
gfg3dQXrS73l1pRJCxo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tQ+G2xsm2M7+pgOpfiIlksWy+/pGN7Iky7cbkCW9SoDRG+cEJm3oahvfC+vdP2NlMUF7A9uoVpnJ
OtXkf6Xzs4d7CM4jqnHGKhZjckRRcSHUDHTYgP6ieDgxTzRw6FPQMRwGmuE24qEqq7mJvwCQX8xF
LbosAn1aZDBBjVsBWbwsimjU7vJiNDclgVCUtzDlYfzJ6hAEnXlFFMrCnN8RZ+7PXsvQ+0TWbgRj
+YRVKreV4xAJqXi3HqC5ipAFUFALtQPOGy8KHDtOunetyEISJ0iNp4bTv37N2ADDoQuhoQqNQ6r7
qYNf4Ph45k9ALccWLKl38SnF689Dn69yHKY6IQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ddjTQptBd0zk/T6frd9ROCsL1LTdAsoMl0RoUmZxfzkn6A9GAWJZZ8oUtLn6pFzruja1oOI+ehrc
h0K7kXMeE0YNihUfkMhydoyXJFRwpz94IXfbHA68vny7kygtFuho3vlH9bT3bXl/gpdGH0A9OJYJ
oDWrxR4TwGFC2ekThXw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UZmNWyrTYWDMELlFiOvHIHTK0kTGBFVT1iti1LO1iEIVWx60LCLB+xMDWkh/eqk5uh8/t08uybEv
BiBS+suIoO1tfYgaTT9pvPT2IByWNk9cLck8M2lbGmzJ/Tf8jksClbtSHg4itL0kW0A8DtarJ25p
D34zGa7/fngpGcaQNmKD6gt3ofrl/d/OUOFFDMIY8dm43eZpgZ8vvXrLJDXTVW0CxCL9cBJS00F6
YEOEc86NHZHb7782Y8IQXqpncEnXF3uqPwhF/11kMGz4xUXjf2tvJb5QDl2DoEQJ8wT875dpX2CT
tVrXCXyfOVDMvw/+4ER7r0Yyw4ES4WCuO9d0fA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 58560)
`protect data_block
c74Lq4wFls8hbeKlaCmywO8fJxtoJDsO/kPq/ciUsaHCl6BMt83/p+KRJXHfo+FD3hTaKUAszQy0
xeqbwJU6ZtYoiH0agKjk0w8Jn1oNCfujrJv2N1Yvs2wsyfkRpqVkridb8otXjOIQDLsqmmthdYgU
KhMK7gIXFpqNWp9ln/knJKwKEcK+pRVtaTgUtJ9fIlTfHz5OhJlml2tKoatKGCTdAcrOgoZLaWp5
MB1knNb5mdP3kKcSz7NwDetQH3Vf5eEUZHL6smREw0y1haPH0Ao1g/P5W5JAWExuD4BE/+MJv4VS
y/qa1qxQuOqVOROstPznVS7EDbpogC1sVhE3nBtHETSKyZnQNt62ciNq6ofMALYQNfO4fNNuvRC2
KVRdqYBwfa9OqJzXphNPFVEWBEprtqdFG1zJkqdVg/qCOy29GQVqhhtecJj7bs7a9XF1juvEFDh9
6Df7Te7a2gGZTRWMy9qGX/pvarCZXvDLVXU1xNgaJ4dzrusSr3k+yLB8M2Y1QOL3UqI2YZxUrMLR
w0HtvZ2nt6ad5WHfOjeMWQ6oBd/DQQumV/wgKSG1Q6Kiuucy2mIYQXMc/onjLZU3mSsfyHlwzJUU
BoT6Awr3Zrq/skgLuBEvvwXGkNOLjZAvThONwEnr7s8SZ8vx9wMla/ac8BvXZ8zisWMqhVUNGZZj
SMwPJEwX1iyteomnE/9cAE8bIlM1F4enHyDNWzMDsFSJUd0iPXLbXqQfcs90a4PIz3wnCoqWsXBZ
rjzUMprfXSuKL9wx5WDoRfG9OkZ7q8pP1cNzGYUMd8j1Oq2niEPgfctL4WP3xkbdtaIgcyzJQwL+
doV/C5ugG8i6zJQncHW6aZXouCFXclC4uSZIEKYDzbrx4GX7NUn2er4/zMmVtra1X1gWV79AZF92
9mb9tq+bUxUCUBGNxWMN4sRPX3mapQ+SHklnqmpvi/zYi6Wa8OJgljVxCHpMDpwvJPfvbPix0H/R
ILUYC63PzPf1giiAe4uA2g31CsSiux9m/Hblz2JdrtN5xkDLicmdLpQ8Mv/ydCp3f+SpgPL4BoQw
ZPWCHxoE05RcV005IIOa2QvTcxsuf1Oank1ywoIX7XAVzQKfeoHQj0KNEugQvBTx7XHfMgfnZe8a
zUh7hMHpyOUns1GxKEh6SiK3sonpej5LS/HGBqOPKsZSCz6bU2NrkYyMFkp5VJPTgeWb/iouEF0A
h9pSbB4hR/SVBsNOUueOQczd8V6sNgC3PccnwR4R9xZAISvcY7LpZMGfn4zuGzLB8HiUbmGPG3xE
idpEVHKfxhu1n4S63yQbR9pwUVoTpHYHrXqnsngqemHaDoYcO+53WkUxyuxH7Tm1e6VP0n5ewc+5
jIH7C7KhSyM6fnxFJgkAUKimnaL5BxE2xyrld9ZYPrG6mE+KA3uTkMt2fqtXawrzJF/3qYiKVnaU
sf0Az+S7xcCFtSKJdk9BKOUqsoZRNAU3JVXRw3T9gYlR7aKLNjEG9dqhm8vlkNvP3eBcyuXkHkdq
FkG1Mv8IS85zShgcgZ250yG912+s7iT/3vxiaIJm09eQURmcFmYa7OotiSGfTVj68v7VlohQ5zmp
CUF+PC0QjVQc8dlTnHbTrA8vnChhg9zH3TGZoA7q+EzZKaYLEZYkTSsNhK/rKYn056sxucUpgoyG
/P8vqnZjrcoQYw83XQ8azT2sXr5aEI9sqCPlwEY93kJ80G4sQFdseMM/d6sHYbS8xLEEAsFRcuOc
EQBPed6VJa6Cdl7h654SqH4zLtgyxLMzAjDJiO//+haXORqECDDoSjVg4WYo9ZU3XQLyCZZNvZ6w
mEmU/5Hc6CyvUCCEplAkF4hAZfmv+bNU74hN/CMuYRsselceQqe8w83HpWt1/w/UKpp+tEx1GiL+
G9+QpgThdI6gfS3xGapqbAvSLIG32Zy4pfTt2O1RsIK+uzjkbsfxe2MywKIe1l/VLhhRiZ//djZw
orQyxTG7mk1FXhrkFf6S8dSmO0dKpC4T9eSSS1AC6cXAe1t8p/qj4JcamQXwEBCdFjv6onkB3XwW
B5Mo1MyV87JQm8Z1lmd17NRC+S4I5ALK93MbueCZEaYJkeNmNjAM3aoHzF4iuuQBaHew+tCzAyEX
va5L4jAZdRjcbdJGcxlW/P9P2zxSpF2QCX7CRw/gQnn4oGb3fS0vkpS6nbAwMM9Hek+l9vICdJdU
N30nM8ytdtEPGugG9HUFc1KIJ38NpsM53FRuqu0Wi98H0hxF4Bkclmd49js2UtkLitlVoXdBiZBx
5r15CAvMu4DZUXsPjuTySB92UfhlPxlQRyVnMym9NJRqF14Ry3js3xunh0QoX4FnNmeS1MJgnw8/
MnuOY+xxnqh0RxmZO1lKtS+q+kMffBsHTW2dxo/5JAdKzdcUZ2eG9mPU20nQWQtbdpFSoLE9Zoxq
re6xi2xYsh/PMMQVSbn6DoBN03RIMOmAePvclluWCOp6JM/UFaywNOhri0Ity8RHow5Pru/aTbUv
EHFIm6CyyMoOgfNkJJj9jm1TfnYZyf1Hr37M4vjTkiL+f028cAo7o5JL8bcajSkhXpVieS6LvN5F
3Q/dXYzQEDyEZ2jrwvWWTmL7XLfBIwg01ZisMmn0T5DnQzF5Iap41jS+CqF4HWp1ff15qm7/ATD1
OmPLWTc4XCzrIWGD1bULcrHleL55lb0Qy70WsGqdJdcruf1fWL4+UxVMAJTk98lO3q/M0TUJLJ2q
dJY2a0Im4xxS23RwY0F1cPpCwAZrIh26w95AiQDeXglr2hsTV3VOD+ZenAVcBALmRmJXH8rYX/LH
wu9nC4nk96WfAxspOZVTa9q5fD5e+Ec6kydmji/8TPBvH1k0jZR7wm8LZ3Ixrp1AiCPSuXy62E3M
BmNiHy6lAgA10G4VYgZ21UVZLVytu6c3s5ndHw9g78e/KMB5Jn9OkZJzOcb3a7gKIAxON8Q/snAb
P7HpXMf7Nz6dsdbdlO5EQSl1Z8vXKzII9pQQbG7vSB1yHqiRvifT3PZTL3jXQ7P/p8jvORyGiWGK
wzdYGNO8uGqRMOmzUgjI2TXTBKk1lbwSVY6062Bm8cYjGD1PJQx+6KfxCgnxIT5AwM8mCmy77S/C
aTtNRpwigc87WzFyDXJwqERpSiYdyWL5QzNHqpwZyXY646gdzhWh59vev3EQV6Mncf0LgSwCRXis
6SNrVVBFrPqR3c+as7cfkX/M2ubCZhkA4FKy8846Evr7/ihRCW6WBrABHIhl9soYHpaUwGkZjvqr
Npu/niVxmeQEBeU0J1NmxTPthP/BANow8lUSocXgubnLhZAdXxUBtnqwUXVT2y3sOP6dbqDrbh0+
QncCPLI7+qq+D5bd6K3YQEIbRvJovRZZzDeLNSrNTZZ/c1Tc5XObJhFJqSkdArcgc0oRJIFJU+X8
01MZe5TH7hzzQoZzE4Gb0jSo9vZ8pckcfsOYZcAsPmDjrBifgsc0EpMlcwn8NyvY45Ii4s4W/BFh
wwTXC9tOwmQuYXDeOjocC9jMq/2SYiI9trSORiSHQhuNyD1Rc7/PmmnKaX5lAbpYfDL/vVCpcDAC
DZ9tnPIvmk39grAOwat+fJganVWK1DY8VC4MITV05QnPaUX4gy/KL1FnwbB3uIG1Ho770/k61wi2
1RQMPBt5Bhr0KbjSggiLicEc+tyKhANU4o/+X3gmWuRfw08n7IA+wXWcvfmOtR/nzsoPQ0hzfL9X
SwPjI3+/0jm2quMTV7RqWEU8gkXs8RbSnXbsDIsyYkz1quZb3P0clU+8uXaiWSn9aHoRs0jw3Boi
ZtaN+7k5olNYZ2fcMUzB11eZSiWqIZEXlJGO+Qmzfz7T/+21g+EeWuJdH11NfuxKzTHMCJqvLMP4
sfj5+gz9ejtHLAR7bo6xiExnSUl93nkZExnw+LK3q1+WyjBV4HR5GOqJmFXyaPUv8OogyE+uDKsF
f0HwpNz+dr176wAYmfQ3vaBWb4PZstOdN70j6kYND471F6DMhO4km90PG597l+GAhwe2qH0WeHcI
q/chSxdSsvf0Ke4Vqbna9JqD7pVRwo56j5lHCwn2gQHEi/mZngPyhaPruN5LejAx1zfEVVYWn6Gt
U/fLWyjRmeI06E3o+3sjVEclNvxANNxpIlwi7Mk7Wm1hDxm6M8wom6VtFFUN0aI17SR2IQLANEHo
02w/Pk+0IjiwKNP5nEhjoO59dfglVHCAnU4I2/d/rd1Bl0H4oyjvzoGtVQ9lnl8Kvnh24AaIBi4Y
Zquru9OMVyrrjUeOtq6cbptFvQXYhQ/+V350xXlkRuW3OcKbiN6VaiFeEcshCtuwhqySxpJ5opyF
eyVrUusbMadikET+81LNfyjWswQqrLls8jcVqInDZ9d56i2AmQir6TXZsCAjnJbjzR9wFXQqnPqY
Tzcl27myGm1azNDHX5dzbQuqX/TUKMu4ZeSMnLCz3tWfKbG5Zd0OaK2ptnl5B4zGecsxdX7ABURU
q/FBxCHcBaYcOLkWKFQyZG4MDVoQMoEva5lo1QSS1ZaQbZ1Vx34yOiL9ZP4aJc7Kj4YpHAFUIw4R
+D82F+E1YpIOpbmoF+YTqlMm7wshJKNNfMwIefTqNqb/WjETiJTnNB767vuIiLBNAnLteZXWju8w
rN43dj3eqDlPM6ijGL6XiSxHthxT21riX4KpeSmthT9rfZ1KqXO1nFmfS8VJQdSlRKlk0Zmw3hMc
cf/EoFOYvV87pD0FpfPi+Gg1hLgxLAPn1pR6JcXz1FH9bMBWv6jY+xREceE14N85ZjIjAxTmCA21
JjRt5F+7W8fUdxE8RwZPksWc+IijNGdI/jh0ggr3ZsKSjV5v0DP5fErmoSCyhMVl+8UphUXkXWRo
OVrYvh08/X5/mZRj8Mtz9AcHzL1lYkVYYaTHXSDoth7Us1brvqnLLnedqD0fovCaHSG8lQWPDyMp
bPFiA76hm6zujwbacHJOYKg6w7aDve3kMWUafBNmpmEJU3kFrecPrqz72m7CA/SxcCRGAxoYWr+D
5Bttt10VGLzlU4UYkj2xhfKoSzUsTcrttIk+1a370NFY8EfdI4IInEPpC7/3zKGu8KEMwMO1Q8D3
Y14aPN/6e4kKiFFO8JgNgiBTp1t9+QYqB7uEyF1SgK5fQh385JdYSWv9fyx2c9CVvPfn1vTNHzQL
xbxY32NpFcbbDZ3qyGQUMXsR4k2MUJYdr5znXnbvXefWZMpP6qM08xmtVQY5d1m0FzVjTwVsvYgB
qgMeJbX4+dO9PK3tQTHdX9j/hMrMokuWdDvYUxYzzoECzA1A6HqIsc9S3OpFtb7oRkgWgGOp+iZa
/GoXlCZXGa2UtfAktefk93vQhSuxoDkfUIb07o6Fm45t47/1dsd9yQ6kzLot2/tqvH/4QrK5fdu3
1AZjxjwCSATdFEKNqUmsnnzxFikHWZthDGYKWwbYbQSH1BCUVVPZHgUTSYIS53MIoMUAw6TFX0rM
SN9iIeNlJd2F036VW/D+V4Fp+fGrLSzzbqI22sbVI7Zz1d3YneRY+m8qVErjWX+soz6A3emzf1Lm
T66Z5BPqhtSwlomkI6T/ycReBYGlSEzuK3hyEHbjcK7P8JGZ3oJ/VPkhjFHxmWC0VQOSExTjgLPi
VtdAPO0rf3vVDJ8AIVUgtc1PFDnpwxcYQ1l2OtUuB3RDf/KbDCFqY3t8dA4iEBTqGANoD/5/Vygs
wE8z29QIfEtvhsLmlAr8+jqZ00erCyUsmMq08k2EHnTwxeQiscCGAoxxYsQe/uZYZo4eCfGP1RL6
wn7KwfjynutBAURxP/ouflpvItrWi1Z9kbTcm6sXx8yweWgwetlYon0+CKD/aY40WxOHBOMEkosz
/TybT1BUs5pUKN7Se35v897+wpOEd+TtXxYf5RiJNa7Mer7iT3O7+nF/SMk2nA6+FXsvpslcaE+f
fp1W/pxFZX8XHEzrGY9bo7/GpfZEOEiexXlCmqDrAQBjjbG8UsKi194RfXpMcxuOnj/yHldiM/jd
IJSaOSVIf+5NHRhqFov8pyg5ohbolS6sGsitnVQL2Ig3dFD40/IBTdDiVYBZiY6CYabwqhoudemX
o8SVuP9J8lEMfP9MyEo43S9srUY7Ez8y4bTgOy5SyovHzTZIGsGIyr6EmBlEumYNO1T0M2SSmGmH
bz4tX0VBZsmhhw87WTTwMe6C/t89BFJFRr7owc+YfHK0+Y6al7OkdZFfkG/yEQBYrDZKWACN0wZm
Ca2MsLmXFuCQH8et9swFpOXVo0q41/kfoESU2lndEm8F10GIhzBx4pKPr9dN/NNM4cf1aea3LKb8
PlbvFadJeIKrUdzo39D7qsi2gj4VKLkOzzRJ6s0Hkb54/tAoauDMDPM/DbQrekGf5TFdmYHx4dP8
G1OwC8OKebo1Tm21vx4XcleW4QAgDCUIyHdT2tm7Tpg/UUCg3BSzbD9kMnFEwQQcnM+l9S87Zsyi
/MTOWJcz+J5ROCGjcUG7bx2xDZ2+xhNS6NCym2Drns+dJJdEwe/fH0Ij65zBWLm4z3wtjQA/j/rX
L4yeXYKAfqCCy6A1R/7NHLWx8FfxNw0ZP9L8tRJN/jG04/p2iLuSDsPzbc7QjNvhu4pmiz6dSNHs
O5XisagR17g9nIiiY9bGrKvTzfkLSOxGJsIo8itkysp5Rop95mIK4ah9IPgj9Zk/XA69xsnt3Lho
TZ4e8eO8L6Awp3+zoGA+zJ8scoTmLODX1y8uwxhDxs7kPd5nU5rH3Q7fHJAMtZuqfDXdjJAFkgSO
E8rIgodo/tNDBgxnNfdR5YHYrYVWcrOq/ksprED3Naww1HzI61ioAejtruZfzaJosPUpCnlzGKQL
Sb967nhLzZNxkCgzmrMuudwmk/dlhv5+OyUXM+wVeZRU4ozteJfpl00GWkAQ2aQZ5X2CNY7eh1tb
RlMK6LLhcQ1P6a69csUm/bhU1djbRBJvhW6fN4byxSfBeHN6RA/t7EdUx/9uOUGKVZ8Ag0s1uqyQ
8PidVkHpKuGbqhnnClU8Ehl28LXNkxSCoVKqJ60b2eKcqxKa+JH/OoV9mxy8VO5R0anOXaRF4mbB
4TYDPNUQ4Gsm6rTe36G7dMFbKb2LJBeMRxicHjO+aApp5MgQESGOdn4mXZbgGrlyxdwVirk89i9K
l5R/RW6mWe7Dix5/vtIovPpNnq44TLWmuOnGCQeoGEmTVG/uHI+Pr8zqPWqBlp/Tx8yhrkhBm/rP
tVHIibXtSRYRjqEPPBDTsuAp7YjidVKqgN5JGOlKsdTj7ELm2Xfz4X+4UjVjLZ64fZ88+NKfpv0s
dNjCbR+MH+C8pkbaNuLgB9K0wUaFQivQiGQ/0AGJNUBWKSjH4Wb05VIGlT0TQHWCejA5I3iXT3yx
P45fzvDFNmWLUh6pQc8UBzB4w5Yy8yHm8oB/RjHxwYYFcwTjW5/R0T2fm5XtQt8cck+qye8XGQi7
1v9QXHhR99o1v+g5sSC1BWna3InlgNgmN7DLf/f7VokulAVCeR5g0Y9br6Xxju7MF2IdZN7/Cmu4
0hBmRlGqiUoLSeZxXzK+LGrbVhMlRNM2YTFK8wqsFERozucoe8LqgoBC2Bo28/7z8kjeNLGDgAB6
79wBU0I4RM2nwipUPyO1/UbtyTomI/7vk/edQVFFuwcn1gAJwr3WSiUJnkB5UNgxoxkIDr9UnclD
b2EC7k4WKTG0aLiBnBR2owbAw/7zVHUsc+AUdhEOv7XPCptfB1MqPyko8a8ehSn6cono7mUhYBaO
B5RZLvpR7iFQNhBmqeJFY/kJnqpjwXKky+thJIK6/3k9JWztjR2sw8cA2gdrxYmqV1M+L9IJXyj+
Ys3/I3GuCUCl+/PG6hxPgWGM7Gz4rv2Kx1MuT3bOa1rVQxJOLSIq6SQoS8Xo+A4ilOge5GyxMpzg
BQBuoFM7plRbaZjaOnWQ+iON18Df9uCk6xjOeh5et2vRGLVSvPCT8Ackc6ufcUeeRrwsOuZymglG
7HGUyj5vSUkrCDm5+ttaw7UMq8aOLqLg6MnlWNDm/RoawB/R95x+KCgFlXvBC+Rc4nM6ExnPw3GC
xL4fHUleg/kVlE2i2Cfq3CKFwBUxiefmpeXS2lipmC1szJRn75/FPEJXc9b+8NGiRjlsIq7RXegG
UojfBoMu7iQlUeTIanTAFdAfaQbUgfXWxif46YXH5nQTou6/ayxM5ZdsTbd9NAB/VXg5YxrRH7DO
Ak7XYwDGs5+PtNHkypLxx0rGpFNrWW+VhARQbf3+1RpYN4/lo/OdWLouqe2xSBIzVoEDnA9uqplu
pyS9y0E8TqKpfQD62mOuVYqZ2H2PZ88FaaSSNyZV8xPBtW0FI/RtNThzIuTPYlyAIuFxP6PKp2XQ
o+5f3R+1+lrqG9Ksa0jMxHygC0YKh5tb158iMTycPD4Lww3DUxsvEa/IeQ8tT2KhgpzTIUdlQrYk
TY5wAsvILFCD0nYY7o4bDqaoVF1K7JRdAtNrcZ5nr0vPVCxWark5NqtVqGgmDAepGgq3rDkeCO1D
wAa+lMz9lXLZ8Kc7OHEvm5MhEgpbL1BvY2CD4urjyRn2clz61kB4uPcg1Byj4enIVFzap9fvrYeY
SNWP2hEBqGLEL1y0FqtDAUuQ/AcvA2r8GUdy9vNufNo8IjkVkVKzPa7wf1AuxQID7S24X+S6FvYp
mo6R4LGpgi7CMP8QjqQHURMgz7J3Cj0cPBKHQSimo/cLf5N1nsoH4ZLQwRnr+BZEGZczKvZcCx8j
72lTEtz1mzayr5qzan2RzwIJ2eGHLgSAnnXEvYzzD55WVYCDTL857aLi99eh++pIvhw3mrchwwUt
Ox9a/QsBU7o63ULIdhPzCxLewpayLbssHy1sCEEV7VDFyY0wnsCPvL4Nc0q9nPUFUJO6WPrhUvpF
7mx+WYEoPLF+qCAkK2Uoxl0PuaerKw+db4CujbQLSVG8819Cg/TTvt7c23lgpDS3jT3fv6Uh+z9E
1ejCbk933QNBgvQ8jX4voTU6GhnzxHtuNVw5Pc8GRxVDVpYQENJjFU4H/iNVNCxCptgpw1ILFDyZ
PGY4vU9fcbym9WG4Ct6AYKEvhjnmRoC/kP7dSgRO95n4w6oYNwRW9kwwXzG2fYWhbCXVEE+EJx4s
CDcHumc7JN9jvKeeTgYT4wpyeUyDYtQfw3T5QTCVavYBKGgQiUp+rBJ9VT9ONta4wBoBXKmrZAOU
7kYHi7QbuTE6yuA/1X5WDM+Upk+67Q+hQEj8f9RyxiipuftwsQFj8TTEkRkPIMSSVfpYk+vhu+i7
8889SCuKY2RlX8kdyMiQaQQ/OomEXZnxPV4Egu8uwYR5FAarObhSH/mY01Ct55wXJefFwdvK2Gmz
/SjoUm1QAMACUn6hmVPamhvfYCmYD5PUzbqMgIQZNhzg8+kXPJJ1edeA1S2CiuoKYh6jGTj/t2Dg
hD8prHxN8NPbuhanzn5Tl6M7BvYhyZZrrtPthOJI7oINKngbTuDDY7N/Tg/xG2KqOGPbCdoT4Q5r
nPWe+FI5bv/f7yWFK5AG7NXRIBjpK03KH98xJb2U6q6zs/wLSsRFwxMcDYKgX8NuPe+yUeJRh8LQ
OrXUKw6AahxtKdSALBN9YaeM7dyHm0u+GdUEZ0sR8SvbyBm/+UsNJ1sqBwwEwtC3CD7EAJZblmvD
l3DcmgH36uhr4nIuFX5/qwpLUNCpheA0CMiXFW3jcOCVfAHzOdHBv4ksbPggZFNkVUT9ghPpBPDm
9oGp3HE/dKonROgA2CES718jU8Czk7HZcACvfSX8x8VRYg9C4hA9UpO4jaa6yAAB+qkJY0KRMnub
1P1rnXkyFNXre3BLmLzp2BRdylasADSplSIj4iC3lgFwtdvau6r1R0/pnk43lkayRjljlgd6FWl2
5dRxl+ctUh+HQT723KcgoH1uBedCZLIboMWdrsTaZHy8ALhH0lqOJUIcKCGhtvYsGlKFfKKJgQEc
TsZ2tzqGo32qGV2opQ5bmhlXymFwqccxZoZ023uTee6jtLK17HCm/Hi13em8LCjvgeGXkF8yik8O
XW5X1j3fboC76mlFCfG4sJT+6InzAf7HYZf6Mpj97gwTXxrvTLKlf0SednVjtYtcioIeQoMTQzWP
SKhBnPsAodTE0M31km/LmILiRoRAX4Tic18gGvV5UktW/lNoIqowPb81kCT7eKuAVrkLuc2Ip6Q9
5t10CjyhTFihl5A0SBrVFYG5zY9I89VAwMw4ZnA6r9ekAmZHkGHw8sZQWgsH6uVPv4CANMbNEr3b
tBeKGloZYzcSwedXTBE1oAcvL4knrPV7vAMP02jvSKGjgDWAc2o6zBj3Jlvf3qI81jLikJikEqza
bzVrqXmQxOPWuSfYRvGF27UU0sEWK7UMQRZQFU8nLRCJvqK33nNaJyldAm2zWJ0X4nbpBgIr1Lgx
JW0Y9jiKdLTuFjfhKVrPXSxkKidxxG9uI7N4+W0IuENLZiI8VKq5IqUxOmqj1QFyNBFg16rJH1Yc
qX8K7jkit0SRVOOS1jhuRDvJ+CBbFrH7ZV8C5oQUPwC8bmD4Ow8bkQ4gE6RXvQVtZccdkNsXLEsU
RRuSu16EfwfuVRynRMQqujs0v+8shx2LDr1sLqBI2LXpQtu5ErR2OPLjiGj/aarqxovYf8Hscvpq
ArI/CmMqqJx9cU8JECUoCaO6ZhW1rWAQdC3UDea7Iw9kEztVGjtbmQ88b+/kzZUjh7kq0GamoQbq
v0IymlAjVTaz5tEfT3TwHmaMce5/yc96QwoIQZJQWY33ZNfZAFz4hUTv4czq9SpKiXqQkqPhy0u/
dpGfzwdUc+lSBImhACV57+d3Xd1KQSqJVXJ36e8kvWt9/zrRhAPFVCtP8cXqQu8pDItTPRMdj6R8
gAZpqZTXfJtDEl83xwqGdyo7GDTQTmGAXjTQpCzXr8spSQrqAK3tHoKdcxPcmhZBiWYvaYo1+3UC
N9lrav+vjjithQ8708mtSVRQCCG9jIc4uSZgNtrBTNBL9nT1sCzYmOcLUH/WcE5HfpeMRS/LjIRT
5tITWZDvaTfodbNN/MyV4eZXMBJwpm5u7MVRTePDPmCMoU2QSTURIaTbdg9u2rGkUSfYL93ufFoJ
+qXx8N/R7IajnkB2hLKB8CGb9tHDQcjaVEwZiUYiplknFSNrXEYXzec8w7R4tPrUIXwZLYPb4J8j
5xXAARR7GOGFkC7J73UhjYQbT1IouYGLnvP6YPnDjOUQni04ExIYYdsUSmwqEIg3cxCZLhJNFHQ2
UnKL+VBJ0Vl9yUqE3fesxww0ffILyrP49t8KOgrk0UiwiXQoFsretLBlgZ/5/S+2MkbWCsumHfEK
i/WBkFQaUa0QsCyR8EBj95seVyYQQNYREb/9j3Aezn2Lpf2XK+a5W7SUZHlQfwu3n8sbfZdAPnQJ
fJseruVfADxR+fTH6BvkV7w65yWCxbMfa2x0AjHkB/Pkwl8QIJkusdYuJZPBlc9OWQkMScyQwtMT
ElkM4/+7cDLweLTMrSNlRgAE9D7NP/wJfZWcr+76Bbidh5pPqjvYEDf9CWxW09q10kGtf/rH2WDl
4EbA0zgr02WbJtoTd2CZdA0xT5I2FygLn3v1tyHAo71EHMJb62iqN0NQ9kHm/2il4e5PeeiNwWVJ
dSipWZHnt7MaVkHzamDrnEMHRIIRlccwAqUOk1OgndQgakM8JoqGjH58qZso4klGPFChjO7xqypS
Wq9ssachKkywi3P+rssPVfzZdXjqlYw3u41NPn1Q2ko2ugS/94HM8LU+6y5qyta/EaWdEScvl99v
qRRq/RA1aGzJIU5cOfo2Hq4uWrRSfVAL7uMNVCbWSeYmkj8R/viYTFTwowkKudBrB7uUyJV6CATM
0zmHbbnHBB5occpc6UW15Wzw0ULYfZOzZbzCK7J3p+yV6vHscQfnHo4M/wDaq3+ZP3LKHpYVJQbb
R17Y+Vv86mKBGqIWmuQ/yE5/Bjxt3fFCBF/98oCobavDKsFiwi9uVzcU+BLxMMJNjc5Q6ISY6OgB
sbw14ScYBZHCOmNZq8o1/yslVdr3DtjdjBGmDDqvYfVz6KCr6E+PBNeuVhLL2tfNKyyc42AYZ938
aIrYbfUckdGRybBA4qt8xgZDK431HkSQpwADZHbvCRn/ao/d2CKGNH/EgU8rpSRMgCE9uhn6KFPv
KDZkN+8IjcRNpQaOZlaGMHq7mCuzkmVIPjUaiFuu5rx6TT4ldRsn1QS8Ku93Ge2R77LQTvToOge0
QHXQEBr5LttMOMyRgQR0Jo3Nt43HLGCQvbCYc8L+IRo/FEqERDDWcVpuHDXqVoF0T7btyhTOpN/0
XsRTa3gbGcV4i1S/WrEn7t9c0FiWa7IPzCx/5UNvVXSlVIbNEHz8ZeToaVy10MSbcI7NVYDDX7/8
S+Cfk/ZCQ7vJGSU+Z5O7ounihKD+E+JwTNp/KSybg+SM5L4SR0UmdJWnRj522W/X84HdRa1K9wtD
gi9Ky2D2kf7uv5P5upCjhWB8KUh2r6xxgQKygvZtuyG66Hvoo1V4JqiBZAiVQhkElHpkzYytR4cn
WF4/BB6W8Q0euikcSxUN2+IuubLvyOirIviAN+PwF9tz3Cx1l63XL13oTNr9RSqJI7EEkUYKEl6g
VNE+f3dnkNvOKYPLPv+dDORgQ8ZRNDZrlqjW0NB3MXwsbzW6qCqd2xkSlCvZC5pdip9I424BPmDn
4N+A8DocTPQRElyS3hQ432gvIvY04I8e2w66HsbndORfVBpbAwDJ3PHoPyOu8g1wTdQjAfEhxJD3
qkzBRCk5vf8tVjaY/VwwLIgOjlZijdjsK/rfLkRHJOwYYW9zgim7Bc0nOJ3cQUwXH5B1fC7QSodJ
Tra1uu9ywver4/brn8ijY7wtEmNAAGJHiFfB8secAfK6L+eeko/PTQKqNAkOufiTGXQelqJPb8Ad
h/XjjV12UxAl7dkpOlxnAtQZSHUj1DasbipZKN03RgEUt8npyNrz+bGioW3YuiO9miP+T77tae2H
dlyDRPUoEuzLe2SDAUfpPFdiQPDV9PKw43P8vkkJrkr8EBYaTM08BC17ucg5Mb2EFc/vk1naGUlg
glZzfIAFSrUg71Oo5seP/qGIqtXywh3yNFa3xf5DQFhBeK1+H98lMoD5EmvAS0e3g7VxAmWfnvil
jWZte5Kvs/Zqx0rRnLJ/90hGbdOzbGtAvmZ+VNOeoSxlXBgIwYOtjjKSWlSPnmUTWVW4x0bPjXCB
4Kmysabe7e9Dsa/bu4BNNThUhBIoAjx3If5VqXAc0golpbYXzRh10uN+sdaX8PTxNmg+9EECwzJg
RDUNqRN8kr1aC30P3rrukQOMwjsa2uk5f3m5Wgn9tJGcEIsjy1bggvxZ1A0uImmlEqoQZyKTrro5
RooLYzLzHruNE2Ogdnmp/9vI5Q+qDPYmYDH5ZEhIDsoSQafy3WjjqopOxSDX6kxR0x2ABzWbv1cY
iy6b0vBjh5hMiiUkHW7vtPV5Z2BiszQ1WEgT+Ur8dyVnq2kcllSHk4KmmYTuFJ4fryz+3SookYRH
++F4BaNs1Rc+21z66F6CfHrx62VIXeUCl1pfF349Re1gqoTg8HGw+4nxCqC1ztfABrHAALaAEYsF
gzK+m7FB2l6GXn4Ggak4daifgcz+xgYVl5KPw0q5GxHcYhQWwcl/U+pU2KeWu6Tirnpo2AOR0zcU
vzT6vglj4vXRwDBRvzZje+8qxh0BkMIOcGAQxfILs0iH7G0x5hj34wA7pY23Wa9gFb89LqXzCiwM
xxTNLDgBePy7JvP+By6RDoMw/6ilrQvavf4Gh0/fH4qPZyOraQ0HBXL6SyIPKZK9fbGZB/3dsQ6Y
8xPavsncLrSkNGnKrfwUn18lBXbJfu3QMkgbBvQqVm2j/IN7y9+QFNE+xsT036igb2Zd4fZv/0yx
bQ6uu4QOCzSptOoEVesA5cPCX2DuNbYOdqvjgd9uKdKDdm9sNpClwJ9DrbSqS3gys4XVRs4GrPcn
lI0SIztAaZXCPGAPxIhk5qsnERqCKeHVX/5XR0jkKpLjjk63bk/KZkroT2oUVj/34Gjg1/8TZqTS
i07cvhTy6f5hiWNDp+g72BMQ4iQuwZzyLCAT2fbbhBfpWIKNuf0BIf3mpzNtXCE9oKxEzLx2bE3r
OCh7S8TDIqfxTe9sci2KVTTjj4spJ/bD/XpOXu0VmylkSxkPbWXrdY3qcz58f8tK5LB4UJ6dpezk
MZpwQXKORfCWdZtsT8Jx0o7qtvTT+6Iz4MNbeUiZtRcH8oE/E1FT84KBgnk+y/8QaRy82NaI3t5y
YOoZCXUN7cJR63Kcls6N4WxtLYTAO5A3hPs+WxzVMctbEPKFiJzMJWD5NgJVaP4S12r9YiqGMCnU
zfyx4x5dcM1t8SXKJ885GEpaRQ0R/gtp99eLnvYqwcarVd6EF5GP0u2/BogTsNpXICe+CM9JjBoW
FdwQJpP8elM1LqAnotDTNO+WdZvhV0dH8KePwijyTGF62DSJOb+XBw5Ot0JVftbFyoDbZK0BbIH3
ipEQBGL9ve9U6b8vmuXblVqKxBnzx8IJ9y/kLb/iKchtfzEE+X6dVX9fB1/HP3mtpETgdRIp0HEP
n2pKq3NlY94T69Szgnv/3n0I1CEbn03TEBgbXHkYUcCmJdRetBNNVx13/Zlj9kidW0T4lLCmry+l
3reUZjyyO/x1RJgyqseJIEVP5wFrFvh18CMV/vjSYn4Jxrn5yoRN3gkUANDSjo4cwXIu5++8t9+P
t++RAaZus5R3kare96CSeYp6ayBYvaWEgQj6fWoQAiKed7xddGxogtzzW3TiuHMtJF/SWDxFJEvu
QAcbCIsJHiXfXiNJv5O7hRTfcObAzJukdQzx1GlctufWGyJ/Blyuq7q9bxLeyMVGoUJpca4QSPGz
hDPoazM5ZwEeLv5S1nLsIntubKzHChHSFzmVLTxhFtGkBbIkmtYeKAA7BtTHj+gNphtCWPkD9COW
6mT4dvAeIR7OyRjg0RPk7qWjIR+2aJsSIaM/h8Ol1nj7zWubge7n7Eerv8oE0pB98ibWcvNdgwOd
TEULKocSndej+AzO1VPtvTIZytDriQbkMQz533w7sF/8Nda5xHZtKQoaIDD8NVmDkDcb8tEvVBxW
BkQSvZ+Tb6dlskq50rT8nIswRquSjrX2ga+1YSFPyJ+U1PTWXxRJUIWtGPjfE4/A5eq2L2lOI5kr
+ts9teu+hp8nE2PZuesBTpTQK7UGwLW485q+PLEKHICWYVeUsV2nv2zLvI8C34ULoyXOlOLQIyMA
sTivrqYSMbsAA8kDlqr3EkDpnLSS3zCwvoTfUbrigx5kQCiywT1OmZFfFIVOkGtN5WjmVYer8fLt
Wabixam5M8MX/DMF4Qj0O7e/ufNFG4t8LJWsoaohxzJUXmp5ZjoxXJTE8PeCP+LY6pcFyey2VVYB
trTMUwoYDQXvC8a2xor7t6eCf+7PIuzd8nKRy1IFEDCY7JP0V/pwRNKWFQ6RKzcV2VqHW02jBUCc
UEo0Pu7HfKfxMGDOXOZGT9NkO8WgpUKSSKlB8BUeOhdsQxfYTVt60j4S26NdhnaS22knOR7dQLnY
pRX3it5bm3r3W4PA5TeI/Shshq+woPkECSCxMBI7H0P5gmeeEZJWbta8SJujUb/lxINWYzL0miW6
0+9c+upHuiB/bds6uPhuGuUtO9EjFkca4uvfOu8sCiOweNXR6Ducki+HlPZlPMhTv9yrgsEnsP5m
0J+eAVtAk5MQHlFUyCMhhTpbWQnJppWJYYR0hU0vltPdERN0P49EqyhCrAP05b9tyc45BaicphgP
/9GtKK/nt5fN8tbQJacH7TdJNvFbCicNR7/OBym+Cqs8SW8foKxC9EIaxqIq89G5N/56SVBkG9wf
NWyJ6EUwqiiInIucjp8FF3eQafI1nbCjUR9Ua+8XzfiEQKC48ncy7K7Wr5fkaJghtwmViFOESkGj
Uekp0C2Y6BonwH22itREHGlekyqmteR1DwbYH4w/CTd2+2r2TKtwP0TIKS+ei1WjDd6nvKi6K04L
wYi379LEuB8AoycjenMj3Lii8oYicrMwRU5I85RsJPxVXo93+ULl2KCvS5PFpcf36C3ypFXlr0ub
qQ3SS6RVxlJxbh5kJbGzyw8GFQn1Ty+Rewxpuh3wGBsRybVdoSrWV6Sn/2c7l5/nUMbPVZj0zL9j
nx1oKPai1AIKLOJULcGqKb9c6LUt7HVspmsoZ3hMWI9SCiIFnmR5pERlvFe3rdLqc8bLCXx/5wru
G4/PQkQOj3i3a2cORIdthLl1Q089/kHz+BPV41dGeIoGS6GGh/UOONpPah94+IxNExxlCrymiPPN
J++hVXiYkRFoLov9lsUE/+vaESIY2puPjZlgoivDfXHHDBhkFnL+YgV2Z3aUlbLRzNHBHIO8itsi
Yu5tqbXGDlGs4LvJ7ifsddMIEvmEcPUGatdbneh1WSqHhJ4OhJioQQcRHM2SYQsu2fA/I9brfjyr
mBmtlSZu4yH+egKJbQmMUzgz4/4dIXmbSQE8v3WJ/37cUAmhFIPx6f9L3fZu+PEujnvUcP6nUFU+
uv/btuuVscfJj+Rfm4pLb8GYVYZ7d4Wl4no0U7pK7T1y4/JxK+Q9fT88GhPKBV7uLDW54hwdhVjp
+DFnzFMwMcVsUoPI+EiS0OnLl6nne5uBp2jKM1svYPadA3NWIJyo2B123upu1OwsbCyqI1wVgMQj
ZexEh9oJOhIBEpjaE4VrpSJ7KskuCXiuapk5jXzRn6x3gDSZsN898Dx94YkrIdjd/Q+gV5L+epqR
liRRCKNJBm+iL10QIL70pJjDhXCWqsrJzL144XIaZkgt87tzNx/8aQAfFnnKETp/0tngrJIhNGxs
yTLpnrOMFn6cu+A3esoJMKydBft7NKNx59xMW68rN9tYFoB2rqllTRwYKFFzLZFORwrgaCKOpoBT
HQS0c9aRZPmUqHkUz4TGYQl5/8d6qVIuxzIAsGOzsV7xkoqwfe3TAoD6HEw730IwDFgNCME+oFdX
Z3Ij2Icl/jzaQ/9gzyeme4DV8iGKicnCW64MW6SyUBpSM4grL1eAhHyCeONtNWfDovorR/iqLNJv
N3Gz1zY5Cveo/JpNtYY6dK7crDq9BGolkv8PufWmDBzAjSVSr8d59fjjATAoMcEgvajYTCQZZRS8
azJH5TJCYbNGo+eu4E+SzODRc86jnwE7lwYlxaReeQyfLTRk6F3PbTBxLvdfZBeiYCgVu1C1sFEn
RKqoSkhI8GIRZXX1NtG50ieRQCfz085tPn/q2CP5kT9n3332wtBmIAhP3UQPNWjxom1o92zYxPKJ
I71fjKVDbYeoSj+hl22fRU71+xPaIo+3bAyL+PJT8LHsVvdSO0j5wZXfvaJD8CQq+mLILm6KCxF9
IEPTdZNRhRXbfoa5FnVNPD5hT+0Y5EUoX9F1NS5ZGqlRrUZap1AVSe+qNAMfyFWlx2fqpPz+VsUr
hQmLLMsnSu/Lj2k0TjrXQ5ya5uoDLWhyLRe1kbNpYUYorHzrO+0ztc47AHIqm46hGsd55IUY7UZm
kzV9GXA1eeFWqCMXVL52c1sjKQtj/qNMCR+AD5kw2ia32CxmbmDonPZOp54uSlTU9xuzV/YYZyZx
tEV4l2/O2tmw4WaSlEWef9+Si0ga0Q+z+bU5h3fA2DyVbpRE1tVXjolP/8pguYgP5s/7xQgUKc20
4JcF5Bx3QyDlH8I4gHAU75QINlM531fnZal57U5XCy6q+s4UbMIswmH92f+NJPNuLtCWAsrXQNKh
DHkXCiZh63f54aPwyWCPSJr4ukCj5cc5Euf8YF+S2aaQYv0aqJYS/MEqLLNG1hfLqWk8BD8zY7x4
36KHsI0Kg+6eKdjKLtf1CpVoeapXvmQIDLpsa9WBH5XnqTuedOsACIU+MP8m/YHqytQ6bkguiXM9
JfjeUlmDjsM4XnaXPGl340rs8r0BJ/do0nghiUdbVefDuWx2kYvYPKCL6oWseqLg6UVz7itsr85E
+Z40iP3VD034QcFPAkllIsewJsP03Brrm/H3pxrb14W8LAEuep43UvdH505lXkcwigHErubwJHLm
2PeaLvbRrsmEjBuh8lLlaTCAYL152WxnVblxVdbv1PYRMcW0Z0TOaqvw355hK51zCrTXB4ZD+Pgw
ooPNB9hJ+G3Qb0XndvAmR9t44bI4tVfySdGtiszqLrMUSReP/xxpkTEq0y/8eVlMvZL7vUQEW1lX
9+M383JZvwJo9We8qEcQX+ar+oGUj4abnXa0cfZghUHGnfInvqqwvAvhg70rp49gBgTXwVX1ElMm
Z5LtFwBB5U0RIqYPJmjfxW1/c+WWSilie9HJHJkucBlZ/ndzGyylGng0HCm83H5s+VNf8I5oZ+5l
9Q9KJoKdUwCu+BucOJcQY1dEjE8Cq1/+oDnCh3RsV6oM+1hpA6lIdLP7a7Lpo0qh9HddlQkLk99S
vpNpheV3V6slHiMCPjDdY+92dYDgeLtjtPeAyLPWkxyGlRFcz+oqzkhcR8bo+M7IeK201jq53gfO
Zne3OhtN/sNKV4vscKLQW4djj16wnKqUV5rFVOgD2M7HJzGeu0NPLl103FmJI26OIBJTUMF13Lq0
UDtFbdHaT9KuTewOdNAbyz4JZMvXz3GeLnPez3MYeUhHz75eJ5CPA1f+pU54e03i3skQOucVFRpV
O1TBX9uRrKHHjPeN9WB2zXH4d85RzBXQfKtTwbPRU40nZD16tJcJ1WrsMpAGFPO1p2v2e4Wlcv9h
CJyTUZxFF7nO8hBf8XymbjsZFP6hHTHvVys7CAArN3JsP+CXO8MGbUbR8P8jCTMGD+oZUpa3hNOA
SZg3HAnfJ7y4qAD2btZkSS8/w0jz96mvvM0qbvga7FnmOd01JQIq/a1W94xKFOsX4DmzmmLiqJ2M
p/oR4x5NyISZ3u/2Mqrq5VGhurKVRW8fXk5WI7K+LaT3M91h6yLk6yEYMEjcay9x87dkcEdrbo80
HFeAyf/ajMl3bC42ChrJ7111DLWPGtkAtBxcrqncNGHA8Z1Zuk/YdPXdCCDU2rGaBwnI2J3G+06a
GOlnVmKkrmMnRzuFUB6jx2TRvKOKx1hgSPewZ6bK1uCTD7f5Ne3iFovUe9mmixwGeDIRVRcAn9lS
04VasP3LDKmvVbv3AtMU6/0q0+uq3fIjIJWdqiyITxSsuk7YFNG+1+wLGsAUrJIzA0v7QM+DSOnS
cpj7fPid4xmOinqFODEKiJIjvqu1V4HcCkJJJaSILXtH/VMhCS48ex+9IKecuNirhi30O4aAFvWr
hipj3dwTevdEmtn26ocOysaaqzVlPIUlDDqS9yFdxJZFPiB/hixi5Wb91vyZ6ksAMkGgjxSScRIP
xioWn2OboLW1dtjsD20fNk2513c77pybM8Tx5Ba2fwUes4PSfcCxnsNjgr999Zp70kOCWBZAHqrj
DabT+KO0cmvWPehTB0MGgDzMl69puW25KPZy8O3snIZba+abB8anF2JS2TmztIBLY4Uu7ae1GbO3
Mv6JhdkPdkXT0u7ZsV8JF9o7H5tVJjPD4Gj86ZQhyy4iztx7f9diWXMT+zuHZ2wAn/L3rddYkyJM
Z2gAa/X/zx/ldpjvaG3vig0FLoX1s7EY2X28Zn2k0lowXCkl4ZQ/4P5iTSh1Fwc2aeZLKH2J1bxD
Fkt92hyCp0Zm0uuHAkQTYJCC0bSYmV9dGf/tT416uJplNGgjgwgvfKdaZiWpu7mQTONP/zGG7bYe
pMoJ3vZ7Gsi9mlLg0YWZwLs22CKfa6UbtyfeSSDX8S7AqrKZf5k1VDupGvSDeTSEg3qHsfVcjTXg
Mo3zSDdDNFPOzmtuNTQHq//jH0tXWtmdv8D2LheLUuL9JIbnOlIb8pYMP6Lc0PUR5d90AnS8dFpe
0J8geGgYBIbnM5GgIvPugn/P2mKGXzXAfHoBzCK+bNBbmLH960PHprok+VffcEpm0tkpmgwwb9Ry
eRsFFpBPRQaRIWJ7m7FvjLSObNN2staT34jLAdvVlu8B+MibwnCOEJu9XF4pJn66palEBLzPP576
UCNXd7Af0PJuOYTXzJW2v73SVSwNydBOy41TGna1ATYc26qfhPGY8pgygBHwMaZ4yqHLkKiIS4SH
Hnj3T7yulrIGmd1ainarbtupFXO3cCyCVAkIWCxZ0M7zjySUZAzqVy0Kivt4GfAOjSLcoMIq+AFZ
/xE/iKLlOSznx/1WLVWsceVwhKUCkCpJt0DqWgvIasTmBB07ASP7D7hcgbJje/4k1ccCyh/oGotx
9ZgfTSv089ZsLw2j2sJLAEs3Hss7cz6JWjHqEWoju21bOa0qVdMM8TBC+qxnRtQ1A+cRXRexl04P
nln5+v0qjC4MNNg8ItdvJxnajWvW/C7CWBySYDpdq0ghgM0FJfxOnaJODqYr9moGznuBp4Xzy247
+PGMGvxr7sWo38A+ew79RXoCWwRLwF7iACwrlVMNHY42izP9ahfgr1B7vZGd0cb8G8aJRB7GBQbX
cryEk8DdLX05x//sSSOm46RdzoZdsFajUD8YYYqXxnjzp0AeysuxicN+Re/3SglfHlCmk/VYGcWC
GrsRaPhOp39cpxXKioWHbUUvRaDNnG2QA6EXL2y9x6FYxyUqOw6Q3tkGQnGu0tKWRGq0sGe9NWPy
GmBV9el6T1sf5+gM4s2CTrnBZ4WPVZ10zkBXjQa7isyZ17XABJ8phnNRfa0RqpgPNmdN0fN91Ygt
WW0TxfGZcSiJZ/vWyHPlgvu5CiOTzkzy8JLD0Jaoc8aBPedOtB6PqVYcy3GUjTww5G+ekFx5WdhI
+UMhbv4H21g49F167vHbiyGXMJrPPpf23/cMnOHr0eE5sVcLFAKrfeHN2CyZl8FijdfyyoIejPvj
4wH7yDsvfDHw2gesrVCW5YyWZf9eyW3nsur4a6+Fg5qtvIWGRfSBAbUJfxwfYNiAbMaFcu3tErat
zK3bNximJzh4zDq/xRJ7CqHC+qLcXRC0gwVNApz+kAkSaF42HIFkHZ1gnIO/WZMVMIpmNLFN7xvM
VCVyaxDl/HlEcSJq9bdt/5uAHv1Ts3YLWDU8otYyzpYbb6lUdndCZh1FFlUM3p+HXpuv3X4knryf
Vqa3HVhtBvKADAzKpE0cMtfYATwWClvtMoZaJ41RKMHusGRq96l5RumMzBz0NixngLKYI3Ln5+k0
h3eLLtX6LxBdtLMYKvt6+B8hckWQCvD+ED9zAXfGhMtg3U9f/w0zlpOA3mjtX4E7MkQID0PyiW5Z
0nbCFw4cww5o2dqL1Hao/nJ+qo4qdrT8ixCNPt4zuZkgsjjr6UNn71RHWh9WfHzoFd2eMWxL+N2o
M+wyLJiv4T9gyjHHx/wH9mBqjPk9LAm7onkZK7JdltLHJKMqrjBicLisKKY4uXcjiw0i7LNWjJ2m
RsKjJl1ZpdltktFXILSWmoVptkm6fu+KWf9A8FNrxHlIftsYwYRxj7FPW9l3m0o5fGk+uJektWx9
cSivzVXOhjVjyv/GC2JqlstKJ7DxOilD5Y7umWIB3K62tnVfMX2xjVbSH95WG6n7JmIHUg8XJP1H
NrLdesBYjgeuGI/M4RaleTrlvPSaEu4VFrWVH3hT1aK7Geft/YP3U6/EuMv27RNriXZi5W7L6iCw
CjDuwEo2iWVKtsd4pQovjIflF70UXc8FYaOEHXSmDVcbdajDxRCw67v1GB/eRQQJAKJN9WVZUaat
BKrsK58Olmp48jI4fby9sqN0US2p5Ch1FVSK99NS//o5pPkta8O6XkLV4tbn3jQUYs+SG5T52ZYL
zx5gXz93X1uzhlYJqAJ2EzjSwn3tKXC9YMYjjl8D+Wfhc71Cfh3DIPNSLlj1K5Ao0fmIEY/IOZje
cEZMk2M5hTF9v4XTxI+fj9M+ZVTvo5rhP60BbzrVrO8fNlWNzTYP3VyGT5PpeRLwQVPT3IserCjC
utnvvZMfqk1RAHG+Ksxn+EHlYLBVG6BSVXdflH9KD03kFCUpeXLBE2xM1i9g00v2IgtTPuR9i4C5
eWfU0iO8fj2ett2hwz16FI+/Eskq9XFPcLQSfHqmQTEg9hhAGzZPU4t7o7rKKJ5dAo3y44Yvy3J/
wwvvwryyM9PntTdaBtcb/q28KcwYDA4q/e2hgq5IE1qCEtLXI2YLK7SNyxYxJnIGKs0HNHa3d5cu
HeFskOaz8zWsauti2IbIJxEky55nl6wfI9qo+YY4fKIdUsCm6wPXtpUoMR4ht03MKBJQvEq6n9qI
qfKHr9fwHYB5btB75DfClkIx9XeJ8VmFpqB/ewWM2/2+L8DPT1x0iymOMvE/uoZYTckBsm2hyN/m
e+pa0HcnmdK4/b9ZzoRuVZdHkXEv6kXZsQDzH+p94A9+zKzajMox9GICZ2KmAKkaDSZP7dawN3gj
/Mktjd+YsyvmI3yFJqkC9qgVGLNipRnSjoCcrauErNhb4op6L4GixJO8rcuuo+J9mTduZ9L1cTgY
b5/uMtyiwbzdPeiv1axbWdgqISyjnM5s10ghKFnAyRqYbJ4J62pE3XaBffXpaMvFEYjdsi9lVB16
Yk0z7U3t80IC/PGTZnDgRj+ah2gG7Bw/LDX23dM8VlGWmq/E4ttMTi95u96kj0lTl2jI5H4znXYO
Fdm0aFj6Feq9VGS/ekOKiWplricvX3sAGf5Mrf2lpEk6d2EnE8VuW6UfGqNoRnvXitA8rodHyLqy
7cNND8qrwOlHohgdI3WaaeZyerRLmypatgVYr2oIzSh8r7xEVDmuaJZaByUgbSCH0Jio5XUzfitd
Kx51aUEaA4LF7mFxMVMmfjVtAEXpfSOigdhPDygGuAHcZlss8VhcBachrSg3g8i6KPTXD3mB1XG7
JIqnp8mjRa3VHHHZTniLd0sNsl4l6/nbjFwVDgFNQGIgN5B7Z8FaHPbZ7f6uEZpzqU7ntlzlUYrZ
IUcZ1R2/LcYw3gUufmbkMkOSkcWuaUEZjvrkkNNYhtmEWLepXevN0hX3dW2sJtR5d7IaPTRcp+Dt
5Yti/QDlJpUUODnjFzH9VO2IAuEegaBRmdeZZaF6fV7o5n9PsDzrv/tYgmer9FIcoTnNy6w4C7N2
vFFBlPS/WjcDuuWNNquKMcvBKzo2a1tBMns5Tar2Fa/TFgEylQ4WxSOo7IcfRLOatRcKLtcbtg/N
Ja4UdvvDWJZVgIhgVKjQbfDlHsOJ5lwHLWSaUQQ9GsYQQYrUmxPIT0GSrHMe5vpqWAw0yj7iLrPN
whrr/0hAjmZa0SKItmDi17EuSxKu1rmKakT+lv1sPrs6j53f2OcZAPwcnuwsyirRRAGZm7xlKXI7
ZFXqrj72B85+OwoaT1WjmZajo9MY3R9zWIui/LWZrsnnvTfL2mr3WYO6SRoDRIYhoRtqvga1hQDu
1NLK1m3KRyVjrBy8rGTwpl9CTZh0jFV5d6BHVCJ4CANkvQExxRD5jjrKmnmJVVdUwy7xrlM/ZTTu
uXMf2+YobcGg+oe1YHVN/C5X56D2ToGFvHyQdyZOo0fsyTXtaviTFXggWBaYNNdjWEqQJCmxdklv
XUI/BTTOWJyXqNGckrXMYVO2DmsoAuGcZt2zjYH0yamb5XlXf8iIyfFQsOxmPCVtKoGAnMXZCfZ1
lrDzFMpbo9oZM8lIh4DnSawLXOj0TMflyOzB0E90Os3mUgZPcDAqjXszMx+LPZZSKYBoNisCz6tW
KB8SqEVlYjTRhItvV1lb+cYGwYY67Q38k9KCxvtojr8KWY9+SgWfoBaE98Lvivlpjg6jZZ6fFkcN
7k4weve9CbO5GvUpx4GbUB2TcuGJO7z7UkexRdiRmZLWCQOQTaSpZ8qsPkjE3f4i5xDPKbMGvDHQ
O/6pxAYC887TSH263xFotIYi8tJVfm9TFFjxD3chuiuvFrhYUbytqEO3l9JMrHv8gAdAxk544q61
u1xD+K4MA7O7OcATmOD8C5LuXpni7AXGYNpM7fb+lA4QcKOZ5w7pL8OIdf1pCYvdX1Hor3PrNf3W
DRWNM9PvHL9gyD8efA0V4jTWzIQ0Eci6whplspvsB/dKZKYRZGNVpNl5zyI/mgdhqEMoYEvX11Mz
2on5hu+VYmS68YS8VUCqA5X+uKnkVYV4Or4md7dEJdYRqtG0R1pVdzlvfvhWUgw0Di1d2+JPBk3N
dKIyMc9gTdq0F+nBiSzlcMHeocTfgA35vz/630eY3x8LwEDHyGsozOin93WceDgubmrY+2BPrw5r
MDr3mB7fXVTwVK4YDE3u6Hk7tsVCwbnwUndv4zaBGzhh26C875fyx+KVdiWCTxXnwrNzeS989/8J
gtfw48MBDLxXsq5U8BtpvKwagvHvce938eaA/8A7FOyKmmDiVpP+cHu7EMtbuGxXgGt1fMJCnHJY
Ve5JfWUJyHAEgXFvaKDCYg7T3rtz1npg5ilDBtpLCNIp8KUHf3C2NFs4hqNzqwb5hkEKn2iCJc0e
uCJVbUf7Zx7yawIiH6qBHEF521lsgvgmGwHCdmqs+wLny824H0F0JD+21s9YjJn6eTKhSjUSwDRR
QuFeXnJ1/qD4nXxzhWmpmwf5BCuI1XWXuzIiWVOBSU8DjKmll8asEgZomE+s2cxa/L1L+ackYwSg
r3abQvwoaTFfurRGSyuYnbOZ1yHtOjw7ix2An4AzzC8unjLsVXqgSEOJM5e6Lg+16tDoTofY57k8
7wSUfnp+2eUo1xi2gKIHUzp7yneZmud8DIyLGjF1N6+gqR4htHtSr4ZJtT00xCGFE2d0Rwu4AZa/
pkcCci7ckwRIjs9eE1rOfkMz35STOezoW6te9K0+6OKgf5zctSq/nTPQtzCiohzbznWGRvt6BSJH
UxGCItL3FrwaInw53mjj6/N71Fxw1FdL4FxgI5Wvi1lkRPVfSAFuwa44EbK7e+BqsLIpeiZ9a20n
X2UZ92Tx7hzqFROj7g/OsYHIC8dR1x+dDDDSPreACgJGiklX8JgXObeUwWUHVA3czxVCFLgOzSRo
hQVHAaInmkr8oDvQmm2dALO+AKljxFScwz+4MuNdJseqgCK4vOBwCJyfdqG9MofLW6RRXSad0YxH
QesbNCAAmLovMJ4zyThqVXx7/HqNr4iyAdU8dOUtP5sxddOikJvM68/Sqmo2unP9DOvy6YD99GYT
oIZrtFzKV4W+Trsbq64mSZkL5+zmfEWg+sEIZk/EXf4Ify7/7pQxuTEcWC9GIULM8fwx8L8kNF01
2j9eDay7i0fLfApIYl/Gt1IzdSsC29hKR/ZDQU7ItqduOf8X7mc8BwdB2Ne97ZMiDUY0bVtyD4G6
HpRSfcUTJRT3CDhXfxxlBtBkw+G1G3Z8mMJJkihxJnkI7Vf1c4HgGi413YunwvEnZjEzVgas941s
xm0H3hA4SczHZmOjKm9pZQHJGFHf7Pl6ZTPYN1tHQgoM1DrselRy8IRNwdtw2ktyHd7H5eRzSYJv
YlLcvLU09HgYiMLUeV5Jgu/VITKZeaVtsXl/k4MYERpZY/HDqzTdXcGd5FhXf5ZX2EwnryhaseAF
IPesSgm+SOs6PYW3/pIxJ2CZH4KoNlGwLfGJYJGfO/Y49oWzqTM0AxIhKDC2Zx9AmRLWAF+DGDoT
7/wLpQ+vMw4t++WmCul81VWW05AyuaEBmXh3CXjnKLE5BzJMW17IW0r9txeaC5kalwUIf9rFpgL4
LVG50VkBoZuN6Yjteilcoac3ipnKa/u/JXZ3mKr0qisue/TT36Cyza5DAOCjZzMelkH3Vj3d/aTV
Z57C83Kq5MOEujYFZMdAOS4hRujVMhxXwRwai+N89uiAsoM7IQq2f3F0diYHisXmS/Hjn8Sp6paG
MNo7JkGagMm1uq/jHSFMEt+lG3Ffjn0JnGt+AHQD6lsvPeCrNVIyqXHsBQ+Rgv/M/YVfBBwZTxwx
0U4+dn53QKFB1Ei6wWIhPbLj7RC84rxcaVREBa5RNmpc15+KyaJCFo9NBLJy5IBlgP7JkkhB4zl5
sstkIuauUxwprs4p6Lo+QFIRsrvTOFrTTfx6vy5ZavWlR7j5DI/iUn0syL+9hh5KgECrdnWVFF7Y
Ot5kabjwLH3xYyYQZt9SVhvdU7cNlNoIfNx4uZFhWdLS+T1I1ghPGgZRXgWHQOfXa+2bQbAPajfT
ktnsfWKFU6QLzTM9K6FZ0OMbE0I4ZKmPcs2LexTxIS64jSmDLwfXssvqyRLqzrsP4QEmD45L4dYe
Hw7QxykgIdQQXys/mlhQrOgNFsubhlELWvbK+zc9zzXzH0H8miQvzcsnI/ShQ88Xu+xqiNBjAmxd
OZqUOXzQKBfkG0BtvNexyZEzfiJsrN3p7FQh7Oo/l1uIemzq9WAB/xB4t6xoSVdM/MIgMWEmnZqu
8jV4TxAlKq/Aa41PKIw9vfSXeeDFgdJA2l9wuCwIfqc2eWwiGfdAbRrGurEmPfEUKZv0UQ6UACQL
akZMy3cEAWOz35+4OoZtaQbVSzBtnSIUM96Zv8HgP4Zdlm0Mq3w9A4cGUZ+mUUZHFWRQL0bu815s
GrzpC37SNGevhbWYPFIu4/CFI1QVnP+lDp8yH0Xq9FospoK++4DuVbRpd+It4g3pBKopIjhJrAuO
qWVIxDWbNXsSFMM9kOg1+yO3a1+wxOvdjDz1UjAB9TIO/eQXYWamSiKXTkfDGXt8LnnGRMyr9pwy
svkjfumOIBnu/vO75i5zaNDjSt9+PBeVF5M6Cy2M4qmiA54R37A0Q/SZ4rx+l1lOiJ2NZVdxmWAg
pBaj530x2zEKnzbv6VAnOGMzhajhQoC+2etrW7hjAnOW88n9tff0f7+5qzs3scQfJKd2QJ1/DEu7
V+rU8iebEP8vFzN1Ls0Xz7xq3OdYxZcI7IhWuNHnaZnfkPlF9+0XYyF0EbQH++QvL9I0dtD4GXS7
aZOyBXbSW5MsaSv89jfSR3VQ4ruDaqLptu2C+pSA6PrB0omWxrtWII698EvAX2kjG/NYYP5kThOl
i2HECI2VVvnBsAixgPjcKFriWQT740XACe2R2gj6H+WrapX+y8KLCzKvtalrmXOw4I0XgsRGedZ6
cMZTulhxfdqIk+g8d4GoXNOycbd3jsOC9b9GZroYAg4QDCqz7zw+vkWhlPRM0obtep9JssyhnOFb
feJ2gXESuAqu/ClmZr6TIi51VkxqBFJpDWNtjwaumeZdkPzWLBKktp6vlNXlEcIvV9kZzwReYujx
TXybojJiS1qvTaQw1ofSkIu8ocBIXJ2PiotuWW4IVwRSn6xzRT/XayiRF7X9Xvea54DXknXHLzQJ
UIN2amsxsOp+zW0BxYfVYGUm9QTFnNxCehPmFRwvqANkpYpbz0Ks4teNDZnxN6Ms9Y1eX5fm2TbU
bxEyqs40VCIlLaqcNN9rudYKfvXPjlw23/nBMLwKTeOdQL4qUU+1teMsgz6T7JwPjRaRSZmv/EN/
a8gIg+4dmJuzT02RrCIrs+zMCoQK3kT6Jqi8ZV95pWLBlNA3DveIs8+GF4QHdl1O6w3sEQzUvfAl
Vu3ervQLK8KMU0Z31kcCk15HS0Mvw20gl30qOxdEbBKpR8NC3WgXlj1PLTilErHdw8rDVgSCIl/g
WI+VnDZ8bdia6nMeOvRh21TJtMJnfcFN2+IHL0D3lqccKaEt68w2HHqtl7ApBy6zlir9LPs4SKz0
qrpcOMguiXFlLZPUknUDkp5XLQzKgrNPcAzyO+OKtZWsY5aIpvWRtD37/ttgq5O7GjdSt1dC//AC
UKpOlj0QKuRUbibdu1Lib2KeRIk3u6jQN6qnABdISSD19PUs5rh7+hmNmr8GXHRBTiwjfRxSycp9
MngUoosSh7nqgKRGU2JBNKMM8q4ro+mcjDYTll4j2xdpAUs3wiFvVbNq19fxKK6MWNb5UfR9uNic
ZlaeT9bd02iifHnmGTYbkSsngfJJMQqtJbfzy8oh3m7i+pzp0DT+/mK8gCST28/tl1lbloHca9A1
iMtTZmMXesYxPhX/W0xHXBsb6klEhky7fjmQJxCwn0lmVbEE6Ud8sH5bY213L5UPQMkpPWasVi6B
XFNWQ+nuZfnSpMgTHMyPh+IszxLip0kYjbwq3ciBq++yZElnixOujD7u5edLwBNo9cDFBUvJKf/Q
NlF9akd7mZUr8eVPcBZ1XvI3VlHTsy+xJ6b3j7O6GkzRUTU0DPq66idyQWjwcWn0nbNJhr6gAe1d
EaHhiP0i6TFPzolX5ytv8KAwZAWQdkjXp3+QfVrfxO7x7FWVobHjWz64l8VCbiYFw7p+BvZe6K85
Tr2LzsyXA4FCXuKFzEy2PZ8tUoWMC4oXnF1xQqs5P3wLiIDrgpoPTMXLtoIgvQCr2u2JfEh4+2xd
mAj+TYlE+JFfBbKP3V/ERT0t2RccfWw9VxUd4JhGU0Zcsrs9o0AOMEDqGIEXX33Jj9/ubZcgtSgL
S+Vw5USVoZ57A1nKO80KeV+9JH1wQMRlp0uM+lvdZFLGJ1g9hItA97qq/m9mt6uYMFbcmCOn37cl
Qo5ASGGCteCX2EvWS52Js29mOFYXsi3uXy3os/1J32NqTsvCGFd+cvNdi9Wcp16n7lcmnmLsO8vh
ZvWZ7bTRSGaP6S2yyMswvelYLtTQ70K8+XdvQg1pi1baLnZHa50bE9wLA4tn1zb1/BEn1hEvrxac
e5nRn5StpfPJk5Zs/J4GR6sh80Ein2p482lAFKRtWSWJST3dvtLlpTsd/w5yXMkd0uDeDnD47ZoH
OyDbT5fv+XbSGz5CEw3e4ylf1N+RnykB2ti1nLgdcZJbWtWQeOGFHYMKvjq76zNV7p2VNMDjkUtP
R0MUcPf5mYxBwZg4FNtSJEhoCa6p2AV5fTtS67dT1RKv8SEt+/5XCPsavTW1lkj7/p+GqtIb2IJW
FJsppn/OZF4Ux5+StW8uyjSiiXT6aThQJByYEj1fCAfDoGuIz6Tom3SEeZIRNJVM0FA8M7KbM+KS
jY0bdu1FviESFrhJMPcboTDPcSOzYhY+6BJXOKnfW4NqGGNPJU6WSE4QQPm8M7YStzgFaQBfp9OJ
MYzdFJpJOVXuej3aFLQNshNedI6Cdj6QRKkL20JM3SNpKzsAfRFLvjSitSIlIvDhoYWjd6bjti3G
l80ps449HQaUTE/bQzR1QFtUb/pCywv/Nl5A4XqrQuWQYR4ZyOhYX1YcQ/UXZDS0CqGXzKhR/jUa
k0imld8IUc/dkxAtKfz1ng23VhqLTMopd6inxcKmRWQnjEg7CeMWx+j9nv4m7UuH3uElzbzI+riE
0xe9Q4pXny0MeTumrCTcrxD7rvHQdQ2v5yZSMNSAN23JpKclVpUPc9tm9sMnr24/rikqHEjzQ0Wm
ZDWOcPzdXBdFCm8BA/x08FKMNnf4Wjm7chlg7DrRijkJuk9pPWoCeBH1zYH1QZapO8dYQU7JLt/S
p7m9qCVuXsXhDc93PZs1UoVJ416t3wlkAeTkzp2Qpj0pBjKhjXXBpq/98TES/TwZOGXSTL3SgmqR
UmXWIFx1m08GIOzCneUa+241+HvEFcL+T8O6WSyO+caEhUZWMfmaIK5yEeiZJOuFSVpHHP7PFmUu
KX5zCqFccYZxE+FKi5pKXeb3iFL0/dPf2SGVqBBE8MUdzbRDyTuSvqr3qqBOSKtVYe7JwczLMZi0
YhOENKt8Ki5/Aa1xNUW0hUdbudA2IwNp9Ap9ITodfTRvzJzBuZFJvoxb4ex6YHcN14zywAIBBM23
eYIBhQzzQl0ffndDC9VBhSIFKMH7YntsinO/7iZudUPuT0Uoed/MLfUq1Jv20YbKA4gcrAWmPUjz
QYMw222UoqSLnx9MI1UxWPgmy0nebei68sAFj43GAZs0Q9q5qAMtM0RTaTACT1ahKG9VJASz8R0Z
NLpEm3CbqoNtEZ65GXyFJrhR6amgnJxhR4cFvqh6wdS9MAFGqMvUgVOHan5lRIAaxDSyHtI4jPTL
Kfv1u0zhOUkX2sB+qqF9lZuC71IJkVrhpU0D1VWUpLrso1yc0DekHbuLZCI8cfxL0nlrE1Ie05V7
nRpb8L/AaV1YW3dBWxcMXFy78OSb3oRNbBwLrSSqpNmgwgSutbghWtqLFiXy7akyaDhu/pUZzyrd
+s7HX58NRpdA7qziLrf8F5yvWtuhhgAYhLSUs+oDV6AFc0VuYT/JY35JB3IKWssd2Mu4YQAoGxbx
miSRZ+sxN373ucfdeDYS/+rYTqn4CshF9U4uJRkXb4yVdkTdykNDJa7b7pPa4k3yujZ1bXlgwkJH
WqylTuQjQSRf1e451AY3E09sgA0pf78oakcUeBmxBOErADnPw6NjsVYhbynxx04JVUsDRdRQhFz3
AESdsZhmJNr7nXdPG67l/Na79ro0ckmOLpjXbp4emwsM0QpO7DFgExnBFElQ2wd4maD66CG0Caht
ZoUh0MnbChGIrWNUciY86L8WWi0uQQqnakR5ltGRvWXqDhnjHG/y5kHK7QfkoWeHlOn7ZPFRqm/r
jPqkPvWUNHeGgrdLJ0tmms9FVky0ocDSnNJkD6R2simMeMGZKj4yZnVVG+cH9qMVVqQAhQZEqIKk
8jtZDHthJUoc6zCLyGmWjhVaD8x+n/+FuPZJOaaOLlVBCnQhz++BQAF9WLOaWruyIvNmTmpOZIcC
R4ZR2M/BtKJJJUoxG1KloTceoQv7nbfqny2vTfhYKLX3wAVVU7I+ECCO4rsgHmQr6BO4r9XrsLdg
3++UMk4vG+dNeeiwe/BIlXHktqCyN4owkH7sAtGqsVkVgW9nfIdcS/+odTrKTXfkBTTrHWz5rgdW
tEhmcNpyZHbbfwqSmouIanUy0w0IGmWmzqqEU+nM+JhaniXXz4FgFjCL8oB+M9yhEA2jYlqyQVap
xem2jiyvVh2Yh9lXyrcmoRQqPSff4k3ZyzTUmrrjb9CMrAgvgWL3BHv4qlurd3mziTUdtgpwEtYt
Kr0b0XUALcPv+zLQa6fNxodiQyIkvxeMHLgLxOGuKH+hNKsC2kLHLQn+jCCmlhmfShu8kNWSb8Pc
7M3a0RB5Z4QENhYu40JDaQHJ5eXQuf7cD+EXaGOU4Z/0XaaWeD7YKWT05GtQyenVGr42fG1EflO5
020Z9cWPn7JrXKP596u7+qBMA/gKr6FuZR80kHH32cgW6jxeHZgx+gNmi53Mu2azGwLmwVuhZrML
VgCJfOTMctY9y6pbaE95tMmoJkrjLVxF8V873hgosa7c/g8HROqnwGkCbpGIvHIbQQczh04Inod2
Q3BQb5bIedooymAC7uKwav02e34Nf0ZMEoZWKPFazJPDZ1u09fHCXiSFpkG4eOKL5cqD7CubafoY
a0902kONMjFRKdktAlVrMoQvEhChtD8+vQTYYQ0Zs6dKlJ3nhjq3ABgsNiGUaAXE+W4ACSe3Z8AZ
JAu5OSUoSsVFmpADWC6o+js9P50F++baTUUCvDUb4HPGJrKIzetr6NvX21DwCGSAGeu3qJnLvzsY
cX0ww7PisHf8aFfVxIgZw4sO2UfmoWxA4ih9xj/lXE6LTlzFauxz/ogrE/DHu50bTpl2RM32nXlM
gVV48CT7XCvai1Sb9jrEIk+Rb/vbS+jCbeJFrdUHosJJhqjunSYtYnwP18ukyD32kJokjuqQq4zM
cUYIsiV/0TfteL/tE9OCzSCOIlLBcmakGGIclfTk472Ny3xq2Dgd0TxJ2kVsyug34F8b3sIgAppj
Ho6LNOggzB5kHnNCvc66w9ytQLbUt7yfAHl1j0zkzKj56qye/if7FsnZAKC37r+8AqFKLwnNugGv
KM2CH1iyChyBFu1oHDwSdUFlM1ItyST/2WABQBJ/CW4OdhzoXm33mgF4NVbxjdQT7f5Hc+CBqkAg
gYCPK3d8IGB6nXqZLEYrZTF48V/YOPRpGvt1DlmpKFpltqJ/SPa+cajq/lK5Dy1eEI4jwKR2FKmN
v6IthFTxt5iee69g2zhNDkcVhLmd/8d+bNaiCOQES7sdHI9hxdt+GFhn1PKFBxa32lLa18rsKlem
d0BZFs0HS+9jchaQnjHTf8M68jhznTymB4/ghONLDDFz4iFRxaZ4BocEj502G83wGHElXCPNvKuY
/cwa6UA1O4sK4Ec1Ll63BXKw5LaHVCexLQnjIc3IRy538H9dPYO2dbhQ1WcmbcXE1S9u/r1g/6b2
WBL1B5eTniujHb54yUx3oOisD2qmZsftz2KNjijr9sywDhyhXk3fijBAv2IAfmGbLmqVIt4JUB7g
QrA+JpBbexdptKtZVEJPs5uqphBsbptdgwiG2BIsBsQmmvgUBq8Qluuh4WuZ8CWlzq8jpS5qX9BT
vlAOWJRNN7B08+JCh9KdXAV7sTbd8PBBbWO6r0jVGF3WuwArEWomYFNR+TXA1z9GYskTv5y3cqE5
cb3toIYi0bY1Yr3PnMFgwP7FfxfFS5jllKtWsskNI3sNeKoLoq9SVaUWNRS5ogj3cQ5aYfpasAJE
OnEofS0fi30m++Ry+W8kPWsBAupHOa4/yYxVWbFOCnl34gZ5OFpBku9Nv5E33zazJrnmmqeiNPGo
DLlbw8SmT+2rd7Afc7K0YQA7kImpbo2Ep2AjFhHdm4Hqn/NTOpcM9/wU7+m1qCCGzB9vmS1ilRhC
LokJ2oRzNuBKbgFi/vah0Th3ybZcHOM8a649SAomZ9zAlzCfjCf+lMwg5JpZiZ98aEMDdwxfF8+f
J49hxkdLfEMrzGTZS1Y3xTvy23CFLO33crl9a6ubI7M5UMW6AK83VQkvLdZT5F9svbR/0WZHiR3B
pXcTmUWb/6qzo3XqMe3CdO9q6qjoMeVhlh+TWIiSGaJdWOY71Bh75roOw1Ji7Th/ccjZOU9zdHkD
disDqxojEJ3JokBcLU5QqDqE5PuBIHb5n7e56s30uOPYTHiRYzg2t7ICWO8NzXssG3rFM4AXfGjC
aDXK0mp/6mb4iFmv9NEQbWCHmdUK2w0mwyP/N9niqKJQ0LgEYyqhOQEhtr6DfPQFrc4QOFvbsX4w
K9ehDYEsyW2xFg8xiaSOm75PcSoK1yTtdG+OiO9Omj4khYh/I7uLV3v0T23dQOg/2r98gu3hnDac
w5JRzzpv2QmjqoVMazPZQoXuEznkLZI+iSBaxsnluOxufL6Zyh7wNJi5/KLvr8sgpYj5kwUq0k6l
Aaz9osXnPNGgMz55Nm5cpW4niVPRkit7Pc9sDYZbW3f4hJy0jnVgTX+oqO/ucHoijAK2n1HEcZGm
ePvBOCRj/dw320V5pvS/xKbmPnbOg9D0ZQdIG5MyUsu4OxEZk9by0li5WZJbk1oBdECzq3ruDozM
D5mSJuIrv/lScTEswvXgfK+zVHh+HONiOe90kbXJZUzmcbpf/3SmSAGlvDwHqEh3scQwfCIFCKG6
ekfwKhLbfaHbgApjHpQJ9tuynsdNwxXwRa0fqR7QSkWGtFRtHTjnNXb3r5PeN4rLoZJ83obrmWpb
bO79HxxMpb26gtri3YhcbPeBs3raAQvSXD5gGVUbqGvDFA/OtM3VQ6B69k2De0Rv93NEEWOpQwi/
1qkcDTXLj75lB1xGZFpXC39BMd1yYn0Vi+DeKqYKTkeBsd5tWhec+DhZJ1VZU1VADzxf+CwmHvXb
aHXtyAmWgopX8UXEKS1yXx8D7v7S03lRv9lP7biqlgdeqrWzq3g9ilPsAJYGS1qkjUv3bx51XQjX
/4oZCdqlFeAILOCLRVlYh78gKF4GG7046OywN+ik63QdVYjEiwyf4ogad2Rtqsr+k3ravBiHqOK9
QFFNl1rE3Jw8mZLt2B1s1CLKA+kLCEAXNB/nJXbbZFIh2A2bG3+oODChrdrw38d+bi4a7x0k2VwH
XUOCZFv0RYqMDeM7NUVhYAXr2P5ZavHWtqcHAuE/gSBSw4tucR25mPdhCKaeQzZdNtBQtsdLfmP6
+VDTUy+ATs8sTkqXcpBjWDEn95BjHczCczja9Ij6SXkj7+CUXEyfjzU+w7sOMbC/bhmKV+jrx5n7
QZxI7pxNIZsRNa4W9tqgz1D728WDLdQqNR4Mph/C3fPK8xb74UnyMpmkHXhv2xQpfm3w0gu4Ysag
bys+T0lpQm1UhaLWMPlW5fbrIhvttpe66SBQToVMFbs0F9pnvdYegAqWIiLVrbtMZxlmSbz5UbIa
/itOLQNukodP2eqn0dolB/hbWFQnUmalXuOFIxdpVk3hh53IOE9ak4XXhhZFrVmtziM2Dua/NpNs
1V2AD6piSMf96rviGy6GjnZ1za9RLRR7wUiv8Rg8A/c5pLCUqatq0c4DVEBd75NW/qUbYQrXFZdq
OTjalmJULqi31aXRzBaDah9drlQz4jufh6H9NQC0xWbNG+8oxbsAqMZaWfc9+7coLlULm/jYyhTA
Nc50Oir9J43UfW40AQH7QFMOvKHXqs5MRLFK/byusROKNUQveaEEnwOv8AMGCDKjy39dWUgCQlcX
X+7uNRmsvCsjhx/LT03E50X+Wg2zZaSz+rWt9vh7Enc9IRzOQVWMcRymgUAGVOflQGlgx3ej0fxL
GEStoMEDBJAnLSlnz8A2wKFA6lCN3OVUIfqmOI/24ay0Vd0u83oWU3U6g3i0W6aerZXVLm8/BVwh
4xbQhjR9rgMWX4WF/sNbqrxEyLQl49R5ntDX+gJdYmzUAgRrFXvBUtb5nZyjJpdbxhSN9Eo5eLNE
3NkbzdkZa/Qz6SWX5AXE4/eOg3imF6JZRnvp6ynrZrIIqG6zB+APo64HbMLW+k8lskyo/+k9Whsx
so69qnY6yS9WMXwg6x6teuH0yzbgjVmP2OQYx1BaPlEs4L8hcnvJnAi1K3seWd40afgdg/MWbuma
jTDaqFpniIyFtD0mKrMTEKZPBJvhLbu1xlywLR2M2ptSytdGCOeMZzXcgUwB3lZYPpzUuBeLEngf
wraOCDf+TCtojLGgv+ojn85oM5qKBzi6xJfLWbB2zHVkmTlJ6KXAoHbrS8hIuwflqs1hJnIbRXSL
ku9b/91sHCQW8A3k35EizOuGpGNf+3OAGrYFTZPqr0HKat3DYWA9+ZFwxCwt2SQ3rGV8/c2+odhs
jRVSW5OAzlQ0ixVfG570onnOkwpPIN6GKOa9jYcLhsus/eimTw12498n1dGvvxiYEfZ2PJTIu6nv
9dtA0rA0RvP7rgdzU5amXR8gRUTVuBHB4Zn25AO7tbMfxmbdvnLSP60gJSOH0loAgr+QOFtCuOW2
2Dcgaav2IOd9Cw9mQCYJ5PvOtrI28nKFOQAoPO1lisVX9TceKfL1klo5jiAET4MDOVgreXBWQBlL
qmVYB0I4btAZfNDiyvQRUNd/KhU1u1wcJbIN2lowmlEScba56HotP0Puo5gzDgJBWy6g5og3XxxN
8DwFO81o+FfyRog7GJSb2iHNz+N9k1yurTsjlgjHvHisJ2qiBGwF+3ZVmovnnFkcBF6CZ2iGLj4s
GkUBG9wRfUQizTFxbIwJiPKA5xUooNgBzqsnlhCAYv4+KW5BmMW8eXFRx/ubBwdLNmD+3GqdCNde
vGUlhr4g3WLT8vxLXI9N+LG8uHp2dV2crzv9pqcEaAB34XjuGcbJ4nf2wrmvXTMgIUuB/hfpkvK+
PzTuo7sbJT51rahJQWtu+FV9ZIIf0hks9FkVhyvQh9qbYe7r8OcB2bS4whbHIH6/U4Q62tQh8lWb
sE6YycfYWlw8B68wzMymi7SwHYQBB8l5jcfUxSrBibEyZMPcZA/mImdbb1v3Ctnl3oOsSyZaenGf
k8jrbtokbVobqwJPI5IrhrsElNZ9quK1FK7dItRs9zzfuYNpHzuNAVxatfzwlPOyEvTWPCdgTfbo
ugh7mVEj6dAaTUw19NlFiUgeEEdteYxtdYg7ravszf6AiG8nYbBEYM1hLksM+5Koc3CikM0dN+O+
HNv9ae1BAp1Bpxk2fIV2VXrbvhIC+VKyi5YXlfZUwTR0Ptxsz18/Q5x8JfoOBeq//ryurhVgGsmn
pkc7z585SqVCtN9s5aQyD9pgMTmqTxrs7p516hqmcJwnL26zVJN/U7jihJIxnHSRHEcr5dN/yt8/
ZSFzCmKGeGhuLJM6JsgSzNeE0myravwkmh0SHdVkhCA0x6tSDCNpuWHdbWShqpx3fI1kfOpvpSIx
EScCDnA4Ng1Gu2FFpnabaB3TQ/eB9dn6YmAtrmXhL0lpeaD3dFKNemb3bD4u02nQWanRA76RvgwH
RiZrgh2r/mFpt/VQEeybV9Fj0o8NmrG8dh0AQ+Zv5Yr5eevmCcXOSOHll2MUhx9lqcajOELK0y0f
jQYITBB0D2ie20ATpk/YWW/wuDlsLxEuigV3j9yvO3fhqvIdeoXK5+PUoLp3g/+o1ft6R6oXWGop
3ulreNpDh61sk+Xcxb+pnZtedCjjtrK+peFQAX1ZXUaYhIitf5SyfeTPvTJJTbUc6vqccRVFzK4T
8dUiil8S0RWHroZDME4k0W/7OXd28dKKylRY0L6vgbDaDuyVtrTfnnW1NMwxS9+5LRUQHh/VP7h3
ArMehmaGLFG5yiHGhAgtZJuEb5AY7C/0lQs4TTMfMijNiAX6/Spo43kuGYJZNY1weiUZhWdLnPHx
4fNGy0CtwkvUnwM/bJTpNdsGMz8Xsh1IPJWAKLnGOAZ9zx3W0dC7hCyUcZacEPPjf/Jm097KO8Ow
XW76b5kpXSFnoPKq6VGfv7yknARqnErPyiy0ITxtpZlMVAowImtwVkh9sPLWigs9kvhocqmQ2vav
PKlY6nj03L8cvg/3XXOPs1VgRwACJjuap8WzGtYT572gnLAXKKjPBVehpwc70fi8FTOdFWmOOUsV
tUTQWaH3VESMNshkg/kSOgFMYC0XBN3I+dnS/dVaf4jZMd9G1DRWT6aeGMXa9FVl14NTIaPKonxd
d+gIMyiyCcbGJnVzbRZZENI2CGQ94WfXjl8x2e+Y3sG7d2NwwWA8U9HTxDu99qgFb2B7gB1Ljn1u
+9lqjAaTV2dJpvLPJRQsmLfgYmg8ZdYuqQBm0c0rsAgoMjnqePWKPFh4wYKiEjGbl6Co6cEFFVo/
MSh1ehzfOszUtBCpKDILzccvxW0/PgsU1Bbx69D/3OXMUtuKFt2VTy9p76dQiLvDOWhWnRNyUea3
DiV7zM+Nr2U2G/DScfW8p2KeBpSxybdHku/DEdQvGwecLJMzaXMhBWD17tYOMG1Y+v2kCjPFsSg7
bwbb74QO9U71AkudKL+R2AzpjUj/RNCg59y0bwmmPMkIcfddZ2nZdR85X1oTf8z8ifQsbQBd4u7A
sUexKoLfqKESwq7n94VZ0Axc57HcQR3oMAfKs2t6Irkl1+zREqxMKir1Rf0tAE0W3PPor8SytiYI
hkRIcekDjzCKIr4ieZr5UnwkyncbMOnB/WoYogoIJXiJd4Vitdkq9xbskGhkngvYsfOj8P5Wb3vl
47qMDmOMh2WY/osbCR6H9WCcoCfo6aUq5hrhVuO62tX3wlyU+gr9VJKuNqGsrbpf1/ulOMyTAMsO
Z9b01Q1sWFdFXUQOwwHK+/m1Dp9NpsVqfDb2NkbD2qJ+cpL8JGE/BoIzi/dRJdL4U/fOBVr1UN3e
QoQOLmfCiZJMenpmTfStB99uHfOGtN+2VNWaEoY+yaF7Szz1pP9GUTd8T9ey9db0oQYlXfIwKQap
YvaGbCVxmIi48Rzh985pIpV91atMXK4QhbFGJa7mCO/lSw5cIWLa7apBcKH7E12oHkUT5M2v29zr
y8+h7AVuQDXmLR8eAqAK/K1xgrBO9rEGAw9VUarp646+QwQFf99I/Be3MTSO+mxrWgOq/MKWUvBR
ZPRLEA28ZWYjOGPlvYEtHx2zMAASFgRjwbGNiAsT3gPU+ek80sQ2f4vzyxXFnMfkMDivFGms1G47
oJwaKU86gET1ERqsFDmc8bOj+zR9xVyhPsR2QNUeI0C9hZsBB1w/3ogJl8W5gnBZJJyeTUZI6gKC
OaIVHL4xg6RNY67A2tLEQU1NVxeU08ux/478AnaWO150MRHNKFRBUoWhGH8eFD2Q9rhKyrWAyrJM
VKtiJUOfBne7vI0vuH1b0yAwDr1Pz/l0nHQhqRf3fjkmqLS9cbm6RlKuJcpfGyXIdnzVe4b9UqpV
QXLXPrbFwE3kz9eLXEaSmtExk5YZHkiGMqObG8cLTkQZ6b7GqDHeoKdIbWTcCWRYNhq7z4x2v0kg
3xpXvabWNVBIV8deoUhIVpaXq9cGRedF5qG47DoVJUM31ENCi4lPq/nNTAQELcnxKbv4zZt/ex39
AyujyL/ivHmySOYhVhFehXFtyT/sd/4T1ZJ87HXgoLKKYHeb9+ZU7D4VymKOliVNGEdFfJhaA47C
WymtHl9wk3xEe5VWNR+VZ4ihGoc2PELgW7e+rn74VodNbVCA8yZ84/qcFzc/Ce9cFJ5tsNJxkz22
MBmCGCJ68nE4fA10YizJoEsPIv1IAd34OzpCWyaVn8z0rh7yf7omru8Mkaeft4YuF+PG9lqTkS4W
f2vl62rNYFU5yVnb59btYLMkqT1FWaYtwWIqW1RRjYXGhJmHul07pqnsmmo9Lykq/iFtYaWZ2ctA
cP5SXE72I4nIfFH1ActwTBGjePvamG116CREMoghFqxRyWg/S90r9mioPnl3RYSOX/Jto+VW6tey
p1Q5CZaez9Pox4IiFBqnJHA9KvAMDQm3tp6OkY1vPMVk9auxKUwe05dkspvyDa3VCyGike0ng7zc
21ic/X9oR//6pHUohDmSWcgEYcIxINiWW9jpX+qJxDcGeIFe5a45eYgqIZRAk0G/hKhk8B9LYxoC
NCzqpo1beAGgIEQb5dLUZUEATU9XCnYMyFYU4v2Pd8esnPquINlVpcJZeUtGBYynhovFLyCBPKTN
sBRDwAlGM/ZIWYPpSeaFaSG4abydeEB8qwd8XGhznguBJOoUObqN2CXhqI70+R7GEBPocKq9L5jG
PJAyOdcYSQGbYtX0GIpCLr+mElNX25rry1zRfyLfdEHcXbebcmkm410MT3TCUVjvEuKsmr04Qb7M
RbjCrjW1tfDhaEuEXQThQu9mzc0Rd1+/92YE/+l/uupO9Dn/S5AwyHGnTocYUEk+vUrQPvOrx6op
LIy35k/Ij3UDfs9GsLfbGSFam24jB46C8396NWDu+aTsd7uNVHNRu0RJCbjzrQ+oZEntku/HOhVa
j/xIauisvOp6TfUMr/LD74YBUkK1Lqk3Nr3Kez3ayfCIVqMBn08fZM3ieTxBxwWRs8JbjpX2k54b
GydZrfLxkX8h9McJeLfFAh0mlBKzs8qzB6vU42kb4M6m3g7L2NpO3F2ackQe2k42xXSkicMe43E7
Vak0EXQ9uYrhjDKMuGAax/n2xRrQQDSD8Vq9hv7FMUEbVElvMauV77ydZifRwq5s7Tx0pEVwT6g6
e9R/8H69ri5cbYpFzSmYz92BRk8NcbwyO+2gFS0tU1E7Obq77ZgcvSypQOxSZNJX3NLWF/4OpXhq
RKIicyUROHV5Gy7nIp8uOW4gIfkjOAJcs+nGfSwyt5J1d8hX7xa4Tc+Q+umAczgmwAcxeQh6Mv7w
ydM8QT7vGehQGrycCvpKCNNaGhUi8Eip8HoNLWysNQOxUtx5UFx4ThoZ69P812KhWA+rTZ/vbDIV
5CEyse29f7N3DbW8J2OtmLscsWsQTIe1B5DHl6od6JxT/Nw0HYXCp1eoKXm5B//u9NoREEnMXR6t
qF+adq0NgtUqocxS7jlWV4vKwypwaf73o9BYYZe7NMnGtZVKmqt7DKbk/p3PL4RtGcZ68gPXX5Eh
ydgdKYD8pP5IwhodRZsx3SCAxj7TMDszOoVa/WebD7Y2qEyAfYXTuIEev2rjpCWiCQySfczCPrIC
ve6y2Tl2VU3pT/XXxDDzwXgSy3i+kb2xuDPl67MCLGtCuHikjepE9Tp0dD8GgN6N8BK0lZtuXgC8
NUqYSvVbVKqiw+VFBX4bpsTN+BgldWfTC3VX0kdHwD/iDeQuOZdsGtwZ9XTwX6q2sBwK0utaIGq1
KRmX4roNKtK43GGE6p6uANPdZElmXDLDEFRj6ULbEGMF0sob4hpk55ne5Cd/gMBrnb9EWEZNUm1l
VOjqKInzbEBH+3r1CINSQCAL48aTYOhj7R8IOMAKT5d9jLvJpVx6x7RKOKNrBchQdnLNGlV5hhMO
hX/efTcMBNvCiY7ookm9dIJjPF301bzJPMNs9QOIS36IkloIol4cnIxIP0ahA7a9+4ijUZvmG9il
xmg8rR9JuvZLclLF9AhlAdnVzNTdsLxQmtW/CddtrwXXtJblcvpsjhKK/KUP9d2xBRrE2Dx0SR94
gdDRvCDgnu4RgUUEVcAiw5pRqjNs1XNjUiNQoI4g3FZSIKYf8AqtRO15cL1jmwJEzgzzdH+my7fl
ueiIEnnCvCmogsZKWU0moz5dcGTIH9DWtmN0+0ua3iJwBWqWMlT4grmniHactvuEIBk3RyssBXpX
1lTBJ46qr039Qrzd0H2t1BA/CW40ItqNAWyjjWWo4kjdg3XumSc95HTtnb9Ct1lYCkGDmvS1SkOl
2TwGp/bxp285xDOroqRrb3fLYdXCT3V+6OG7w5srGn+hDwYYfzlB9M0myhhxwkFyh4SQ8v1gtf7U
ipf1Utp216fzsFcbbYdusYc3omqXDMBXG0/g1ajxU/MWbdOmg3eGW146mnn0Buaok0j1w4a4fp7X
ICgqiWQGc2uKI/nFxOysVwAfQK4BEZ6POL1h1cGcabMNoZv0U/8i+ChbR95tY76iGAIKVA9D2uAn
uCHA7hHdbxSoi0vgVaid30XmjWGC5NMkKwZ9atipAN9+eAph/4V08k9mkSzreUI2MoDmrd5q5NQQ
nT6Ow2SXF86jWiSHB8SkLWMjmilAGVwqVlTvpx+pT7mApm0Cov3+ry9QLCVVEeCr2LInzr0zdnd9
4hecZ/HgZwBtDls3eTnruZ08eqNIp0UUhYknmxRM4RxEVJwhXheUZnn8Yo3FOBRlqO5dpzdgngPI
AoyzSnZCkL9dZtk4MRocngxtrVpkaGcC4HBgUsY6ASPy4ag5a/M+mhsAiWRUxt/t5fBalTFuzpZS
9GqWCxFduuqHwKA1R//fpmAMiL/chcmsiQn1FeinmhSFYEKq2OtgkSak0fP3vpl0szaMRbVMomjd
2aRVHouSbT4qdXoSAavMyGaAb4QCaEEWDmsRQ4lK4nP+hgL/jQ3S0FIB21j96s4SauQIH9+QXbv/
1Jkw5m5jMeLfrtOUwxM/QBc3eFpnA2OecAKZkiXbPu5zlcxZIeffi3D1XfigqYL9O2svQVedXigR
RvkgZfzSKikwGNja6A4KlalwyhUrMomWUQsvOihKrogqWkyFSITY3C6mAi8Hu/S2pCHT1FEodPqT
lC2giFYa8ZMqj+7GNzVhUZrKoa9uNyO0mo7BwMpqO+A61zNaVsRDPuQKgqozaUXwDy6O9gHw47df
GTWhwFfhGp7eebJL1B+yBG0PcThPo3aI8uU6RVEBio04mCBFvOJa3rLmx+4BFwgwr3kR0pXBXmeY
J7zjeXffTwzmS1pm9PUD+kBAAO0C0Rod6n38nl6myob8ZePAEGEjxpXm19nLuf6yOpC34IyNXDMA
yGjGAHdz0wxoPHyvYyb7mGyFCC1Nswdz75B3Apwc74Esuws71ZKS5lKwoAC+LKUYXapl9mz+fVM3
1uYb31nxS2fOX1rTOlv85aw6aFtAI7hKcaDOlZzH7pQVnIoCSCOKWnTnc9u/gGEWrbpZnak5zHPJ
BSgOXm/RzTnO92zF6dX3sQRFvPmETb//FpVHQOe6tgP5/+xImAlhSdVT+zrpCChEytBMR5iI3Osc
FCkSZbkx1EXJqWLFZEXG3M5qyruaOc2ky+2Xyw+o7QEhgBqtXa7BUYwrPxGvsBGOBJ5uPgvbzqS+
EtSk3DFomrLyehWTrWXDIiCc4BjLBH3qWs8s5X0p0N18oID7pk3s3FgAy9EN4u973cRU7PS91XdV
r1QyqlWlyZttwHZLDKaYkP41yeEWQsoaqdDLwN2/VWmCayI0gpW0Kr2F5lh6j+GvTcuKIOSHdKwa
G/XrhVoeADJISRtpg0PQpVXmSXwXuZ2qFu7Ht4wfHA73rYjIgElx39M1nnir7F2sJrAPDP7cQ2gY
4Zg05Ct8PUaw+M/j/5CWXUdvRVNPleqpAD+w5qLfPb9yvGEP7ekw9rODndjsA8qayRBksY9cm+uL
kpoMlKR/yjqPKqlPrV6agRDGKN01+O4Vb5hlMfjt/is75U/xwGhOKJobB5cCuCIwdcrggKx454F8
rZaRcPvh8gQAMmMLUrFDwdfYmXVZMJT4FmqIkxNITrthaYAjSag5ceuPtWtrZPUwcwK5TwBLe7b3
Kq5R+E0g97isrpPd+aVUvO4ealOl2A8W2ama2OdS8vJnI9cLMLa1bmbtBKHXsuARMe8r4Lyy9Je8
L1D6UKeaG2pE1UTp+9eNSrD+n1c89JW6IlBd+skRcybiL2pkzYcpMxVUOQp0gm17nZanpGfdVO9q
u+dw8XFhynNj6uGmDHF7Stc5VKDwM8kCaiUqy0/rXAaCA49ZHVxFpOsyHyH/uZMgJpvYv12e32gy
AravpDcGbIMAPx34XTQj3yhiFmqahrcQXW0hUeiRUuUB5EgmtqZHAUHs6wZydQTTB0uvf3Aigxr4
VM2TZcpsTuSNvX8EluNFkwn8JPizUl5DY87biTW1rk8lrAMtI1lMSnhsYgDUowCfm4k4/vB/LAM7
7A/Ygpditcf4G7prkNhiP06NRvN1IHiwh7KcMxNHbxdHFCT9Hs19oqVHAxKU1t/PwqKY8iO15BcJ
bEsLcgKPabV4IrvFG+4q0tsfIQ5H6N2QT2AnYz9QPm7KAlGH71JIieI8SwZS38S0Xnuz6pTKSmI0
1q1KttpTFEbWuyUpIBiNot0MhDg1q/lVg/a+LigjI4910xWQVHpIYWdS5ygtJIrorM5VBQ8e/1G9
yIWNxXPBX3sl9FCn/H7lT0gm8VFhxk1YXpmpVFJ6+bhPIVgwpLDrz9DTfh2gEKcowAveNiGyIiXI
cSCo34oN+4zfW5Rw6zeDT4T2gVbo/3EVJDPg1elQv/w9Ax9xYh7fxMwOxNhGoBhN6GiKjhpA/TiA
vy4Cyehn06qwqbIoKSpOZ4dsHRh9QWEIyvhE/jLuvPEeA2kT89abSMHJHA8amY++s0GXJXArSMzA
jIZ2b6gbucRkq1zah52jqC3E4z9a4voHsG+2mn+Y21vwCZk0qRwt1mCcfCaCid3WL+S8IuwlqYkT
bSISJ3mDPsxuU/llZFBcayd2HR8fja/YT6xIW0ByeXcAKLRq7PYXoS2//NU0EIsMiknMI6JfETHQ
DFd54sy9XExuGmIoKrslWRmn1jn0Ha4zKLRyhtrQivNf1cl9JWWvmzNf18tlL7FJV31tkANy4vIW
SQ1jaQZKS+2dF2vqXStHtrJDZKeMk0vgRB02xiqdcS5jlXb5aEpay59L6wpyJKLWdABwFbvYy+bP
1Pg35S5wtvzz3zM2s1bhuTDh/e6ghBhLz1nU5nfN1b9L7F8aQxPJdSqsjqqR2zmziR07TL6y/FPe
S73b2ZCXbAtzZZGk418qR3DLo7miJDzSa9iMtqrovXE262iwBTaHBv9LT4HGh0/ApvgozQxWeo7A
BKiAxFdE3o8IjxTgvUPgM88PTmchVRAYrAz7ZcVBOohFACvm3ERP7VdtYYljnKRlzVGKAjTY4BDo
AsQHHKzQ/HAV6sWFQo8CR4QjDaMNmwFh+96O5KJEL6PTUHuokaogGYcOhOxNy9BNNdY/7JfbIMHd
iIsaY2ipA9lDr9xtupeE+cG6z1kLahCzXvYmG3IoMPh8FLhm+oVHZufVPeIL2B0t4zFvq8zPHN02
wWsrIs2nLyWxzfj1R0iRa+7umlTIZU31C8vQzRzFBBOSWKD3D1xIqQ5t1lkJaDtBaazK1O4bSR2s
lB2O5ro4WH/f43yaSRrbo45/MDfFJEWEsgdw95fVCSXztERyEsu2GMwizuBL0BqATGi/DaD4UGUr
vJyWG6wCCT421ldDUZHGAijK+QMDBMTlcCE/HHS9kKhR7HR5Y3bkr8iEwgwjoolUf9dRZs7Lz17d
mhoqDIavIYuhqx8VY32lg3etkgZPy6gHIcG91nLQD0sfI+uOyCx/Sn5XJWcVvpb106VFjSC4jPgO
M+Dc/osodByBfzPadXk0ooPKBd/naauKEYuHxgEApvdn8xNDw4qZuO7uffBUZSlNgKTL295nmioH
pzzYBfsXGP8En9kKyazTHIuNiSaBFTyx21/JmnH3lWUihBluSnpG5TicYwBWSPUvCqv25la2sqHW
04WPVZOMftge7LBTJs95RrSbsqcS11gY0R7DqiDcAGybNqE3GGtqvq6s2piiKGyogGOMnCBIxyJx
higMr5Jm+yagFwv0abjKF3xwVlT+9DF+EWKnIxY4+H8Ov0wwMFEXbqXzBySJM9ggKe8MPEw0Fzx6
WHZNq/EulzHbfzS7njvMy8gL3JgxE5Kqv8Q1pQ6iHD98EMEaOXtNjAyvKEfvJdAc0mFAiueSX7PP
gWfSUEDo36j0ozQHlAiJTNWZLMBtoXPvaNg9tJltjClazLaLhzAY7fLbVW0x7X3V6vJADa2DLOmi
CzFuJ7Cgu75RP27MhuBdtDk7oOnn+CV2BZNrW6VYGVYt5yq1sdWiNZVPQxx/YW/YZ2XyzWOmNhjb
ImRlRX6dstub1jHuBfWAoRu2dT6sxsmgcM+IaoPdTrQOMcDj/5SB2kuylKkiArbk1JWeCKH37IkC
oneDy6Ou4VJBMa8LSBvQsK4YbE4l8XbpNhg9YvzUJIWciwfsTKelHPnEloF+GNFGmC28ndEPERfC
eP1sfOq+oExkkuWeDn2Nwe4OeALsjHeLPp7HVUek+l1YaQlre9sef4Lqtw3kWce5jBAQhFFEpwu4
KVkd0qwk+fos1CeEgXMXF84wqepQVVzhKfnejS/hMTgo9ktxyD/yTaOxenY+n5ur7vCuz0uYjIRA
a94vSWH2OzVFiP/fdy9PqrB1XFyc8ejxHSmPX/00/AtJKaoxpcMSoug/1Tq6yECOD7K2RgE+OjGF
UHLKu13sIbFgjaksN8jhJ/9n2MwyAdHuJibQkQhseEmh6S7yqHtdmFhGcKdD0GATrqYpAgi9GHXp
qQoJ0WWO4qTtdNXqfGGxSO4u/tGr98hrqfo8EDCLJQkSlGT23orxv4yo52qkzdDCA8IMSjTBX3Si
8JANe8GFAVofrB8segfnoqqQapyrQbWtCrppaG8MifZpKUIMFBAfWxDvvRk94G+r3pdVrY2136ae
YzreNMbe3vfbdOMCPePE2MwGUX4LSgT74kfYDTnx+1NvRg2F/w0LqY8F+dLr6aYDEvz2W7TLiBpO
wCvuzqSJ0oNm5JNScjaAdOAV+9ixsiK/+q4H1+cA9K2D4/IVwRh6FIg72FzTXlM6qa0kiAevaGmQ
iiNkgWliq5ULhFPFdkU9IT4okQkUe/fQ/qUqxoIbbqbz5Iu95zrLLDiNMCRgy5sO4C3HGKDwOg2E
ezoLbeh/SLGsX9uoJv6tgkL75kqb5Cwv5lXZo2qfyzFVWk8zJ8rz/G66hAi250T+z53/DFFokn5K
si76nQ/29eZgq0iyIT/fT4gpulVFItyIWRl4vVW2/rH1PHfrftXL+TS5XHYAk5FW5+EfxptCWIfp
ljZByImyzPQFUrcMmTFyiplyLGWHEIKUwOmp3Hbg0lVosqC+dMfNA0Ps9rNkl+kENQKE916WZCDn
YL23gDSeezucndlEo3A4uqy/1ZH5cFB/VkSXIm1qElgWhfp+0irxpysWjGYB8BvhS6MzIuMAkR6Y
JZMb4GBCtlJSN1/gOp8CSRPnzwXNCTX9OC1lILvNvBMOLJx+ZaRyW4ydTQ30jF5c5wB9DfqFBJrM
wU2U22TykVCq8c81/vQziqA/ljTof26NZI1Y/f0MXvkZoHgiREjA3331w36gU8eYTq1TUprG4uhM
+6imiCw5IWiiNDX2tqIQSnCyD4uV9e4I8J15Z9Fg3TGZ8ks5QnMqbMDNr7lmkBpvFqGSRtUDjadW
/5lqac+qe4Pm+WfDeJCac4X/1WW3aSzo4/DM5uvcX/bBYT2wiD3Ra9FybaTLzpvxOmP91NZsVM8o
I6T1LDK2+yY5DVvHFxvWA5HmUe5utxCvE/c2/zkdstyxVAns+eW933DVgKTEI4rbqPOnhO2wjIBP
rYtvNq9fC7g6EyqNNIEdxHo190b4/o6bvE/eXfxNFQWDXZucnX3wCOOcTlmRaQAFIYRir1V3HZ7A
mDaS40yUqS1d7K1p+Dvw0wxBvvLl2jQkXFjxyI+qWDU9yHjXoRJKjsg3DT+OyWWnXxdUeR8UDWJf
AuM6oEfho7CD7WA/Cj7vf1MOfeXE+TXqn/KwfiZEdFD8csuz2t2QPMv5jEBqe5OWgeVqSbY2eWHc
8J/2ps9rAMDHyA/TstHRSthYFVxki/6DA0pSQlW43ERSFkmPGIp7M5XK0n6tY0MdQBD/SUgO53TP
j1U1EGXgWp3hm104gjWSEfzZ7OblRei5kR25GeBZKWAZf8EO05Dvbj+orLTEbyQkUGSrBmblzPi0
4JKh3jyEJoQIedT5Oo7S8ZbnZyJGrhiXX74LTqCz0utJRppJhYDKUJjYKZDBB6AEwWrzph26MF23
5H2UvM+MrRSYyMmMeRNDgn6628k+WOMjIX9r3pB3WyRaDRHshIWE5a2dSC0w55klKghEro6sXLuc
zXPx92rTVwnjLJuUIKMSdsCPZot0jAv2R1Wh6DQiUMeILN9ql0dOnequ287KuScs8wnA1Jd9QDG5
eq7n41YrVDpBKPVvalE8f+N/MSv0gtWgSUgt6qCo6PcbXsYTLxL/G4OalNhicplO6NMRKUDMpqbu
k1i0vBUOx04efRh52/Hg+oz0lsy9faIzoPrmixnDl2/dlKd0VhZq9SnRY0za1mM06hiyVSCKZzBB
SauDhQjZQQEVWnqellQqy16ETaii97Kc5bWy9VpKOZQrlK4O5yD3DOXGb0WEyh6cXeJN8cP0UjO7
y0ZMFcqxqDtgJpscgK7F1jgy06pBy7KRtYTX+BBWwUvIYPY1s95wWlkUVg5+HIEwE3yBTq6LYEZ6
nNT2uXcU+t42qOh7leaa5DIVP+IdGluTtLex3jAVLIR3OTs3jYDTCwHtnAzhB+iGY1WxRSqzD2Ut
5lEFPc/4W18pgv2Qi0ZbCsQgl2qBRiP3SrEcCbnCmggl+NLSA9tX7c368iBiyCzlPohg31jnXIg1
3Pq2mh/ywv7uBkuGc86bHd48STeL4s6qKQBMVjGwiKjaSgukgUtNrhynO2esQB5cp4KdeGTI/WAA
uUrXGeRtLpN+UdU17Q2Uh1VEsNvUrnJL+0Dm9NzT4mDOx6i7//aJh+DYV/k0MgUFg3+vlAMVna3z
9buqG7RIHiVAXUs92iy5A/ZNE+a/4/MgV9CfFJ4kmRq6bgLFRB5xuJmEmU+lZvPLw/caOEEgkhAb
j8VPRRdhINmf4yGMJdF+p3u1QEF7NJXev1eSeq/f3XvvyXaLgAk9Gx7v0rRXkUwOGBxadgFslBC2
GrbUFvOh9t1+ey/QAfon64A9G0TKpzKVnKlIYOi6Nzoe9tT0LwTDyu2DO84BrIBX+ENYCbEYWoUM
x8pFZiJJ2tq02lsH8K8skJ2FiaqKEHJcvkp+4DK80uAl2C87LmTPPqEVojUKPNchGD8PccGSuTMJ
dljwLnKSzDQoi3P0NQg0iGrjEbxj5xeZObRrwfPBoIuz4WptLxgUh84Qf+ZTL6fLByLFxsbC77kZ
g2N9HTQ9/lk2igyHt5fgjJvNkoqg4jM45UOtx/r0I0eWB1I15iUsbL2cWL470Nm2gkW//1DHQm1J
ZosunfMvkVhvjTJRHMlXERfA/FcGTlhw6oqQSTrr7mha0x6HmIQhmsv1xuflgmc990968rMXJWY9
VGE1mF58s4olFyvziLlkNvUUr7uDhWe3tR6jtOn3HYAcTBvYFWjHmRs3s4PtSO5g2hi5yZ103peD
eLUxFy3x4Dk7KtvqVXXvezugQjDpDt+8haHMGgahDhBzxVkhUV9vyDhm5EUxmfEHsUwUA0pKdEo/
yz+iXvbWOGRaoNIFKjYCdI3dikx6xqj7Qja0XVO7q+/jovzVsFTBnDyK4tZ2XWKPVmGPpHe+cvxv
szH6twPR6sqT0bJ5mKigwExGviOUsTqw80VMy19gaZENYccgnX3AefK0T9qY7gg3aCwe+GIt8zdl
qf+yyreqY1GZddOmpP+5icf1CjSAmTb+bsa41PuOfVaWT6GSuVtUIgC0nHnhpffX6WxpqCtELwDv
CIDxICLPArawMOryb6wVTegqdVFxohFZLi6/de0rsu94qJV/1UqgxcVTkWrjWNQIZHpIaPtWOLxA
eOewfv+sfRi4iI6chZnx+hXxmjQSmS0sz175jvHaatrzT+e/erkC2upNngJjLmwMHj1n1qxTa4r9
nF76qkGe9qoBWPM6lTgwmuqe5eSGP3PJHH7CHidRIdew4CCPd+dINXQGEhixqVbGXvY+QDJSAmDb
p9I/mtTTP65sX5/kLodmyfhHRFeJxLfKIEBM95crpyo5sq2qCKr89M7OaR8jVtaPFONh/16rHJ8l
/kvimWWUFDzJ3LW8TXz0Zc8zlk5sOFuBKg6JVrRDdvafL9AIQADfwFXJH2exgjvJuxak+Q9im5Jd
/0Lpjv0S5H9IPB3SI+PhBJkmE7BJNPE1C/aOU1YRFy8vlyFKJZeoS3X8YHc2e8ZfnjkMo6x0M6fp
9HiZtYLPYOnAMK46DgO6+a6ia3F1yGY278yf1u+4cEMl7PGVL7PPQTjQn+ry3Ky515S/9h/s1IPx
Bb+iq9UYnTBP54KU2qJoeWJype9643X7wftK5fYJOsXSEBml0+WScIxtOKNyVITw5qqR7oEOlx25
IIEU8D1Q5nDkdAKLxg23PK4jKiVHo2sa2ukSCiW282qMllqWIqD4WVGaU2GqZ1bclHvanEx/AtR4
pefS+xbdpZkEg8JFtzYD5dkdDNGSut0loIXry3t61irSxxqzjdnQmsIpwQVUFNTGWXMXseRYyTtG
594RG/FSNc7Qg5JkD5klY4WpwxI/8/Xy6zK+VlvJIZLil2FDlY+nj+GzKfbYLxyc3zsQRuwOiPDn
6F+ItpbCbWtI4bfFAk/9AmuK3Oey/2dZiIMUQXJXLVWR1QMLl4QtjVXOdr3+heU8j3wY1pAL8ZE/
IKJyO2B0h2A22AAbfliq8yG1erDSYmEEw9fPlkY+TBashQLwCGsQ0rvjvZo7Kz158YDNhucgypVN
HQEvEpreCvwDa642a4xZblh1uMZdWeAiRrenoN227ehIBd8/S2ABYmq8O3UQuQZdgK54S168I2Zn
MeguLn19jRO7hGdTNKFCEveL2AWNzbquv8pZbuyOZAHK8vB/h7iDXtkkvVud1430Ey3B/uPZzS95
4S537foi2zxXRQtWEjsAAz4mAZ+ooYNu42PCtmvctyqlio+LVO65ebmPwMOghXnh2MEltagEK52t
VGHAZOGh/XBTkZWgSkpm4GDQGjKfm0sPN5YIw910wqEDTdBdkhn+PY2zGQD9BqH8nvOJxCAby+kO
crLJawppwDRpCsxyULf7Ho4Bd2FjXwUN7CBCYJ7oTIQFmOE+VNUSVWvBKGjBI4nRfMgQJ9P052xd
fbceHgfhd69Hce9j+ohLFUKzjwFVwfdWB3D08DKFiKNrJibpeVrjpY9kDjUP26rORY1IA+uutcwA
kJauDa6DAcP49UKF63QYkZBiVhYCr+QVVSinWS0Z6wZqiYMPZeBHEJTZyJK4kWuITCt3Eqhx8L7R
c75Sc58qYNyQLYANyUYTwGzdY17wU7lafsfyHFZpafixtJi6/9GcrO9eTJzQN5E83pJF5esThKuQ
dGppxnsOKxuBWAoO1suS/1fSSqvB0RpFAuPGAZGkxdoTjxrVdLU9MJyN0RymSj2gAMuzHCfC9KzT
G3+0UKbpbTlfkwlVqDgn0gFfYgJil23jl1virjl1GNpK/R75Zv4OyVlB0UeX68Ym9KARJPL+oW3K
iNsreLBpYZN1C8NU3CnClkx7lzbu6kAxfHM4086wZxxPOC0PPjw/BGK9eVeNvillPcwqTpaeuj1K
GkK9iP1umyDy3bYdWN3lyeXPMibqVzzvynoJxYLDZn808ARV50Se/aQGB46hW8hhUVEmBi4Du445
H9tj1H1OHXHUIndmLVNx4qb8B7+zoiA10g+HPgEzM64G2yVqOKCsh4RJjpntfIu7mQs+xv4vbF8t
glP8ZrOmbXyfJAZ4waHlSh74J6IAwJv0/yfWbwb/8k5BWK/vaXfmLx7AG8uQIi3mXEyNdLC54LoP
rEXyv7V7Z8SS+9QJfAgN/gGXytH9Y9207oVfXYXLTVdtrlGGh+SP7+nXNgr1UZPTUdKm3mKVE3CK
0sdVbidE0YZApI47+YoqxZjRbWi2fi8ZGTGpADuy0tR7WmnjYZWGEs3dPWK3c34M8B+jq7pxFHDc
0qE1dSm+UFxDSPS8Vn8yHxynlnBL+CVmbkZKZ9AbmJHMS8oxTWFg9T1MfkAuL7njBiZsA1PO5tfq
LeAO3M7BnOR5uPND4QyaZc7X7KHTVpvFuk8mJN/vdVQmPqqurY1phojkSKSKWwUPeyQCAo2lvOen
BpgRkY5Mv2Gc5jWYueHbYuQgvEKAaWzisiEVqcae3RzhjukUADY2JRWQEH37Mxz5QPiYGfMwvhe5
Jxw0Zndv7YH65dtLDWzz1l8sS3E+cAWLGHs8YKMW91TpSIA3BR6UByyg6489kJplBiqDaSMRc6GU
AaysD3tBN4hqm8excrFxs7H3ext5VLLPeEDPZ22FUFUcvmrhEwk4laxaiVPv/qmr2NQ7XrECvnI0
WYPmsvBKJC93jmyRtg4zgfk1jXk/wcbcrI7tFsYYjg30KFJd3duXxfMr16NXFo861m+ToOKSyemt
npkWf65WxXOxmN2gukhdMdhfjbJR6R7oNUbDhuNhfeCFdnWgIVbHEmWM5mIShQkpmUElaPWhiM+C
K2baUWWLahhV5oA2RDQEhGLePsAVXs0Ocezum+WxO+TKIVncNM4XGKNVoVsOc5NGoEEXaeh3sTdZ
i6LCc9GfqeBp1QpmfdSGmxdzlGhQ6wTQNBLbPAn3j6ngvE1FYU5tD3NxkwGdCjI+0Q+Ix030nHbB
55iV91Vvnu2Ef/yS03gH+lwuWGkKOdCOOcxsEoms+jqa/30W9By6MkLQcUfZ2Z0h8ZZjRYv/cXao
jTUYmFWwpPYFwKmBWxMwDdXSk+KjxxB241gTgThcQzVF5K1ZqE8LEfqSZ9lBBSYnG/7OERcQ/w9b
kwctLlIDB7AzpZKryhhfsTCo88jZh2CPjx3nc29oN+8VGTQDuxoVOpqYEReh/gtwroefevaeAcax
JX9WIQllPhl5xBczErBbGTOsrljUjQYg/uO/NuOUBUC0dD6GkQ1Ccu6WeLd8BBV4PKXzTzlhosKv
DCt3+2Y/HsdQudmVw3hnVHNWDnWQgyp0TC57oWL80TSPqKGsl7BEyamMtcpD6HKA9RUarHvygwUb
E+3GtfeO9GY4tF8ZIsYhpgUOvYvQBTCANDOnzUIdwoJMscjqiJ9W79vgU2hlubce7TxnGCa11UsA
zUs1AIcDWG0y9gRV+XyWRZZx3uRyyE4dZVN/Rq0WQ20pTLTC/LnXkcqtKohIqJt7Bahi11Lnoqch
VUX3aTprwJ0Lah1B7jOeMD98TvqyMB+RCSOul8wXMaWN2jfnV9uiO+iHX9tvwgSmiSWuL5CBfgGd
N8p5/4Mzk7JObe7e9YZni7/09m5J6zO6ZAfQAkSjpSnDlESgoQh8KP+FNa5AHm9eKDb7JixRMoPL
T33iB6Z53tB2SFbJydXMsBpHsC5TWcy4p+UoffTWKjMhv8WIO9xX4tkwp150WEbUimBvATwtuCRW
vWyIPsTnHp4w+OASryEcRs2mS3nqiJYBPiARggXyFU+/7Lhvq8lIoJVXzWwlbv5L2eT1kMTOYUYZ
7kafiAluOjATxgpswtEMQ19zDU4sNVp5wj4g//WtRF+e2iEyxHC0Uylj1zgm35fSa7v7kEPgamaM
oNDZqqqIdZDgBI5r7vtSKxRDZ8K5SZuq/bf9q5BMjp0m5LUP/xVq1SImlPo8U1+ee4pX2FBRJJJ6
EFpFzqmYB1V5XKWsVIu7SD70uHBGGoPf5/wQ0d0I3aPDJW+oM5Er7IoqryBdGSeOqmxeGMasyMo6
YanzTrmD20IbQD/FGl1pN9lpUliqeIIn155qo9LRjWGli9IEovWPP+CFxqMAzQzy9XfhmTFiFkXY
ncyN00Uvs3Tkl6RvHs7vrqPLSTub6wdsvZ9lkbmuimqfXuXmxJTjQeHnv0uhoZazuGxBhodwQCjP
U/chH+8kUmgQ260QaBBpWWOjIOEIuWNuJgJjGoa7J7XlacjYaIUopnpM2BrRAystGhZGHO+GBIzb
HiwInqb8umt2acy85HQrIU+3wlby5y2C9YGq6qzz/KvvRQOwR2BWEJm4BI8WvRdiJup9GwvjLO4O
6k7LbnGKn/A3LIdN6/Mr6ke+u01U6FuRkMSePLk3ocgvVYwiLWfPBeTjV/zF1OPQR8bWsCHqiJII
sQjj9X1jTIFW1GM0m429SfhMnV4SprtAyZBvNmowiTEJqXsP5CTX2mNVFgi/LoAkDrFZkAGm9rf4
maE80sJYdaWAvU0ZzdBcYDZOM8D92PZXiHlSEfCra1cgMYBNOGKllhiLSnutExd1yXr3DVtBW6M6
CRsxbY+N5ZGdjD4fr5r87x9AR3wM544srzbxe4Z7DcujRVYl152oEEUDW1FzUeuhqLgmlEQHSINs
IFrKhhvolxGDBiFvLFsFOoPYhsegm7pdt1Sw3GLIftpwIvi7DN0YvmIsWNjy830m7gI6wsKaj9xn
5Y5YlnTcstrJGt9ZYYWW9L0JiZV/ctbgwjfw52u3sQwsEH3YwM1Bi+a04hxhKaMToW8eRbD834E4
gr+105sX0TGosI/S2sP3mScvscwKGeurh3rifsjEXmpTw/FNmInjbFgsWNSGWFN1TTvWMFS4gIxg
oI0o7kig8NQ3pCVA9jsas27ufMbbsnWPuVjO2xB6Iy/CPLXZnZELJitkIpDCNcqLJssqT9toKOcN
eoOu/QXtis7+qlwPMfW+K9+kxsDVuDPmxs7A4t4DW63LaiTgI+7i7vxpW+fEy1ZfyM0JP+yLg+Xs
Mbsa61BEqn1DDDCNwIrnoicE9+wgy5ASHJ+kwPGViO712ifxUzrvdDbvujBD2ehKuIRan+KtUxz+
3AlRt8BIUoGC/qx4oj9bfEN7GfJBZmzCw2z7JZaCQ/H4EpFW5rxQGnEJNjsaQW7PYi0hPFFYWZtP
junE4IZ6yjD5MYvNbnCl4k6huTV2lfpKgvOPnKATdjCxWrdftzPiZs8yNRVow0aJx7Qf2G7CHmJa
K0n2H0+6I/c2++0l3xy5s6TVj+HR21VpTWNQz8C7bLX1eoAVG4/auJbUrNo/L5Mg7usXjnWV4lps
eC3wbYXm5sgmhMyouaZ6lFKFf01d3tbnFI7SGpyCSkDXxDV6WvWbVyKueAJZmQXW3mGmIhu4Ci2j
CbB+zvjkZzW81B8+zoEi9QR+kWHPX1vN9xxDOqUZ26fMHwZWfgOr3GuWjHw6HpEl0FKB8ARO+pEs
mNEKw26/bUDqgRWrZ56gSa1afibDxNjfY+JZNxdJ1fxklDn/mIPmMNMHUzn5brtFaADNpFF36rJO
Qa4OXWmdfp/sFwrzY8yncGFh99gpAWhROG+Tl7ZtIKFvRV6meT85JQSOiSXQfKOiCtT3dHhHJtDB
cPpxytN962FnKxkFSryeGsEZFedaDBsJ+kfEJjk9j4ezy1on8zf3qjh+n3e+y3NPYM/HMrxXt3g6
eYzfMMoXeT6PFjVtQl3WGWZlRqt8v2lb/VXFklZGzKIm3DWjWm2CxUj1NunZiy+c2Hv9acUHnROW
1nY5whfXok1sbMYyeA55Ft7aOYFXi+WQLRB6K1tgX8Ny2rrJLnILOySrF5+1M8yQ1ChaoSIJxebK
CilC0gS/XCP4bZU9CB19/IRHN3etrUhU8gt4rtmxrBlmPXd9FauNnGAZ6KBkXiLmcbyU++GDMf/m
uHyr84KbDmHCOuXtrJGaYHyTaNXOXf42ljKtr9PArrOpxUowsS564PmsF5hO4O7nj5VCSd78jgeA
h08Scz3c/jTua7ILqfiU1/gIuEn4keNFaayz0zMmcfHDvI5hl6LnsV5E9gCZKC2RgMPYSf9dD489
c0o9ieRkUHzFP3KCdGThDH5coqq5VtR61WqbH5WUi73p0UYWVgA7wqIe/2Q3HpTymlq13i4eCXK2
B1E3qVxS4/1bfYBr9pDgl/umE8tmL/w74iRwCtv8vxTtjhvKCVA1AKJ2q/OZgPOJckty2a+ei3na
REY3d4n+IzKXWdi0maI2zEiM6yyR4FI4SvMZ02GsE4Mb5YBQWjdamkPoJesn4a/n4p/HQFKXJQsL
9c7GhFBlpQfQz3XleXMV51MwqG/2ed/7VwIu2KIU8IGlamaTUVbK5sTg0KNqnSha/mRkPJzEguPh
deqMFe+u7VCNVradsKg25EuNw7r5J+CfCfKIF68NVA94FDOrOdWECxPOFYSTV84iczNbThtN5ToY
lwtYxyjWmIZgV+LNkIGq19+6uZBslklOvD+77wMOPsiXFnTntGynp0biGPmd0jOIw7WIdTT8N0pA
zKaC92JTqrmyISBr0FyW8iuSajU5I8+BB99ZiFwICBo9wRjNA4dMSvXw1wSZ0SeNcWKyhZdJ1EM2
k4u33+XgBdK9otwT5fN4E+YJCmczC3mRAzwOVvn4WLPa0oMd5qy2ZQ7qDSyy+9EFlsBa+8CXYibd
R3+4VU5DJExZVo/UwGBz//27z8QGsRgUnwEqS5oZDHnp6E9TouyjTUn44wALiyeGRkDUlsqGeeKC
jVBeiP7GZ/aNRglEdPx6wkx0VGxBiASTwelT90XAlCW/yXgKbmkyaYOSP95cfx8tp64AxlSDIuck
qFMRXQKaAznobQAWqYvyqc22Y4KLjIMB35jOyn+XQV7F6V/10hUElZmLurO6rqvbLXUEElIqjEn8
qgbtPfndc7PMSiOKw/IpvyBMSMNKaNpfq2rhJux7z6+/Xq0NisApMgxCoulqzYaXeHwU7M9nvHCL
UEZoOnm1JVJVSMvrvcmw6h3msp7SbNG+v8YehANkQMkxfi27zp26uS8gZ4+jzvb8COvyNJgxGqbT
J+IpJue7OEysiTy3HQvqhPToeBJgmgl9h5wX1AM96Vg8k0vzMkCCSaOdhYh8stkGzXNXA7w9hahN
7fxrdS6wlZ5J9tlWf6UyCrnImzeY7eTRXutSWG8q7QIwo6Hj8X20GEOTPU92Zaou+lGaM0fq5sIc
Xf0ZMW5PACrs+/k1xKWr9EfVIDO/zlQIKqFKgtbi0ArZGE4fW6L4MFL/2BFxM5JvfwJw0+9tv5Me
IzuGC3AQQDPpL6NOv349Jjk5tAITgZfFHppgmzzRhJBijeXPFiGxjIeXPOw/LbvdtLGpsU+tavEN
2yelAIhXDv/LCFtb1b3KYsru2XZtlLox+pSnexw5iFY5AbG3BFz9jVjJKWSIch7I8dcU+Siiae5u
KIZOU+SwxyddlKNfPjs3p8KhAYvIb4kp5urGKyCW9EeRUdfiA0ghgvffuj/6MQuTq79EUZfsjfej
LQuXvbQaiZdFcYTZpk4vcdfWeRUguUXXrkkHQN4fe+oZ5TpnMK9ChevDhVFzBHlGaDneox8R9YTf
WkyGOaDPJ+p4JTjENzj8sWc5cYaNGt5FzKGnO/hDpThmS/bWus/kepgF6ib5HbWomdWNDYr6UrhQ
k6lhd/mG8vHN+NaTlUAsHgxrBCOuuhqo6tbKSZzntido0s9lLFjIx+4vb3AVz/Pv6JJkeHJmCfuT
0l09ZefnKBnLhjFMsqQKJfKnN00VSnNs+KMp/5dcSnWyQyiYW03hKYN2lx0lUOehY1jn5YcaI6R+
zvAvdrvtdf4+/kXckNw60JSV3MoEdtLpMICGQNITbf5IpKaaPme86mB/l4/KzRlHGXx42RCu3sfs
up8mIBF7Bpma+KdrlWRc35nyjOEdpdZm+fbX9lXidB6M3BPDTW2QuGXcPGVWIoJNU2/rxGqCC1Ew
xTrUdDv++zVekB6vmNqOHUi2TBSRY6kqH6ZADKz4wOksioE9itpi8hi2dz67rObzezsKM+kpwrt/
qI3dZfFJu7YcRRQSRfZTMO51yo1w2t1c1inxinY6clVwtoPKsxzqIOJEzcsRgbZhRE9OjnXFFb9Y
bj6xtfk/jpMLKDZZvTny0Kg7D/htqc4UudeXv+vqzhQ33F0VprGrEdtNWETSYpM8LJy83bs7ovyY
Ns71jbPMUirlIsAlr5gkd2oLlIwaGzg+/I3EF8aZgomFTEp7FUV/PBbtmPg4vU6ntpRrrJcswqeR
wWmWpA7QtH0b80ZLO5rJCjBYGKYsTAZq5dmGfx4XRpkhIzXJAS1tdm6s8LDF2jvRDwzD9YCEC1bn
CGN2pDq5wi6bV+SZn7eStqpRIJtxEyijwYlaDF539ra9soUgtnFMzToh+nnzBOyb5D8qkCLDl+Q/
VJo1j4kSQKxQOjBwHGvi37g1UMFAEqqguroXEY0fPQA1VeXJ7LJd1Skk7sKY1ZYlRa/xH1VvR1Je
gU/XFa9rLs+y5KWiplLEdh2/z2Kk4TScjKwYCQINdjJ9/+MOATTVGXjW6S2r+XlV94+OPHCG7toY
T4szxp0iSRZmC0KdiWaOO2E4QECwd5t/gPjwRYErpTXx6PjWI4+hd/x/T72hLhrTHMAMWiGGzpXn
VmQYWzdFDoN6vyu7Cm4RCxZAZzTPDgZhv0q0yJEPDD5dXd9tR4u57l9gQmnzLiCIljDWlyH18z4o
5cXXINvmcRGx4xj05Pk+zafshjbkPFtFcoh0D1Us3MSt2MLqzKg/cfRozq1wUfQe+VrAlU450qcM
CASVoPWSxxdl+5KslihmdfyFs60JnwmQ3AgIwzH05civjKdN4aAmi2HLnvlw2xC2Ni+lx5l2769M
qeLDoVQdjlBFoK7XqTnDorSQ3rRlmGZmit236dB7CHkYW4Z+rQQQ0r5r3ZgJVix5/VivNz1v+Au9
EkCP9VD8Tqb+VZh09b51l9dakI43RhMHL1iz5A7XrWs9TsQbt70jr8Izz6okKghbxpJoPwU1KS9K
He16nLpZ+wQUb0YCVRDA1gLL+ZCcxWwOR/RhJCNIZFD8AgiuUfIMscSoYl4nykdJTxLfhu5Es9sM
R01KRMDVQdhXe+UMw5MY7ht85UdvladRrKL8uAzvL/aSBvL580xsFBv/rGbptXANmgCCmNTzemIY
jurFV9KZjq20sYe4lZaJXH9eb2VlNtoRDToCW4811NtmJrryn+Irn8x0z5tRVMMb2qs4dIbU9VeS
uBUw9BYYsoD4Ii5G4eUyvUEE9XQuIF8Cd85in9xT3pvJ5r0RUpVTbnsWnvlnKnRNRsUDnVbcl6rC
OGZs9hsFZ9pua2HIm6D2PjunbEghYf1IzhNRrGP4qyr5FBFML5Gd81j8SBZCDvtpzojYKOgJqMyL
Wea2pH3uECzkUe7/zYrBaaGH63IQS4uhAuzE85MtWOG5+MnJXDWXBnQrXf35iouyiSR/tW/A+iSK
rc9GmuOujTOxviPadjL8AGnLchpK8YPj+BsnhANqYlHDuLmRlvkscNl5mXFV0+M9chgGp7pkbHcw
mfpPrzC0X1H5I+pt4u/gfhInvBJX1dGadyxFFU6deJ1gLSpDBz2EY1i0yWI9IW5DlLOk9cqy45Mj
OiNsMlfOoQjwAdMjy91n5gYGHDr730ghKv04l7YFH0p/RJhNksfpSyYydMgruZOfv4/9IVHqtBxT
Xbe9ii3w3CdZHJo2SfvYn/GW/h7P/WOXEdzvBZfy9nuCX7Zbk+YHr/Kyu+fKvXBNz61dvWENfXXR
CCoQPVqApdenkzfpd4ImcVo0krPV1W/5zt+ggIJ9E2dIGasmbOW0LjfQ/nNrdme14v629ZSnQyK3
a5d1VRmG/aNuLDG/ZO0qnjOfe7juu4Whakj1TIWT0A7xJ0xPrdHFK7ODMqcX/kl2z/CHgPadYVLG
bevftyAxrGClC3qeZiRziEzYyGkGDynGlL6m6MZQpFZz72CEgpPgjhxP7a+Utf54UpR1H+9rGBfE
8IlTKL3UGgwJ/0olRMFDmeDD+Y+0V9dkvWe6qAvBvuUzMPGUS4QI3paB+NgGHbub2/W7QjyHy9Mf
YQgj41IwK03T5z8z5Wcb4B8sGeMkQIyqRi9MTRqiGhYE8Rl4O4mUJ0k79JL7aPsWDjBsaCiymgoV
jxn9acUtcg7w37a555A8uikuVdw65xwStF9m6Ve0bDunbMFWNlePimAh69tTdu39xnPYvYkpINYE
wbFSpSijXZsk3bNDJZqdNkvKtUD0xgvxxwNP5YmIIGNCPKd5QEh53SPgdq/zxQgXXaEmRMaGo24m
cO5mw8s7N4I2h+MOHMhRtQF/4Q05um3lH+L5H/9CYjf3pdK9wHEBqwJkQqOAG6Olg+/zG9fbzIkB
v/1z0eV8niz+GytD70+UmbaTO0SF5ggZBnZOrg+drWHe0eJu0F9hDkP+0d++ekYrdpLMS4peLoLU
QsK8mUePCRQZv3qEwj8PuUYxIbnVrsIPh81qdfCkr+EERmFg1HSfHUKlmzhP2YyI8+5MajkS7RR7
gLMLRfo8157WKAJQbhbrCLJEOpmjZKMwS1gBGHcdkhKFufG38AODdWbfH5WQpBUdt8GCSibb/9ZY
d7WvcfQ8gji8Ac/b2b4/6YTXfUrHuRtDKAydxCLhaF1YUp9cKwS1cUx63axHA8K+YkFMSN3Wmi+u
D7sxWnjZ3DHUNPcBXjY4xUs5020XcKV1nBECndFlrNnGl2dZLhFK6bBM0NOXknDBoThcCQNGuIac
aef9p3oVRqVqTwe6BABBi/iwNyRFcgLhFaBLuHBeoTp4s92QfEpzYQWcniR366IgIN7Mzydbz/2+
JaO+wSuKIDIt2vflg/pxIG3MObEh6Py44ButEbGevP3x6xql0ZCsd2+8dPHz4cJ2F+FOAWXRllB1
/O1VQkPRJBuaCYZthlfCOERn7rIvPwyPp4hzYZ5IOun2ZMF01jqy7nvQMT+Z789An3CK1BPrSoaL
rWI65TbiCO1WXHp78nfK9BDsnTqrFQ1PuehiZxcVL9el5A6P+oGTNoYQ6kuUtqA8k2orck5F5dTp
Hys9/I/ltcuDB/kaTy6EOu9aNI8w7sxmtbMlpInctcAC0cau0PE0psVYHfsIYitvAWVc2N7XzOXY
aguQr43qmz3Y4Zr+XsadBpbc0Rao+N9IA3IUTpJyxEgbZNkA9c0EiGHqQmmqpSzcQyT7cDfZ8STY
4GoGbNFDCqZlB4XgExQdhw4lwf9RbxxWIgwTDl8hQjr0TBtjlhYIETmZ/XYaIOHfYWzPbtNaiyyp
e6RStmogGJacfKQwqkM3GNYYezcG5uV7ZoOeKNAXZZtCI0z97TUy3wIn1pU8ioVqyoZHakpPwnC9
/PCU6h10u+K2HlU03Mgczxc2jBmpm8MZOUN/e0evSxYn5T31upC/JkG160jTlYfwHfgb/MeHvpQo
7mIa9r/eFNH+M09krF9cv3moDD/xa05R914QSd4kotThMPipIk7S76FduAoKLHieI5q2b7APY2wW
iq6GvPY3XB//OEXUWQIbaoc5zof8D1iMIDWrHQY8U1fWdsoFki6VD/Onlhho9FOlvkjpCNw7f+Ya
fjo/OIiwlr+Kd/5r5MkaZCx4efpOl5It+gJ5KZWmJDlfCFux1epMrYbQ3hy3WJ4V3zzypnBZ1oI9
ZgvFV3SknUlp0EXPqMSh4vDBYuwEsAbiRvc+5LJy3vMpde3FwLsuZio6Ikt7yGSmSHxHnWFYTY2F
BqDCZK7E44gJBl103zwcSEb8UarOdYzgO4eTKmZR4msu9bACtv4kr7cQG/ETQe2XdnJRNgOxiQd0
6cclnXrPNAAhyMVP8NfLL4cEW7FIGmzUhIU23Ap7YLbe56Ub0r/FI1BjxVCnuJKZ3pti/9UOcmBn
IkDKTAnEgSoIp0hAfdmwjhEsxWAhxbmjeb9fHh+bzDCueljv8UgeX2+VB++jUs8nJVqxf47e0gzN
nyTjqx/D+w0B7fFgag6HTylNPMlIBJyLnoikP6J/l5YxbjTXRJ7fEoOJ210Na2f3XrEOf0zq2M++
Tg9eRHG3gML57DmjT/mlM2+pJDr++2T8oCso7uld2rBU7/QhpXxLPT/cL75xWZfDZQfg3h9JpCxt
3WpnTuETT/t/Atj5ZPWj8P8MoWsEYDBOCb9W9PZvZStDKNBRfYDqJM8lfPBmNxFeMVmFsB/ydg+0
MMnoatXKcIn0AO8Ap5OzQiBkvZ0P9C7CowSz15udZNbLLXPDonb61FmBigH6qI2XcTy34KcJzspk
MsZ3YaE2jyViot2V3sj4A1Ge4brXipETEPy+bWYyOH+BNuiN35/J1P7GM4/NnYgemoeuEN+V+GeW
/L5FVE7ZAL+L+xHERDtE/wTaEa3PJHTkqN3py7B9hbfxL7/79vXmD46j9CXXPdTP0pBMhIXBucTA
N6+sQq+A9Kvt77C/h1HV66mUYqHffYZQFkjaI9cGcZ6yvQz6yJSoxqMUbwrGqzuQWg+G5KBe6D/A
WJJGT0d4V2hvchtnz5KVPMuJMjkKeci39f+7+OikR3g5GFkBiVjGX5okKYvS1/VTrnATzUP+oviZ
IMzUlcxvhKjQ++ScGGeKIbb2eGvhdFUou+/VA+WJlCq1eOlYuV1uNgZI8+QM3xtZZgWs5f0mBEYp
/PXtgkDaiGVyJqHJtExT6HddYHOZpdjKBxWF3chzMj3uyWvjXJlQyo9NmiSvtCfu4bqQS9DLrO0X
V3z5C3rC8g+BWv0SOVj8EWNlQ3SU3AY8lZ/L7eLA2gRMwPWcvsS1NR3vyIoo4vDzVO64ExhOnX7u
Wki+QxFFj1vQzhJ8k8x4zN8Muhu8GqN49NYfEISZuaYYl19jjNSyw/08t/VNL8NbLALPRlsMr6km
QUuX9x3g3un3CpPKPyKzzHiZ0waEBvBCuwT2R/2jZvlKoQd2hhVuqTUXAPZqS7f8gqj2rGRTjc7a
UWP6l6sveVmrq/TAKuQFFYTO2ciZUSKJu6NYYGjPO6rnryPXWfA3zfZLTeE26TCX4cElgj+9acs9
vlH2d8W5DeNLHBi3EV5ot1jf24JjomDuX21qcOHHWkVV9Owc7aoZExPuIwu1C52vWkEr5UDwOtSq
6g/kb0UMfxV9P445UQeh793BN3Q/KZfu4ZEYKoXM/tP+R3DxrTmhfsbQYn8Mpd++CRdBeBXrgYO9
4qAboNeVXZ3HgzlIQH7Zze08UQXHolLEPzVU6fddxB/Pp3Yt7RyajbuOvbzsmI4k3lvu2KSBzlvs
DnI/AtXsMHBnbz/K0M8ccxUvMlhl2MPQ7jprtFD935e884bvxzjtgrIbH8SJeVt3rslw/LMPRoTd
mWSPoyG/Ff0J+7OpFnKohyIETYTtCegpdZlmUVql1g2hzY/OelhrqnXWh6ujeaDXjclXM9xpevqB
OpjIlFgPSUJgnJve7gPVBQdai9FQsFeU54W/tKA1m1/FZxORf+Z+PVDq3U++5dTXUoAqTjPecVw8
Sm811jYXJNnqRKN3nghyOtc2RHGvPzYS8VpQQl7ExnZ+ozqvhLGDckzSqZz4jSGM4d7FNY0uyxgq
SFyXQzuYHFg+EsX7YpZMg9OKzH0PUd+8lfnyBnrZkPCiv+FeWi1rUmvHyhTh4OalnJVuZGkJ3KNH
8CIwKobc8vdccRuaxHIrSGb4UukEjA+KS2gC7sRZmz1gfNSkAxJb/5dKeyAggC65M8V5K6Wt3yQZ
3k65wWUd5+zuJFwktNUHCSxkHnOgRIecfH+zSIArEb+OmruiFWQ88h2caeeFlaRvOhLmxPJmXPIv
9F01o1tVEVftTlTlZpaVSKCwPvqsO6esNgQ8BMamtWP+i/GFHCm/y3iOzL7Cd4u0x2Uskf4Egx2u
nz3ArNy9NVpgoJkEZmLb/Rvf9KUaJY7daYYAWal7/9i797gxCpbB5ANbFvlq1ky0WJhJomYXTQSa
Qb+kuDmNUVg7WTpfVP0MecSeQ2mHulK2GocdiH7qKW7Nhl166XRKLECR5qOiJPfbiZRyt0FQgzVy
0rH51mDaaPImAJkA1keNlpRgUyx4CU/xl6UxvRy8/OUHB4S3BbQjgRW77fuAZsS/PrA0LzExi1ve
o07JWyJed5saGtbPAydN7MQMg2Ogxe2WYeMWRgOaBVQuxN4VrKe46Sq+KvAQWftIiaIavjfmWczN
ftL+nsuN8Wt2ggVRihujcOIsn/kXhdH6ikGgL4dLxEUARBlcZ5VBiD+eZxO9xBQFx5rBHUJRkYED
r6iC/wvmTTMFDrsmX0aBj5jz+aMPuphzlNoNBkLRcXtlxUg2QXY7zCTbZH5ZvgHBRRFHg6lIoKLD
6AtI1+v5l4kPEKzDnMRQf5gGZZdRJZ++7zr2Zk6tSSh0OmwIw+IzT0wjeF9CoJBriuQ149A4K4Ya
g7AtAUuoJSoSCJ6KUr0w9xYQPnZBZV0eGSAqalUkCAhPSKCCNvulwaoTRShGyK7NhotOECQ+lNb4
I5TVjyGru8uXjv+ndC/MhERPrBz8ag9+CSF4okfKn7wtbh+YFhVKiALejTRe5mizIIeJkQXJg2kl
bhzcjQzcvDuRRfUdGVM+x0dirJHzspHdN3ydk2r6oEIptmZThFp3ZLbul98vCf4zquw9bAMkVacj
kSBcBDSGlRxz0gezqe4zxnaoOJ2dFig9qxL2DmVFVdJj7w9JYO3f9TQtRKUXWFbIV5pk9lHwq6Ek
s8T2WOGnTwyCmxp8iod/lhH0g8YZdSfwh/2DMJdc8KGfD4Wo40VlYclVzXDtXNVAypLZGliOOdnW
SVHukrtindbh2x+MV7I+xeeEurupdzoaykV+uQ4P5EHInrHQyvuAj3soK75IJUwBjQDPcRRqHxzB
qEr7X3Qo4Ue2Mi+Pgf0jvtqCc2R8EfQfrkx3E6Q+IGJ0rfze1vpLjFjJdI6aUsbo0VZMXyXlJ6Yw
g8/kLn+g52Y4k6H4JImAwOL/7cxTRKb6hflJSjOm+gcgJqDX5OQABPci5r0UP447QrgIw/4YLYnx
cMWScB2PDI0yPk4QSb8OBy+U52dA6NKBihdpduyW6iUi2Wtv1PiyEwdMk1FCITDCmQ3ot40qlUeu
y0WhdyfuwriUXCZV8FHJ9lfFBPKh3U1B0+0ktSgx7PsqMwImZElqTEKnt2xCw415vqxedu6XvLm1
dlFoswCYmoRsr3nKwLnlMKkgR1HaJXF+TCFr0xVhHD/Z0eBnVJ4JgKzNYCxTxgi+wErge0nBM/Xf
+LiUU834BqXCKod7rrCIs1StwANXvsIwni0MWSkQNhLBOtqHJRfmlSKDQ3yeBEfiJc14PSROHQdD
h29lp1vOO104Lt/qSHuKhgMbtn9mxpqHkyLaaCN8OcVmwEagVN/vFLzpb0bUK0tlhxFjJqCQCNJx
FHaAIYwhOfrOUhmvjauYR+MsUmmnm2qGBrVImiDQ5QC/3TIHFpQjukpkwDsR489W4u3pJYDH7VfV
zNUp731Xkki0MziSV+gvvpjNVzaI3kP44TSG/PiySv4Cv5tC8se7+KmWaa78Jm0MvDbVwl0/MQQl
+9hw6XOqS54WmJW7Ztg1jSs3ol1GKDrhmRFkU2usbp4LFKM+A6L2af/CeKvrm09BrAq3qZlbp6Rj
iO0DK8n/VHecuFz/7JjCp3aLdW6ygzUCoP0fqJbm9jHGG1vD3ODgfdf77Pldm8WXR5D182SELN4r
F19BA8Op3zYiKNy9R1P3ARwPvH5KrHOEqQaf7VEWIX3rx8I1S480KxY16IZ1UsN1vhC4nyC4Oo3E
6IGZR2mbAaQmLkS5kgBoAVu3H6hEMnRHKT168a78cM8T3P+hf+et7yAqQx5alIeLn0fxSY6gPU20
eGZOyZwoLQzfCPRc8b8GI3gX0Wbj0SMkMCNdxPKgde/QCgrpyuY/DCCjatMCfpd+CRFrXkmpaWCk
mSmELZWiQoz7rpnKsmc0bILqHv+qfSDPLaGxerCDyjbcjFl4F59hxyy9vJeSyrA9REjruh8dMzp4
EVR//gJsj8P2YylDTDk7xt6i1ozy2DNoZ6WgL4il9yVjDq7Wxh1+ZRQWGZqC13dZkuJaCbBppVP0
MSI8iULPlYHuoJyMFLCI2U3IjsbJlreGcLkgzgGdQb3fe/SI3xzUIE8n6Fewe3R5llThcOGX2uF/
XSIksyqqZDhE77AW4iV5LseEmCt4kNdU4xOm9yM8yBWiVGBOxmGy7X0kSP0fkhtZRdQPRAaz1ZhR
lzqDMPLC1dU7NLh55AhQmzN+zZy32+WPLp63xuPk3/oPCng0K3r4X/JdZ9UNHmjExZ/qo/imP31L
hphaj/fhWm6bUIAioyufo00ASMgvSxVvSrl0cLWnCo6goR/QTR/1S0wDxeuYTOY8WVsxxoL4JaW7
PpKFZFRCDFfEW/oy8+KHii3jMZ06xj38o+DasOe6ziRgIMo8S3slMqHKs+LCzyjLqZ60l5B5Y4l4
NXXwdXI2NWdDAH+KDmaJuGTxCAb+SHOVprGfbg6OEqVlIzADATnROpaAMVKW+gdLuQ+P9jZzn18n
AZlPLfX70CR9Pj+lZ4JceKfYIyINGPusGKKkNsKxAeK0GwGOBpakzcqkmQpW5wnVpCjsXnMXvh+C
s5rBCxDYIuGFYgOSJ1BFFBNgAxyz+BUYARClIYDZNg1fgIavcXajuPjwmt7VrBDit7TDIsZMUz+m
Mv5WXks8yTA1IpB5St2Ue9Gh7wyh18KUwT43kfQDaKmO5n9tnsxMjgdtqLmd19Np61J4t39dtamh
Gi08oQZm+lHePFx4CaeKXxOIDmmkp/tY4A4iooS20iajX7xbv5UXWKeTN6nw1JrsyzyyM1Yr7H8N
tQCceyz0oEPrbRG6G3Ve8HpE+1yHh7yxvfD6Q+SXb/q8BRFRuzpwx8VifBAy6hftm9SsrIXuw1D4
btvzK8DBbJFyYu1cciZxoQloEl7YgWtmE6FBh7NL1JozoxIK/oE7LvBAxzI0u9rffq7q1i0xhejs
TskKMYe6qzz5OK/0M6npJxrjg8/0cwxa35UCbud96gvGYPrfkFpwGHBPBZLgQ3pmVi0P1lA2KAg9
kIdMMnza9xJZ/RwHsPEoYNv/1ZYckpBCKi75Owr8kcNlYeTp28hWsxjMG/ihPmUEk0JVPwHs3cAX
Zzv59J3xUTCFfTXN6NSmDLRlNUZwTQ1e/19hVxWS++bxV6UJQWUJPazTJWzVa9SR33P+4GzinTx8
TpVpJaKV2CVJXLMech8AbOILNtdA9QVAK1cHig50IGDbsXdeHCALAKd739FSfJv36SLtyWpSt+mC
1GZF/GUu7xwIII+sSQJbBWKrDvK80psT5g6NeBwSuLTHop3ZLl+sceFjJ8O4IYXLFLVQXC6hQ9dO
Dt/uJNOyUCK/0zuZ3osES4pc3AyKx5/6UqJOwNP9m9Ul6Y6LuYovLDBwrrpQ9NVtCzixsIDIUcd5
DmgbjtnL3brVjPS4j4fkhJsoQskfrT9dknM107mzrESyRCV6aKV0TNeFXcXRmVKfPLW9CGEknYtz
j1Hdzn4iMQqzjAgbyOGiE0JwhOyDOAvmQP9Mu3vJlVOh5Nag/k0wGQsc9GhYSH2ho2F8N7zdboUP
pJornkcl4FM6BrJ4tZ+BW9Hn79QtvchxAoj45GHDS0iHXc/qVD9AvKMnzq6LJvYejebr8mWnq/L4
Cc97KVST1jVsoGKhVUtIzJREuXZvn+H1vpl1kPxbBO2WaYK/0kimCkeYCVhQOEveu8GZh/01jPc0
zyd3ESXoFgcm0HdOadBbtiAbiitwQ+F0QpioKPExogIigDeScU5dXSdKRmmQzN+oGQxQfUobRGlW
zrYYLT5eNbOXi4BhEC+hpMeX8yWD95mk+42QHQ+qvW7Pr+r9Teqxo0Ci7SHCWroobzb1rU/rHKuR
lM75SqrEU1OHbvBlocqD6oJBOtKiw7FJauMXDNOylM55UUfbs240irYyaF9KY2P69GIKCi9UGoW0
ggoqCOIRGEPmC3phSHv6E4fndrcJzQKAppXp7pooXBnunWkUop83gMrOSsUACZnIoj9/iz3wdkO+
jD8V7VEa2lLcYcd0FreEZrXKYBgihRF16sSJ4GjvN324r8YMDcn8md7FCJqcACJYpC6bk9l7S8mT
31usupYUA/lnC9KXRg9Qm50IBhYZmCnOeV9VdqvcSMBF7Mi/5V99iIhJb+VZwa4yL55jX6ARbAp/
PLCDhz9XyIUwQqVfYWIyk1Iwag3Da+Cmu41pnbYAoQ8BwMdD50O/8e70lyz/Jm9jN9XcDCSrz566
97ezaBkdvGUAstDRUpdn1D3zu+uO2DkiwO+WcM6n7NuAKmx/uYF21XMKan0Pkm6qFNSm5iv6GreT
1ZrFFhkSH6KEU5hlaeAMgzA1RIw3E+6yZCzU9ktaMDEcdz5jQevrUIS3aTkvjaBm6guG+2i6qfNC
6y9f6cEuIrVVmlHRBd5UPNycf14lBsTtXSnTdeLq8vj1jUYdezbj2UExhOk5qodQVmz2t65MxEnn
EcBxSHyZ3mL2JlIzzD/07DDiob/GVEbXw4UeYWJxaJHdHXv9hBGGqs9bQvcgtD0YCH3mVHDkhsx2
TUD7pyRcMbWvpyFpMBideLAHV7fZp0MbkaCtJ04gA/uFjWRXrmg65p8jGtuiZ1MJTkePafWBU/A/
EjqoGHgJxPe1lv/V2THlwzMJCf70vLDtCYe+5JBHalMiCv/wISfmBcEHErxJyBgdbhVyAwZyfkTh
fKhu8Dwr/oCUEE3Pyy7kaW0Zf74UDHx5SfnCLj1a5u6udccznJL5flIuuvdYZx15beteCgbGDv4/
J4kHQrBT/JmQJE/D4wJZUGxgPWxGTH+keqJh69+YfsS/XcxHJGK/KLDBksNcbSCiImOubmfhs966
PJxx7CBdfOn6CMV5Z9RAi5McMjLU2cSxB3ueSEsFD4MtCUQIlO73rzPSOjab6zfeWMNY++WHG/Oh
3bLh9llieG4ztqekQV5fjI+rQI0sNfr2UDkemQi9BikuEBEsm+3f6aUBuot72zGhwP4x5tPtGBhU
zOmIGtQGPXZSpe5JwKLsJd9F07S7ilEZ2DF3FUa6uefkomtW7t4JQ2CIN5Lw/fiHbsp5y0ZqLrtL
bJABLahK7oUcvXfmJq+jnzIYyWiukjhm79mRWRaNVU1zFHASFj3Fqqlluas026OVA8TCnrgSk81E
yFEaYfxZnXFYv857Sp5eehHLyyAPGKyoaOziYjCk4mKCMyc9YXB8+JiV+SYCwB6kOrbAujVulTW1
k87zc63tixOSDHH6ER2hWTbN6CUpIiRMq634CzisaqPMC9cfJMcU56QB9R/y2jCVJC7DLGFgty1H
J5Z2O9ouWvQ8MsgX3Kz7b0bA5MDYx06O0lVdcZV0UKErpqrRnAqGnQ3h2CXUoUML+2WZwdfSj0G3
VNHbSw95+hs/UD9Lf8vy/Epv/2JS0HVKtPzaLJirmeDMANHMXek3AEKfglYIoyiIdhaDlw7YU6nX
NjxFpB86hoSNgVX/jEP028XET5JLk5kHE4cMR9UVYkWtS+sfmomvDwpBih6Ebx8WZlpD7g3pvpZU
LlbnDS1sLpRRU4fPqxLW/9KVU+AHA2mr54GvAQxi932P8J8pWBsqlv8huXh8098UNyKUyQIfejsl
UanBi1m0GE6ydDs2sNI32Vl1Cdmk1f5qDT4ERVBnsVqD4Zuo6dUurmfOSbZTvTZ3ahl6MdB9VKfz
p+XCQer6Iho/O8rf82oSVrC5dfk1Xko3G0oTKc7unDpHLqR8Qkif3xX84uBvcH3Um42GxXvPHNbq
MvpPCMeowUBZ8e9uc5t3RvYUX9ihmcS1uvbAwvdpsRzbHj/DIOhWlOiAgSKV9tmJG9UvfZOQRNH4
bRvATgq98Emu3b1MEebAx/IfnA8g9GJDX/qbnKiAdSiS721MTu6c6HSlHdZPJFZibt4ZdQHr0ndK
zboMF85MzXz7sOwI2GdpQU2nmvUnpOz1WH7uawW6XcuY3mSiAcJgJNpXwyI028O2DpQ96PGGyaK1
dL0CnchEtRXjRTwoP1N7kZwGzMym97IyICYKWDKgjfzEtveuI/gO9+H7hGQfXs0trSyO2TbR7Bcm
l85aUetqox1zRqfyz+Dp+ARnkDUhKoHGhocF3VDkQ100YnlNyIQjku8SGuc0qDiD4TeaY7V7/CJg
CIceGjeWxQXJiuNcGWwKIoxiH+jTKkl/kdlCrb7Lsuo4IPks0CoGNurqFploy4jTppuwvF5ilyyq
kJWT52BaAZSLDunBW8/zQOtfaWyN/5PStu9WHRvQiFlPNkWBeddv+BeDosoHNYoZId9Pg8Y90+Bl
uxG3vhgZ3nzdAKmB6B1/7La/IUbtz5xW06T4gPSsiQT/lk5PEP3T2fviWBI7AhlBe+o2yIQQ+dY4
SW4JFclMWHW11Z9+nHjiPipGh+oEimAjIe1gU9DTWUbkFNdozVHYTN9gW3cV+O1MSPmymE1/CX6j
EM8m1v634tpeHvHfntvQCs2W8oDhK0ZwvVhOlHRYJ4xGq6zOTcK1/NZWKCTWd8df9WBuZzqaTEYF
4EdtjFA9UM6QW9dsEyxUWj+71zTFdKMvZzove3ZYEPsO75Mq4i37es/gwoBvq9LN4fx+Wui4xNYq
sQD89O7zKoufVN339mxQKASuRZYM5t489FMJsCinrd3DYltx27o3xo3DrTO0IkeemwVcggPFaQgW
vjZuCu9XHJMycnMSEod7FZ9viMEX1K2JEQJoCp1tU/6ZlPM8iCl5ZlnJv4+1345VRTqP0Kf0uDVq
kt5NAo4YdMNPdr5cZ+6VflYXP+LEkzC9HNq4tFbXfxWwFwc0A+Kw0uvgKjEgYnCSEuUIR2fT8nH+
aO16LHB8LlwfqjhgnCiyaWrveGbAyG60l30/GkEw4wm4x/AWaAsOlUgVyf3hwa1iSf5QTZvRjTY8
utOn0rcxsIqablgAmNJ3HWkKP0wV28LlFAxM5eA51WXx/yvOaRe8CPzL7B5w+dFvvRNCZFW9w3Y3
qrBKKXF7YbrN+VV6hCZWPF4/drM+pTM3NHrXbAo8rXpqVfPNdkWfOmX+5PbcyuqAd1aiRUqE0wDG
dyCr/nKc2EJOBjUIeELQnAoKYCFg59kz2dl0dUhG6p4+lq3MDlnhrdTgpuuZEwgoD2w4yiI+f9sV
D2fJ+yub3TUV70Rmlbn6QZ3bcms/EtWtvNWRgVpHEb3w2GCmcAX0bLjR5BKnODAyh/jlOtVDFPyk
B3xL0yucpqcgPSe00SFy8ut4fu/iiWoV5pgnuK9Goh2EVNNx6o4sVCFBuM3QhcQ/j5mDH2Qll6wG
wq8ejqZa2+zPrvZtFGOZF7GVWERrD+Xa8x6uESdexZQlcCFbbNw/HjPlUfROV9W5xKuCLJXxSLXY
G0bCTh7fxJjfhoy4pm57nLXfN67cDoCg6otfnvFyamTXEHg4rZxKAZZaTd/AaKcfgw3QLQcYxJY/
rsgEE3yzjBlsFFKA7CpAZ4lX9epLCkXxPu9fC91husVi69wE+RF1grynNgj43Qy/OIRmf4mD8FOq
jjJOUSP5CKoMmqBuizC8BBS6m2GHeciI7rWuqWN/rwnsBcfl3FgvxrbCC4vtaVqM5A2A0FEBvl0u
t8sIWxZ+GQREqAuzbznhC/AfkDHckwkKg43uzrofHk3FrB9maQHqabRaJFMrDdb8g/JK6nfEy706
We3p6PcNw1nK9sRTTNvImMDfe0TTWhKdakp5YKNExFnPF3QSsDqm9kCU9Vxp4vnV/h9hn4dF0m0U
9I4UTk76rPbirmMm4s4zA/IsJ22vvbZZu1yDyOdPO8qUA3+80rezXzJpK/eIKjTmGauSgNBW/OE4
idyEqCd6Ur/NAp1eGaGGGOcRUZMTD8OChjpK3wARJJbuXb7JtHFExPHdlGCDq27tPvAq6pnZ81Hu
SvTr5RqLLi2zCRwdrGhPrlwjDnnNKoV4HDc5KwKSIWZrH8bmdgbnQxeAYKry2ooSjsYd+1tgqVzd
DeOiVx9n9kSBAV/vH4DaOxQZ91Z31ktLpr1yoSo6xheH3SBu0yMRyRu9jlYdJyiukinb9gVgUTYd
80i8kHw83UXJAasSUCWJsRrLp0pByTs+FG+K9jxLQKXu4hdcdKkQqo66+EA9aaMWj5rgN+cy2vnS
5UjSs7+nW2zB6058gLuSZSoopqs9MpQXlLsCJmkV7w/qcohio1y79ej5qwDHqSHG0leuQjGHbn8b
98PKB5hrpkTqm97kZATlJIdIgt6lzyVKTw9OfgWGPQf/OHL8Xlw55r/kVUXrFpEeJuBvQvQGIIfm
evnElq+UDJeJV1W8CWzvq6uenuvGfwCBul0fjtu8CaCvCDM4zBc7spG+1VNttRFwiX+1rgXeuJW2
xymvij/vsiq8dbcWMOO+8OrTvIRNvGyJtGUHdMOqTQn9O+udZ9cm/qC3eMpL6VOdz5A5a6kNAAGl
ouHxb7cjh42NIvCFVHDczqceRwUfb3cNHdnGxxPdZI/nXHQDWtWFwkhO7SL6pC19EV/xHj02HM6M
4qw1kUhQ+og4zCdYHu6ibkN2pu7IuF3WwW1PCuwAsUjK9o4o2+sTIsCWdc9jnDHlLqB9GHLhsoru
XBiT8dALSawFOuwbkNZpRLbFFEwlmZotGxr/JXbgBE8SSUa6JeFMQs/rbpeeBjGjhDc7np1FJzl/
d29QMC75+8mqIDrkPO56hJ5O4HuAV/nC5bRN7JD7BVluvIGVPGxzQcc1bMd6+Y138Dz0P2dNQqnm
PNHsyi40V6w1u/HLK5FbwyG8o8O4z0uIS4npFijUUvDI4PSUYILfONdaJu+3Fe7dgIbAcJmHu7cH
to7IhUQ98WSJHhZjyOvEi8PbRK0xZgawK5QOu51iuTs9pXuGXT9n5pQVq/BXTgDfX3uiJLldHhRc
+VCrzcOps68hROBNY9mHPTy7/Cqs4Vxdo564r0jWwtJdYxM6Kmq0tM04JGE6LQ1fF1ocfTccBpMn
8IAlx4wn5jGiXk2nO0StI29EaSF7jsKABvWfxmTEKrA+AoTL5z/0jI9RXzN0AjnnYziSW2sN52o6
526ed+bVWu3+eGA0zDuA2kOQ8crUQoKC6NccbWv2n2cIIjaxOhCSbiwgtnkHgZldEGyABI2kzkvm
NNQu4foAZF0ipF5UUdOQSzDbuv2+1uqz88KhKcFUFP9Sc9v86F9lLC6cVc8a0dab7emuIhZvp80t
TvoU2spkvhN7Z9rdhzNpnfKB5wagC6xXHPWagb1AdBfaSI3iLnOT3TEriVCrG1pW4kt3reOaT2D6
/vrJK1j8cfv9+r2Dg0BcmcfdAL1STmLVjw28D2ZsS+w1ZIKNiGEdIMCvPwezaDj922CNb1O0vsjO
I7+vPiQtULb+7HYveqs5pG3ZQvrRCxeqSebfluc3aJNgSV9Mm54/Rt3zjxAjmHTTWxnXC4pLDTrS
O++4m95z9eCEG68v9r/yYDN6KMMRbZ5JfPcyW5sW+ckZp1IUywksNvigLA8uIfGr9p8pdInnh7F1
iIdM/f6jmaXNrX1227W1Z4PwGMrtJJhbi7XHKKFW/lD6Ow69MW1fbQ2k9fbpzUTWpqdmdtdfCXG1
8vkiwLxWJ6aKmftbmOEXyQlvuComeR2cHoUbFR0n40wiVNqRaImz7h31n4okoVAI8QWWBlhdVdNl
vlMKSQ5lklCBLXUx2VDB1fKqV6yewVtdF29ZVNh5q0j7erh0xVnV6JGgm63NVtPTQVguwZ5wszeZ
ND7+LGrVuomvovqV5JGqQ9D59V4BzkTNek54rofUsit51wLzI1smUC2hTZ1eVoa5wVCK6uHFqjAJ
nC1uzcoE6/a71UWnSfneySsXCwKW/w/cd4imbopydduNAVYEm4qR9CDYBIAUAyaJJ0SE7nk9ClgN
m628lcRbqBZuttbF2FNn9/UdzfdAwCkhCLNV8x4p02tRMfEU2KBTD+9kVvTNNzaeDWh+ohtYZCLc
0suJ8SA/ZCwWPS5cCLxoYANAAP37pqOd4+MJbsMZgtGDHzcurrDe3uD5eUulNRrIxTmr59bT+dwJ
kFoBjMS1HrNIGYOW7JAQnkez5bHxlr7vVLduxLRnRN2WY3aNDhpb2CXiX8kLlT0wRJgS4AutkHT/
u/WkqFuG5DCVZq95JePhnEwzVnkf1lz+CYc3Khw7S9ObajjABcrvf7vUYw6wHRW6adRl4Skw1t4M
Tkm3j+rVDglneoT4M5hUSpyJfhEMDunUlI+A4fgj+2irIBHO6dc9CRmHW9iTDqjb/eELGhiF3j5i
IKGWASDGXZV8pUpXT4OoRQXUy8IIuGVZAJEuWrgI3nKxbUZ5a0XeP2/rEiuCDyZTI01G5/YBNLp8
MtUlNuoiE7wut5c/V/rpYydKu3p4cpKmviXEdMsYLBVIvrbi8WK3YfIH09l8UZ6HyhC1U5ZkxBCV
M2po7vSeQnI1UzLD6zi7VPCAopN0znaRSyqrAzXu9cS6bUZ0wX+liOhXKxAJcDTAS5Nd5Wgr1ATc
dOMfOW8YCNog7pAK1UJlxlMymgwbCCFnowDfvpMqUuNvbrjfaDrZmHA4E8Kqqk7blPpY9C5Ojpvc
NxRkZm63DnwATJuDGo3BLcVQRMwl2+Ta+z49H3bT3lxOMsxM6tdZTUkrELRF6bSeCRpYQFxmFm/8
/GnUMG3Rq/dNjF87z7oS9DwoxcVgtDRliuGxaOwGmtWfqOlCJnKvaWiBOJAQ5sZ6JRwpBNmjHeHH
JlUYBX2qUVsv08tdNTuLgUSYT+n/PfDeaQdZIwPIQSeCYocfenBh7zfaCCSK3vIw9VbqlpD3SIaJ
gPkftVPbbZ8N4ZU7ja1/98KsFtVg3y6Z+E2arhhX+xah4kDhtRnpLyRDK0upu3d7y4k3uh3gPFYm
s/MLA6imLWfhT8F585yhJmTdEm6c+lvzJElvVSSgq39V4umjGLyRE3NhByZf/CSnViwPM0i2P8n1
UQlCtiR5nRO3X4qyV32TKmbBUPPknYIFzpbzPTen4dIk9XWMFdsTpmr1f4zPID3kROmx8iyMGYdY
1jxjIlAtmUTnZn07LIPck/th/XFP6S7GB+wk9RlrLq58YpD9bW/OYLyxg8X+iY2yCUNWqtUH4+gX
VZl27IwEIJkL1PNtSjLV5WjGO8cVBioUH0NzwMtGPYm42utvPTb9Oolp0zx0HxzMJtoaXZs2+WtS
ACAwAGX9q9pxpzEUi94ofColQaLIxmNdHbLC9y7X3Ul0Uk2A7aYmtrc8IuiZXeBFLJiF6c6W/nSo
JxyH3lJueskKppdmLcB0d5P4z/gnvlBFly+1Q6W4aQJ0oa/U4pQm16EdFx6TaywuJDOcaVeCmcCA
9Rj2oYEjhzjKrxyRtNoYdALXxX6F1xezPNDsf9YjaFGiOHqOEsZJpP1RQ+5GbBH+A3NFKn+6IKm8
SgIHsy02kvSeQHAO8qdKO8U6GU9ycNkqWrLunLhaPpTCrp2hqPnoINmK/hK6ImUuaaqt30zVckNh
/YCbj/VK1A9wxGULMdQVYcnMZg/On19G4BfQbZ8IV1xW/g5Au/HDQQNTpWjyZg5dnH64Xor61auy
dtQgimvepjUA18qhqbym4uz8JQX/dIfmDru+Q8g04qbPLDHsY3XXSjM4hSbBwGlcoos+j/XuLsrA
DI7Rvdh62sIFVoSLmIFO9oqiYlADhuP0l2aEGOCxfJVeF6Bt6qENOqhy62YOMjJ8jJzsvMZOj6sa
Z60YNAIH8BTK1JjQtG6T/mC6sW+WoVL6AfAkkKis22BQjusWVBvvFGQmDAdmWO0kz/YvZhemjdeW
N24DKezitN/e7K4A4CQjc04j/syvnVHNx/s9fQbTX/AW/D+pAHEjOJ83lXA6+uDgSJnqMYXqDNAi
YNfXqVxbIN259iKveJ5eCRzuPobe/8bw4vhcXQKoi5Am1kiMdgieXUz4xBqVmJ8XjQoLCBG6Oeow
yUKLhgxZi5JvwfSIA6bHfxtA53QSQJW1udSLLp2mmp5bqFAYoCLxKd6VL4YHQy3lqAjo2v1WL+Fw
2bcqw2yw6pebtSAjktoxl4ApJ2XTIX/KknhWg/GZMDM5D8Y3TfHZTXnABOhDzOXpvfoSKu7Z8HCv
EKOL4u7g7it39G9wd18NCnlJ5A6NNRmHQO+1Bc74P0Fuo5cSBYjvwomhjetmoz54R4sonWEx2J63
rXHRmZnsT//xAaqJWg5eVbiEV/ytOGm7cVLzIUNj2IVhnp2yXXR8tRsFz1/t+NhckI/AmvN6usNS
RiWJsqIo426rgjDR0DGFyTEJuJrQmgNT8+40QpfkRLiMIceKQfekPeSJvq4aAaV9yUypIWtyBrfN
DQX3RYOVAsnW8aCLChT2TXIf5bBBfqcZut066CYfiK4H7ZfEmiCTC5ZZBSTPZfoA//cvQ8AK+O2o
4RTvqGh8ESzJH9e9Firq51fpU+yO/G/9gPHCRxIelUyU1cbrCa0RqK0sgALxJ2enX/N8RHhS8WjE
yQgBxlmdWSt+J3t1cCYxP9mMDdWb+nXxGwQ/uyTUr/Tk0BXN6jGgL90yHnnLYQHhvpy2ZClT3ezL
5nB+I1IiOtDVCGze7QATtJXH5ZHn0cifDY2dW+iQj0q/Vl4wOCjDCoesRIx871S0x/EYCamK2sAL
5K5iBnl6d521SAt5dRED1+MgfdHXDfsfkxjQdywvrgff51AUWkiFjzGeThXVyrjrvAG8pM/yGXnG
KZbK0pdosPIXsoOs63jemPNJH7sqIwa7X9Zb3qGk0tKACULFkExr9FjdM2HQbn8QP9h4av9sg8m9
jP+Y8tK15AOvuYl7D9hYNRp8k/fiRxl516CEBsC+bboa7Gv75pxBn5cDU1H+EB4/Q2xLHoNxn0RL
S7Qq3yYvhtpno3ORpGILJqeroBBPbcT4CbSGXdrj/OzmGFVM7VETSd7eungo3K7Lue3bSLFQsSj0
zMgEau+0Vp/2fO+Lay1uVtvImfx1Lnrz9sC7W0ScrVv2H32AWAkYoHmWV1XF/4litrbRYgc9PJAN
Bhe9tS8+HpPkgHUAaFJkpLXmTE0aMchlO7LP9h3TsTKXXiXAFVOXFOQW4F2e3IT+uzG73cwrk4P8
MEtYkk4eQCs8o42K7k/UQ3AytxY2PLZDTxWHyqWK96QRcD9yUs81W2lMAJ0xQ6JaoFH3f4sjBVjI
NB0tX6SZrWkRm2mntgcpe1d+Acr/QYlCOozo8oU8cFKVaVPvBQnOM1l86lg9b0Gs6h8jmGlp94vK
r55fL6LtIjmeJxi8S7L77ctBJm0EsXGdS9bDOFCGGjQ8NiI4EzgVmnbwwbbzCOutR7v4Q0r1zVj3
zIVIo3x0pfjmWkzIK/R0R/MpIKrZnPoREWw0bVBvv7m/705ZCXdXDwF4KkyPeAJl7pv/JcXhHPzl
HpFwp5wsR4FIcDhLM4UGOrEXKqNhK42hN3yJ0P2hkXQ9rUNtkO3BHipvfWy3BB/EunCae9w1o82S
ywcHrWHQfgdWGxoukWW7JN81qLqvR4BU7yAviksWtBzqAZMsnFaHuywWu6a/HnxxOrrZ+nCqeZoU
FYBzFNuoLtp9uxLxhQuUbFPJuDjC3blwE8GGKca8XRG/d0luInvcz2NdpqvyIbla8s0ahTgwA5rb
TUcuUGRNhsJdr9ManHGWjO4CNsfUsJDH1N7gcF6iaSF6OywMjvOmf1MiXkgHm0KJOfASaC1saHGK
ebv0bICPBQtNuAHXEzZ2IGL4X1W/Q8i5x6/0gipD+XpWhm04BjFxxCJPnzWX7/2sWX+ucQ9zXyaS
QjQHQp2xzmw51blWoadZbbm06waj8m+0NqqjIfB3eJ+BV+Pylcbb/kL+ac6QY5vbPnzXsETzQadG
dtI4c6/1BJjn0+XkqevKRpptdIMs+N6WxFnsXSX2gWbfqXwI8nwrPPacjRlQS84ft+kQZRS/P573
QDYmjroRvnaisXwd2Lld79ZhNhBdtVT+3ZF1jjNLCslj1g1d4TAlATt3vBRyzUB3wIUDjcbU26wU
vrUgYkeVxINg7uCpvT1+WlkOH2il66L11pFY1LHEIhSuOhm4pzOi8KetnfGOVnCEPOjaXckLglc7
WyRlnVuQpqk0gmeja/3j6rpfpxoPP3J/ZR+oZEXnRkj2/UUCqEvv7EriWyzZsVnv/tUADmHkrIPP
4Qxh0I23vF+F2r85Bu1UaKdgXkwCvm/dWIN8iKd1d7RNbXDh+HWy5k+5ltIl7l6ifHFsn5AK1rI0
F4stKDxnFnPUbrtGDHMM81xCN36XbPOYHLpLVQJpSeSkPVu9pttgWGqyt+5zbj6EJGFudQglJCnP
j+O9oYk+PfcpuUI3HCUhaGHdZa7ZTXsw2/clR0TEdA9jGqttdV5qHMyDGZY1zNdr7882KIh69x/0
YmwnCMNnxiUcvYL+Hy0IEJhx7sgISvY59mxRdhymNGgm8i8lWo+x9bPmFar8qTiwaCaFTlN3Y4p5
Hmo3aCX7l5sTMij+ldE/GJnUYIHj4xgjZqdmwLACyM0UbEpvpi0AjAbc9Ssmd/UrkfP/eamp6sym
ANYLKfbeBuKVN3iFx3vd5bWN0DFxj1kLj20j4w8Bdr4h21raO+3iKaJGBwmbHP7xEefDaOswP8wc
69gtbLLAJ8ixm0IX+BwyvnG6WrIIQvd6PAoF1yOybi/KxKTSJv7KtdWNlcSWq0Sgr8hWFCc/SQ45
rPJXYAsn8VRF5DkEmW5/Lk7gYb56S+O2R/hasQh2IdbdOZdv0gPEYZ7eLLkEnRArF2/f4FbM0wL7
Dkl2OiTRCgcnrSbT3WtE7EEutHGAsBLFcWvUt+4iKfKL/y7qV64/XUHg3V1I/J4mJmN/sJTwD7k2
otfEIs74Tkui8pzzQ7bWyhStmJ52GIyu04z5EwLGaBhm/g2q2qe+cqKgHSA/dpp6I0ZT4XXoiFBR
FuDRez1lB9YxwIF/Pw+aZf7f0lrSB1f+by8GS3b6Ed5+JAdrajrXTGuYtfj1VaOXKDuu8N4Of0Kf
+dd01NyF4nKHP/f3VDNwgJz67Nec/OuuQfgRr1tmWmS0o9mZMRWRORPK9yhrY1cy9FmTsyUJfv1G
2BW52m+pBTJCtJotUfAu5ESdN1HbQ8DsvBQA7YVNUTd/TpIe0rcv0gpAGh3lT+bbyf16zl/kRMwt
RlyYmyWsKVRuvQwP40yb9YtenICK/0tPeeT4hs0gHBgvE+i45NUvZSzQjc7zaTSqgJTzLQdaWBcg
6F7e0e+E9GVsrXmsX5h0jBfjTrR1vD2NYrkZT+ZJYIzXyILWWp2u6xcC1EG0GQAm1ocLeOI7UI6X
GFN4eOTGd0hZoo1RSEApcHVpiOkJvA2RHAQ5Hhl1c6L8/f1VeDaEDM2pt3vEcVjr0Zt7xlAmTXxf
ZEQK6rhAA7lRz5nSDG5WRWKCbinfGIQMYbARp3bEe8fxoHQ+Qp8NuHg60EE8by2SEkXjwtjg4zvS
n39K+hE54bYfm3CSAaBX6E6srAK4k+YhuO3+rQnTBSgLFDAQywOg+LDTKltw56fXOebHyX7azJm2
GYwkhICM7WGQsKI3jPK7aMxMeKyKGJVyx9qa9PeaOf0TNHTL/A/sd8I3uX+6gx/ugVdhf3W1vdpO
kbjhEOngHn2SQWCcdVVoJJuWsROXxLkrPyvTAy7Wh1nJRUwhtnkdzVuFQK4R/F8HhbSi0b5eNJaS
5B41F6GgsoMN4rpEe39/Ykpv6iguzfTqcIiv2RWbms8NSRghvo/5ych+lPFvzirIvhatW0wle+fX
tj2mKyxyguQVjVy9TZJx9T/JAWJ8
`protect end_protected
