`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
locy8FvHPdFgeTlTZto0ajtMqY/IhpJRAqnLXddjrU9orRkY0mMrTCj+5VMYgCflwrLfpVo40J0d
YrQU2Do95w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LYwUmKRVftfwarZtnLVKz4JXU+aoM26hKalkln4ZJOXVDq5xJZYLc7rqXJhOXoZ0/DgedyQTluOC
++LZEiR7qct1FckHSXan7EN0LIuDR1+6kR+C6pY2rQX5bqu4xK7lVYNEQTWQNBahWw7Fl4DMV30T
V0y6FdiocP8A+rM3hO0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aZcdwJP2yawcc2jVoDxG1yc7LVg6XfQWoKkhD7E9DfYCqaCQrsDrLJdA9Efcgtk7sg2XfWc9bDO2
Zk2PiFC763XOleqA+/a261WbEuh9wP7GL/0R4qjzndrPcdXy4bjaGFFuUUhEOj7OpEnhHHC9EAmn
tjh067q4kgJ9BXn80w06Xt8tmkQpiL4+lofB45rkjLcxq8zCi63Ifaw/5Y92gHtjEAKDYLnShUU0
uNRjnSt96RrwFv6i6Ry5zOeqov6CJapqQElgU9YywiAl/9jDEEVnjUkeEQqpK87UlmDdehjtPcmb
gXKg1Xf6SwslmN4HdWMi//d8rhdXhsUFrslTtg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VrOWgfhisrPEjDlVKUVi8ab3R58u/OdlSbdok0XbNsMAx4d3CKPZH09c5N7On8k/U30aDljZmeOT
ntXVgk68PVRioLY7rVDUBSIevkGy9Mwo8NHOUfPuAN9e8jVN+DiIWbMJD8GeEiB4hQC4FT3K28o1
efzjIBVspG2NybyNmKg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PtXO0Xo1Ly+41w2w1ppYJHHxnNdyst0QMrPz0vTThWJET3MP//SLLwuf3LLEhEKCWYuZYykUjAwJ
RY1foRqktcPnB/QA6jW3+yIZUttPClsqZwQ7bEiYucB51Gcfz69hKwwvYkMED41aAjMc6wxfHuwJ
RFd5CfBPMFedROoj0fBBM1w5SKgtDoD22BdJbi9DdKM4yMrTyRiM/NlsS8jZs4ko6xNtYtaAX9X8
qXuFnii8QczK1MxA09/BMEDlTJ67LH4VjS/WFcUP3ZSrklDxvZf5iZFzLapkO6uW9Y3aIbu3Wl1p
Cl3viNrE0PyqJbogMkAy4l594yXOw3FkOlK2Dw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5248)
`protect data_block
tWcP3kLgyxQA/ubWSdCO70iwtqrJBLAKQb6ZJtveBAKXh8uX35lNf28O5nMCoNzNRfVDJ7eQRMtC
8PPE1PbPYZ0nKsaLAF6HfREMC6hfIE11uNu6el1EDAFMamxrOuZvD7YoL8v9ngKRV4F7MlREuBFi
o6EC8G9dinqK0rvs7fxThoSuEN99wgucF1PJ4oM9oIdNvjd7OhQwAgQFtpr60sH2mb28LhtxgIlu
Wql3NXEq7TFZ8l44e2OduxicaSqm+530A3AvbDuehadzPhFWv1TxvnEKIk7DG80YMfnef1HtWJhQ
7IZVMMnBWuiVUG3p6EBMcD18mbh91Ahz7MjK+4+I6PgpRLr7/lNNSbMvQUxbsvGLX1/gVnXvwlbn
L+JscfBBnclPCA75x6dx5pmd1/amIAp8SGbWIqukmHZcMj5CEPF9h6wFq2As5y25eFhkDJGjmGVP
jrYz7SI/b2GhDeSCcVAp0YTQcMDXnF0PjcxxNGxaHj6P0sFCMG5jgie3uJ95Id5meLAYTBtwBbPS
RYwNU93VojatlDyefksZsAhDBeDq17UFV3L0MaYLcdq+4nT8PvKLkaEQ8HlbVtUjqjVFvx8vcV4Z
YAGPU/wVxNSRL6PzH2i+TAMpSHjJ7CSFZQCzRzyCzLVtVyQZpta1065lxvwke7Yu5ETyHTg6FJ14
YcRpdugnsix9jL12odiryu5OeAYWi9NY3haN8FKBLWFpc4FKG0OnqwLF31pNOIvVI7YatKfjhn/3
+2WXlo45v2M6f6erddm1f2oI9uLevQ+WxujaU8ShXZ5SgJz1sxRqADE4MajT1XE5X5F2ShpEGMH2
j50ldEOMmy6jIxF3Z6uLeLzkMxZVYyx6TEbfSq8qFKIzAk4mKiPcZXhqguyQnBleHIUGiJ+Jb0Vd
jdA9bQ5bnIyWrjgT9nG8+YlTIWlmyLN72yQqF+Z98aSbMKg9CDeTYZCPP3RvpvQGtpt3qovUK140
brNlolAY1KAK6Oget3JpndotgEfHMx99Qth6Ocmu/CdaDA+kY/3bQF27p/BYMZ3FK9eh9OHjz2xz
cyuXHmRrMQoK/VQ/PO5iugRz/PW5HkMXhHFptu56wEnlEZJU+5P5dfSc3QTW3Z7GD38UENRZT66g
3DGW3GmYdJnfd0OIKGZs+uZ59HQ+mlO7yFUddtrzrVP5pXCinciLxQLm7ndrvRboOA7Hb+N+qc+F
Iumb829vpZ15Ex3UHXgKW6f3D2oMfftPXzmg5IpejmjUxfQWyXW18T50MzCYQWDhRYEXb9AatSP7
20Jje9EwpFceZTGP/3Rbbg9LzxEebxhFysmrU8V9v/buXk3+WYm17iQ5OTlzt34ssa+me5tiLpve
gJbE2TPvndDFKr+HkB17mn3b69I72iMKnJneQofZXfxVcqvlCN0U9L+mCLIiY+pa6WBBxjxFuaHt
rrtqryZtkZZt4GTFdBk4Z8u7h2Bp4h9XDbIgSMB/VoxFJ4maQp1U2vQNqauO0TqXZAeGn+GGvT53
t26r4jlMfdRtsJYu9Oyzwj8EMKY0jaf4+8QHrcJBj27OcSumm1hWrjjB91goHGuU36X/fFt88uME
/g4jfiWNqIKb9I0DBVt3udALCgqDY45H9JrTt0RMySIGRyRihTO0RLzh96oVDgUBXLJM6GzUP4vJ
mWOn7wx000iy4t+GcvDp4edk93mehufXU4sM8DreI5zPEFOiTKPpp54ogJba8wqD/Oa9sXyLOsvx
GDIRnTJjVU6TzDJfvH+TZUAwcrjTR0HtXr02LaHHTmTsZcrsCBGcvAy9y+4OnejOFDxQO1Fqe/s0
klGai32EwmM3P6ZdqpUZHo+Np9KPEMU006GEP7YSKJHFu0CXykgo6xZTLFkNURb5l2J0+nBH8x21
H0DM0hHowzWzb5AmAz1ZCU+Ulo7ak4T42ERE3Z64KOGHo2rzgIB4iugNQHOa4cix6bbIsxu0jOHa
kAbvLDIj+zYO370NbrTcT4+NdqorGETiGQzHBUHCnH6ZxNM4uHpy341A1OsvXbHKvaaZo66RlkRq
Ao3KQ9L9G+slc9oGNx8Bg2RMPN/9lj+9llKaD3OE4yZ/HwArzoITndCsn3FjNanGyjHIxd6rFgUh
j5WrFR7lnfGHWzW18J99lG4jtM4Invb3cKIU+ysUfXIIk/yX68Yo8rvTmvwUO0NjyhqlTvMl7v2l
Qw84OF7WeR16OEC3slML8ERTRX1K1ekOa693a9izZML1mpT/H9gVOs2p+20SIem//z+1//lL52RZ
pokSk/5BgzVg45Y00Cr5BvdSU76i4S1GrRcq7cYw1Tgs/G62lST18aROZBpW93UgU731AovIoT3p
zyd5cUgAD5Sv1eySTxxj/cgLlUBZxWAIirApjc7ZCjOgba0AecSHq3UCF0lrbPNF62k4ch/qV4LN
Cb0lXLguWBrYxqs+bc6xSOdAtp/AMfu7gXVLhtD11erfwNb8Yu15Rh4zy8b4ecZUp8zq+c7yTlHd
4lsoSjyKgZg01YeNOiz0uFPs2kr689TihFGeK3afiGXMI4dPdu9NWVKcHSjHct9S9z4Ha/CIn5iL
RkwyRWat02541YOakZFEchDiaDtlwEv3iq3kNsBU39l/tr4Kak0VGf8DpArEjnbtZyvqS/f8oSx/
uwV56UYsrY35mJ2ogQ56e/WMxIngTwPCBWxYU5GGyh2jwSETD+r1xLrO3sqbhV+zGpJp9oiETySq
ksjd736v1JrRa0Fw2FIVQsi8C0f3jQbavcn6+PBTyvB7tBdSYdBckRF70z5UkjLwbOWdVWPNlrer
qGP90CFDsxfqf3r9vI5piqQpqgDdUDx2Q+eJdNaxZijamoOcAiKJheLkqGmknxWCMK7u5czbpWIR
IdIEZvHTUqV2Y0OMsPqv+VvKjxFB6QSwWlWSDhGCc89CZM1sWqfP+XD+ZO3A/ox7R+DhQ7fP+MP8
7FkbF034xjTu/tnDEslufNgsnUdb+Qzboh8/UdoPPa0/lw2ESOg/DO1aU7P4zwJpn91mIUjT/kCn
PGXXSwDuprPdeaNpSaQKIU57bdnCFHDy269mJbgRfiS3kPDs8leY/bah9uuw1VWyy1BqUzaYTfce
3HwmgI8gIbb1qrPKl6dpNiFK6gVayqIr+WADjqlYpNheZkpSifneJxc+Swi6Ck+C5ozOl8+y4n/E
hBsNx29zjAMUFXSuMf3ddtP6UxEGr1u/fxtKHyzkbxDilSC623JOkcddka+ycJgAT/74trjQ5nb6
Uf2UDstO3pSf140fSy9feHnR1tJ2THWv5HOOjagVpCgO3oNS8MNQ7iPuI1XSd+yOTQ9NYCHD9lKK
WMcEpotPpX/DJ9VY7LZucepsrhULsrkH6a0NOmUc5Hx49DTuaoTACLkl9omoWW0k23qvpQaB/Av+
ThsyzS2RgWiHQEycDSrAqao7Rf+DdDE2oj+blIeLtkSKjRI20yVYk/igS2wA88TESQFyNDeOJMh8
+ig8NYBX7l4uU4sa2CevushQQ3zjNt8oRsYjd2BVXdjM/L7hPZxpb7clBimgfGSYYr4mMXNlCoj8
CrLyPSTpAA2yCgXQfkGSZCZsFy/nDpWV8IOli07dZlNaAbXvUJWL3EpAxmEQKnB9Mtj5sVYddRYr
+X5T+msIMP5MXnFlp26eCV2UaIyFailVkp72kVdXpXGCSlifOlvewjaPFO/6Ev3AhS+StsKhtz8Q
jwKma/C/1GGFOPRo/92g44fqcONqUEIFpyAuRgliSJ+fYm/KU3V7MNg1ymBg/jXYk2wl7j1eRNYI
t5f7/38U7Br5AjiMIVUs85w+Za5Wlo/g9+fSwzSmfyjDMv45njK5gkA61bSWVAFD6SWXN+d/2kqn
7ICtDIi6PmIrN7wM+2dUyU1JmH0j1JtSsVaVFYks65nJozRQtKwpAS9CsNlwJx0JFiiaLEuKGYKr
I7PHUI9U0fgS4M0oMWo9KBbXBhf0D5vPBpQzwduWFfBPB/5fUJMY1LZsWeJ0Lv0uZ+PLxVU3M3ri
wMk4x89T2fMKAU23eVLabGNYybCdjIeQrZF9a4SvGBTD6I3X3IuZMBGrRlQ4E+Ct5tzVl0/McMCm
qonkE3CbyT5qz03j0ZlgmKY0icJwjpveT8btujKIXFmX0y+1Tg7dVBMb8DnD3m7lDpolXWYCgkIe
biiAVY2xlkdub8Xc5SqA4ufgKX5ZINBG63a3xoan7fWhUBJjkuuBs+wA2crDtdvokBv0JGAvcOAM
13GI6kxzpjguqMwzBnpYFvIZ7frO6F/HlmBd3lcxWzZ84c7Tatlj0X0TffG3gxldS9MSKnAwZJ/L
gnY0ZOy7oTQDjzyzF/LK9pBBOrhGYUbJCkdyNygBTHeu0P9Hproc11EnklIfp/W5BSfATJlquzVl
rBJwJjNj58Q+NDFs2aj3Fe7kycGawAYTx4MuYLQTf2yileAWagjWp02NOfz6lwfx99JYhLAUPKg4
YgyOJ7hWh32WKSbXFBu8XEYhRIPikqo/jAQKQ1IeSo7xWfMmKUfjDpe+3Mx1ZMhFPTIf18H/N2BX
dAXpxXeaYGyRMIJT8Jtu/K9+pmsnaxnTJE36xpujIXza1QSrNmo/bE8O1OmPDFjDPtiDi02+cgUi
Q2WW28syGUjRwLxki2js8fksOEGICtg3vMrGa78wNQFGN7iX2HW7THQ0gzBP0Q4fqjHcYDGnHf2a
yRkY80p+rO83+NX8+NgFdSxI0uoGNwleCN85cANgy5DLk4pCixfesU5ov37qzLG/ZicFAthYZpqu
A0Zp9kmGX2EhrQH5J9IgWPcwFmlPkPSfIBoZTrFIDBxXf6t/tqIoi03b33L3cPh0OHd3tWWd9tdi
SBK91tHm5CrQWm3DCY5a16Dnno8NGo9uSmt0TqkjvDPDjXg9B5jmBByPZYNaoPMokC9bRmBO57xS
tupsL90YlRMh7jH1DEPZpl3KrPNk6gihMzrj6Jvt0OUyoKlNcd4i+T3jAxmLxrVx/gwjZO7Q2ViZ
svGYeSpa/dKiXdA33KdhfIRBX7vvAqK7ujKRe4HKiH22MrURkEKR5xNg7W0q0wFrkicjWYBZIxvQ
UFyvzjOc5V6ccnEIW8wsgs6MiMBAmcXexWqvTF3eGRtoYd9NB7KtZz6cDKfh/xTLep/xnIZEEGi4
HkIe7AxAWrZeNX8h2ejhcri9cEPQNbp6/2xTRA3GWQGlzwQU06sh28xfIX5I8LfVw+cioh7hK+V9
cPKBcAozU85FqiD32Zv5PxwRhfo/0FpxbEYQF9bFBGdBjIGxr0YfYim5QAVMTqWutnF3mJX9VrYL
ZjVUanqtKYDO2z7UGF8m2ycq5uR9v0FHUEzgUgK55SKvK9VwRdUsba5bwmtX4btQcZI8SngPCxOq
/epAwvotnFWgylS/1QjNIc5JL31cQaJTbPkD/1Unl58TAV/2yUWGidu0p2IUow6i54imxM0jITfN
vG+dViSMSN8MI/AEEV9ClwC5fMSXTqK2+fWx2CNQCHeSrw1gF3IAXc1Z475SkhcHQHoacAAgabBt
XJKmT+dmUWCepm/pZC9OQpqv7MC+nZTejYraQujUP59EGppDpzdTEMXT9jpI2ICGpkfuRwkA6wMk
0IpwKXG7FxM/x/K/hDqBAqQBsmttidsaWmBFwHs3Mj36CVyMWYdCHO2ggvfuq/FJzKgw2eRqLE9j
JnAX3nXgsGoshZKS1Zq3YTvzfNt5kWtwpsa5uzIwAq/Racm/GE68kTiRbsGG70OPgowEsviRDvWI
jN4T4GSjw+Vel4sGIT+DpM6holfA9Y4s9QwMMlqKGR6UHWE8kUeqlSznQpCnBPrt7Ld3SgHHwz07
NuCMeOL1J1d9DZ3yLDUakHnsF6k4tnPWh4jegT/plcGKSFNx36Y/jK6MEOJL5sX8Uwb1mC/rOCU4
4zTXHL/nUd5FFvxbakCbH6Om2zw82WT4AI4zK8TJ46JOxye7ZWc0dLImfDCoLGv7Vdz7mNq20uMG
sfNBcitaAuOTK8ZU0hwTXmup152m9tRdMqH8dHcMWwdfEVJhX8UuLWpV4vdzfMdWKWWbA7Ci01eH
jCjPpXspY4vaXJ41NHCgB0OOl3hLLYMiiLTkQ3YfMqUazyE7R7TShvZEhu0JQzihrYqh9113eCFf
XQ9QuyHLPDvhgbVqMJ2bVcoeRGsE3r6ttC+llNONbnPCQ7qB1YnHLELvr0l7gFExdcYr0yx9rKYc
fGp5P3pwULGl3RIFCXlUIAk4XCmG7qocG3UxCrkrY3xVuD7zKmIWy94x4Q06rDnShZTnTgREpNqz
/PlLhzT5QiaRImPRhzfzCoYDwuOARxDW3vhK0gHL9VrjpRt86gSZi4B+0xZ605We0osT8k85jPJJ
0V3P+DAYY/BS5XOy9+NKVVE/CTPPUg3xV2gRajza5Q/aYDlQ1/45/o4fx8M540//z/mFMIm1OdPH
6x7IwWFkfqavF3alIbiBmhnvf8lEouG6DqD+QLOGaSIUwcC/dzYzmfeoRZMEGy/+C0x+U3okUzCL
5K8vxZdTaYSFJOGbZgStuPkmDoDqkjOLAQMKFi3Uzqun1BGtj7cbq/s7Hks7+pp9J283L+j5wezI
CbDIP05ZfTZPvP0bBE+5006nRsUt1UlqgJMISBzLv6Tn+j60s7MVVINGFq1jS6v/WwKXBiGrvvyR
ENX5jiAsA9GmXp26pWhaiKK/lrV8NAAGcRPYuobwqcDViB3ZnxIoEtL4VX4evvpUQ59zThr8KTab
zJQhqRQ4MHy3nWftUxcr1Ne6JT9Jod8++ZgBztV4MGcDBPSfoek+253tOCbztQCRYjvMsakng9kS
/JFFryzz7Bb2nltaxLGDMGD4r3kQFujrQVWgkGmM15wpRDk1/fap0Xf34BP//dS7jHNJvH7fzTVj
rf1sWlJLPNRmJ+6gDQNi6nhO5n9aciZf5Lng6yxig41bs3RS+OhWZlJJcLW/2UT38t/uAFrmnQJT
6CzavQ==
`protect end_protected
