`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hnCZRK4wsQU13zrB4/5979i29XwKjk4+VHkzEeFvbw15zGcKElzyXw+3u2raG+jyKcNgY5KBH+or
XjZ/iGmEvw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aNt5ib2JEm7gyFIUh1Y4cTmp5HDTcwIWjAHWiaHJHP9TcNRi+kKt1izQC4t8scMo0Mp5fOWZiNC4
cX6NOkng01UrNOdpe5/GwZiqVLTxi+H0VJaU/C7KePqKQwSNooBV8Ja6NBT1LL6s+8pbfOLOrjwe
pTnt3ae3PNIPKNB1UWo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rzb5SKDhpsUv0MuN0RqCsxMkmf13fh+myD3zY2SKweuxjEmZ9pznEayRV5Tx0d2Z6qknNaOKPdNw
z7rHlnEgONkmuTHsdEwMJLfFGPz1/xT+KcFh9RI3zpXffboW/+aKCL2kK7bs4rcOSaGNBwE9Xt2E
bSFMEurlQlprASI8b5Tjwxq25660SoYKxCaqYVtqnTKcq+Q4XHBwA6om2TAwrKLTFveJYhQ8BgY7
H3hmu4Ac/uquDNiYLCaxdwpiSDS1mbCeFfDDoM/Sd+vbtgV0gf2+IhMf1CpzT4O7L0nFwy07OWW6
aJbvcUc3H5RVI5yR1BqOn0yckd9kvm80xcSfBA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X+vFLoATdf4whEoYzBDdCcXlO4vGCCVpulqqGuDahhQkI5jGJQkDp6ET4jz6Uq7lf+YPtZdhfod8
l+3Xb3iX8kK41r7Ydp+rrLy3kpJnB0mealgovPOFTxp8qtxKYOl+6UKkbOKnxOeB2j2CiZ31PNKy
cUkAQnKBYApHkgIPHr8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aJudplVCt9yrmhQwJxIv4K9Hq1/pfFtpbtJH019MEY/SCQQcO54BSvJ2XE2t0AR/Je5FjFT3iLp0
DQbFor96Rnxu52HJq61z+9kHRuDud1w+KHqNwwmb1wFKFWwVnt5FEawQFarnM5gPB1MlzGjGwkao
96LDo+JgMKwmeVHwy/ZfBbE3ING/eetSLy4KZtId/4zTbKeYVdf0L4x/rxZ8MAkc+SrVnYcH7s02
B4oufzVPXRKu5RIvnpNPM5aK7dHBJXG7ONW/V99EPB+SWFD7IJA97ceQJBQCYGDYCMQGx8wmlcEK
GdU8ZfufEEjW3Fo0KmAGVJ4O70x8AfSXgVJXZA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25088)
`protect data_block
/AaIlSjrqmiBQMqYGhEUy7BOLPub9DG7S+DxMeylu14OX/1D+6Ad31a3G2i7PxRHeFK9SQbKa+uD
Gz6lWkKJ0y+RDR8ElzkLZdO/cF2Xy/3hlQuW7ZVee22EazgZ+UCAUdovVQ5Kb7HcFSKoBGgzFuK8
cAX0up/7eIZs2D5UeEFioNze9UdZGw5Hure7gKSJDr1B6eW8tSU6n3FgcreCJpMk9ss+4KJ2WUGT
PnZwkuNdtEOsNt5td7pnprWAbK6LDEPEivNQp3/mVFAVg1wFrrnQNzU3w78SL5Y/D6uGXBKjEvtA
xjLt7XJ57VrN5yWvORW2XXK0bkKVJ6shmoMIJV9CkOhU2Y158kRNVCezl6dvv130wPraNnazkzU1
zux4fpBE4Ro+3T84MbUFVsJrUZuy9hj6vRd+XABOOdK/XavWWGaMJdnUGhrc5ENp51oPeUdGmtw8
t3blOtB+emhoBrOsz5FQjmOWChdoXKLliSchQ27mQl9lARk4z0sU7MHTuRfMSHujUbHQM0qTbBwR
qJYoc0dT/3QIp18iHsFWVb7NOvwdApfYZLHr2rlql5Llu+DGD10SUAGUSmr8lPdhegOAY/9GkjTe
iY2C+Nb0nTHWeaNqOWeJ5xIsjq64Nee54VllY8yaXUEkFySeqPRCy8xo6Hg7uQjpAVpeS0//nJA6
GgDa6W84+suctX+GO2vGs+I6SK/aYij5Ybt0xuyEOUbyKa4I2Rff6iUCXf+E5UGApE7o2PG0QePH
/lPRzZIEkvzOU7CRH9xcH6qvBCLU+FIJaZZbTVrGQMSN1qycAkNJojmX9tj/IrzodWVuTaCyz3m0
dzRpBFPtLCTVvYgaOQoygfmdocrwDB0/jVhMvlpK+hAU2EiOYUkGWAIgYyPDr/kcXg8wc8YU9xl2
SMMYxaCWXfi1uPg+rkX7ApMVbE4wznOt7+FY7BWTIAjspgVrad5xslFpnnQrye3YlE6cMEfd9uFp
Z2rHvtW92pJPX0ShkPDm5YiXRwh0mWQGYUc+6pFJTi+Q94Yq6wnXEEt1RI0q74eTxmY1X+YhWxG5
y8wghZiETvoRcp62zVxTV5U/4sZlmmFe28m2QKARmurV/fkJmMxX0q+2Pzgrfh2whTjaZce+LCoQ
DkSsmWBo1e/UlLtYa/Kf0DE5gnV0ckyDSVyzZ1uH0SFiI5Z2J8K0p9lfT2Fao7867Xwo4Un7F3l0
oe0UibLQAE6IwsqSf5cGhRrSFL7TNnL4jTZeXWptA4eeQI0u3R2GMwtYVvvNk7pAsci4YeChg7ZQ
gP5Erihdl++nPL9kicrSBjJf+VClTzdPf8WG7mnIwclnQYujCKSUF+NDL24SOJrci+Z9GKlJbzFh
C0DBJRCWgrpxu3kiTBZw6ZJEmxCFKTB2jehaxkASU+vW6KVhYYrHpl1zvp4Amflqeh+sdCqO855x
4nShSNuWM6xBjQ/hVMfEtYQ3G7GjObWVvPfK9OgBFgwCm+Oqixz6UT7JHn8TcXeQNW3kTpodixdQ
8JsWoSW1pi7cczsr+4n78VVBr/Sky3lTbhf/GCTpGOQ9M4hCO4NxlVRgpa5MRdJ0zoQlnC1R+uRm
wMF7QqUL9tHQUA2Pi9y5suOg0QJ3nPoETkWEkwohZaglVw1ky/hhramlD46fEO77+gVWA0CFniYn
dTwgrunEScI5zKGgeWNEGGU4P9KDT7p2FglG/LP/XicEl0FLS46gfNyhqObyIlNSn3JEpMWKvoka
cCdQ7GPLQwQv8AnTzUcXRuFva6fNZgmWBwR+r0PcNbvsM+9HPcCJFNkg2Hi7CBZp+WwyomQJvT2O
+PhzhdOQi7TusAtqztrasoizt5lbrhHZi9PAKdaWTFA9kUicB39izqNNGqMR7mz8cwQCEyTxCKww
baULbXuyytztLhA8AAZ6m9RyMFmDtW+wHb0QsfS4tRzTHd7J61YvXlFfRAP9BmryAZWXyitAhREV
XDcFSUwBbJjFDl9K3mXVVZp2g4HyF7SmIsNfqzgQtTuSTiyN4waSZ8YjE4cabMwhF10U3vN9PFcx
PMMhudG5qUMXLyhbZR7+6JwMRiRYVDr1dOoSy6qBzKYrwPhSZB+5JA1VrWdReo3gGJJK43TUwGra
v0k3KhwTDwihNMZEu3//uWcgblrsZ+DNrCIMsYm859QCRw8bQoRDfrkNejz4a8q7J/4pVs3S9vL5
3HYNCx9mi5ADM92fgnI5LWsN1Du0gBZDqKXeWpmotpnVYHZyYDvd7sdGhOZDXOR5ySKWPtIgfr/l
0WGw9jO35wehkljd/wyzNZ7iZrHRJIxzlXsKXyGQezqm22CDrw8tx8J3pa+55AXsyit5DfGB09GI
f/nP5LsyuP82wDBEdc065a8vk0PSftgZZAcLWzUwkht0xqyO3VfzfezaFKk8qiey8YQ4VCxtPbNw
UBr6icn/rVMC6xdgkjOPjQoJqM1yb0dOuM+78jiQtwN32FmPtQJWM2Q6OJKaYSzr5qEJHxJ9SqUX
D6ooQ0FPTnnyPG5OZSsOI0e1XSgW6ML5GtuACUTiYfbNRzHfEBxhNnKtJaccLv5JP2CcQwNfm/pl
teBoK7BbL1QkHgouHE6OYF9hdNXjQ7IKWvMwQm8Z7J8ZaAXlXZWsz/cd5VpuB7W5xqZxNKPP+NDE
Rw5bAMsGNaUmA4B1+1qFh62IwfE/4qNJBOCupabhPI1nRREf1pcII7soMbvFrTEr5KXUQ5BDOUMe
ac1oa761PoPuqqLq/3g4XAoHcKjwM2uzvFE1epQjXdOe7MoqWigILVKdS5Lvc1m4DGuwX4OBls2l
xJXehwd81d7SW0GOtSR80lxs824aCDUyrYtUIvD8B+LnPrPAkMpufcDyDj3Svh3c4FrKAy2LngWA
CMbebd3WDUVLdMyg0M4zzRFsK2OxdmuI8dsvbHHlVDWA1+WZ3gHyYCCpWKLw+o6tNwQ1EhXSErht
KVhiSD7kVHgKQ1KaV7iA5oVq/YsW9byXA6p2MyJ2RJs6fqVd9bsW51I66P3VqFbarkXNO0VTreOe
Lbv6Twfe/fVkAnEO8OzorEJuShrA31bxYf0K37h8Ik3QIfgzTSuo0kjK/dFKED812haqIUrX1z+5
hTAhdLBwuvsIClq44d66cskHB+U+Kh0A8b6lWs9IfNFchz4KIQ6qbJp8kyByxhxcmiE0yy06oKHt
KbKrOCRpa8EmptDgwZijgXllc6ZA7xtz352Go1FjzwE/DTzSbadUmfg+c2tQ4cc3wkDRIxkDVoPW
oDZNv720gW893CjtxMUgB/RNB+rdMlh061q83q7GQaPlpDC47cj3mJ6eABILKwzkdCOVlobbVhzz
uObBvIXiepukbI84Zjy8n0pdVx0I91GIwLf5igGGqHQQta1bpSLu9URQcl2GQbPHeI9vWrUtS6g9
+VP8l938GLzlF7XcTh30NPm/4jWL5h5qAu8WPfJ/TNnvrzGPGFjDOx8/gQfABuxeGwazvO6LUvv9
ywoAaemD6zJzNyXjbDRewh2lWucteknaLPW9uA8M9rVODt15SutWqe8p90oz7UDvcBaxClrjOj1d
zHFK16eJ50aIceAVS0ucbBfDoOi53Tl+VxPeVZVcCO+iYhcB4JRvD+oiM2SbWiTgKXTIHJlw81qg
HYNc5B9BGIMwpzcmnpmS3ELpntgdMPEY4xPgiLx18TnEElJZkmbzak3w6nvNC+C6XTNq5FXzIc4L
54+oRXppWCAIfsJ0ydoXwbus9tO+yKvYWSL2tzj7fJgv0PklVxKQNW19XTSexqaHJb3iMMp7V2N6
mFRNaMfwy7qoJiWjtn3AeA6VeMepG1gD4lmcuinO/CoEFEyefxdEPSRManuiWfY+02w77CaUAFeX
q9vHwnevQPlqTio6dhAsL93pfj2iLmkHzZvagjTUajytT6ebeYBfde9QDiwZz4zOSu8pSh4/Qvnx
VMIS72gdBB0g4NnIyTcWUNip9SD9uh5MMrebjah4lIQ1NBcA5W8651nD++vaxZtIYUUImdfdbIhz
ugJxwAEf0bLyIese1AGn+zy5OxzeMAbk3xGPB0PP0/oPbkR8v5nxZhQu3cndvkX9nOUWKhqwVM99
Y6mc3VV6Kjw78woSWVStRA0JILvQPaGnnaXpHaaYfUzSNwoGG1dw6L19ZGh8hQ7tbKvsluB2tsck
tNozmqp0hZueofPe+DLPOGdh9OC4HVs1e1Yi+cDfOPpir/pbZY74wCaPFBuxMVFH3Z3zSU6dYd77
MRxQwJRzXeRaCcF27yvIu1n7FRhxDSu0oyFYXy/c/vclbJqRVRRUJh0Djy32/KD9CNT/8D7yymfO
VWcmf8u4/omQ89qIJydAdqb9ZQ2aOhUjH91Ul/SJpACVP+7XTEZCJL8pBCfESansNv+BUe5wnjzS
/9jvMo/+D4IVc6W2IXdPgyxU9tpjibaJ85CIBpH5nBADj4DncbmG5eEzdI4IihyUzrs6g7P4VdmS
o2W7/uzytrSap3HR1iaS5uis+nd2NR8eiCGhYKCnuzdXKLft/czf9drZx/jHY6xs/thmMtB3ylFW
X8KMGpAvyPnCJocPHzlLvkcoGEacvfYa01xY7p3WHRPJBCIt/sZ0cIOPXsfG0tvKRtBSMAgjWT5q
euyDFLGGGIhJ0YQEy55G0dVMl8j/YMzJsPi//YMkzxqZEnIvJklTo4jjgXcOfnc6EFMDrGsgy9JU
0f9ZvS6UudoyEUvqG62Vi4voHqZKp+vUEr+R85hmgrVDdRTf8k4+C8Qli7N8GHL6Cfzh1UCIpARy
x4rpcr1GQxdgDKAUxdBNcb/2GOhMn0O4o+EoXZarmO0c9NtnzkCS88ckmRkoffel+aOc3jTQeACZ
9VJKz2DkrOI6DA8ykshUKG3+/98EdevO/aaYYAT4TWUCemYcnd+RNWYqGL8XREhWlh74GpvRcc1w
3EKVnPU+brvElouQn4IcXhlx9w/85y41AbNvS2jXzFaOaHuaZk/Dk9pcag6tc+egroGN0cuMdAY6
Vxn7Pi0jy7XzNjFThwwum/QPcQPq74b/EPt+0+EhjjIS7jq+WxNDhGADqeJVeWzznGz5VwUkFtx8
BSG1NWYWWUlcqVPfZ6ruYO2lk2o9KlwYRimn2/eY8xVeMgIOwWwW2gEOWMtMJg8Pf0yzVEokU25H
ttG3Q54VN6zG1UvSMIM6qSZ48buLbaYkD9qjP+muX83FSjYYEDnSLaCawbZ62Do+XXjH45BdA3Tr
+rsunQb9URCyMFyravjKIfueepPw+SdSUeUG5vCX7UF/6IdZEhFiqKabDElppXrLlhIboy4hNLCu
GQd4AL9s22wXtxHnCVVrJwP9qQyjd5QCa0hjO35l7wvKBOcIYBuiLQ5FmSzvNrOMOk8eQx7ys/aT
6d0+F8RlIGeJFywjviMwD2bDj0cIo+1grAW5CfVCwBiYG937k6M0AvptV8+Q+NXTHnKsnvJGKS6P
ZnPfwT9I718GNmQCN1aDv/8Db0lK9+gcdxPIpShoVIL6ukeLSuHeiY3AQacPzzFG838yXgOggxSO
Jn5l26LU16LpI6FbSSLAjyjaZKvsbm2iJqKU6W8BSRvwhudPE1pNFFZJCRLu3oCqFMUc4sOxzi5x
v4tqnoWt8V7q3XH3D+2HtZqlZWyhyu101hnfVxLrOrLOe393uTqYSkQnXp4LUsiw2Jmu+lkr4cn1
3z4BjlPbDUc7ZAhDfQLUyJyxAIEBenzROJNCBDMIKiEwvKbWoCFM4C1OWwbuXQi/tGV76MlLgtVL
o/+jQxta7mXLGkO77GvPEPKPj4CaBZlTWVGK7DnxxwqcWDW9c9rP929wW79QyIirYwBfSDW2ubAp
gSFTRHhv9OO4LuqAN1CQgqN05cHoPSVwijpc1lCtmMX8xEMSd104KudO5+urEsI/oDBITJqTKVDk
vOYdC+x0no+z9IMVqyAwdGxrvtvue0f7Y6pDFXKRzfucwzXSzIwJukcv68dtP8FZ/3HNEml4zaSO
lGTinJma/nUov/jiZaMetEjNDIss8TDKfVv6ZmOYJ1KkIkNBsDd1ZQ6fRdlsbokgFllxUHz3FgiJ
rL5jSgMAJtA/bCYwuQmmaHsZM7LPi45M1/zv1YiM2V+ZSMIyE+OgJbli+7KzsHHoZGpYL/sI5UN0
fkviegG/YXBqIclF8/v/W/XdFQGNg6QWIbWPX/sdPky7T4/KzL6z/tJxKhbQSNJC560dvW/miOoq
GUjFM0Ix9gXBjJn4CnTUa+r/0FodDHO4+mIEtHKsl7qA0ZNBQuuHqixpt/+a9mlOSUvsc2CVw0uD
ai9fDo+rxPdHQwdaXNaBFgJlUFJMPHlJgVmsUjpau/SKqIfQGXmAT5MCkaBBwCR1SUylW+HeJZvm
hXke6rKDqta3szVZT8Km6MYHGcpCy+vXqTNB3PLNu8Yy+BOdkYucsYalyuEd7JXNc6Dz+pt723/2
BK7rh/YbEhP3eYy/NX6mTBTYWMtVDdNC3aZ4500ANy4kVtvTYrWZN2IqnYS2KCF/2w2mCMW5KH1r
F0T5SY5q8y/YLLIySYSXQ4DC3/fbZK+kdexcTKHafQJ1TuMgPTWgbqV8+Q5RYjltotI2vdE9k5LH
57iEDvmxKldxebFjI8JIziwbIIJdPT8x5DwAkbfL+/1ivgQjhXDCXSPkE6gW6UCnu4fxgEImjyYr
A2pEivedbwBFeOO17m32jFN/+11JfTAVqNA0gUnVRYEb0QCAwH89bBJLBgoZs5RuO8kn+7p2IaZP
KJRSodt9is259wOInBb1mzF19QhwymYCYukiRRc10Xyd1ncu09PCILMQHf0lfQ/ZrtqyHV8/HILc
Mub4gUq5Fp1P5MxlfjJgKGq5/KYwwi9vxJuCvg0y6YkZjRs3gtm6YkXHa54VFnyeBhksKimZk9gK
UMhoRlfznbDZivgj7P/LLDBqo2KxwSK9EZOyjnsNSU6ihFrvhHorwRmn/BG00UEZxzGj/hkvP+ZL
iI8ZFrlApYxeu+NsHi4rlyjgkZu+4F62vpA2TAGq0HREBD4cgJ+Ja6fiDrQHYog2OZTS48tJ6Fva
2paS7swkHjn/Gr2JvmCZXrlqLIDf8pdICKXJqroLo2ZlWCf9ob4ERjPFvtCZbmoNXmfA7RuLV4OU
8cgOLbt+QmmOMm1OllcmCU5j3Bbb8zfd4XpqSU4sbmbThkM1ii39wc7GA0G6VbL74f2pG6FY0QKK
jBJfgnvEDlUyv908nEatRvUz+I436eIazkwHh50FZsJO1Feu5L71Kk8xEn3eKjky+p/akkzNCueE
Pu1rbtFv2Zabg9qIE6iC6QRuxRO00gjZnkSd96QQdKdm3yspWPxNxwM4IwqU8oYrW2zxgUtUomZ1
3Fq6iWLWmQFxGUazToPp6mq+Q8j9w5bRmXx6GkBmjJX92gDRHg3x71R8df0iideXvCV30dGxpOSs
oYkmRClOg5XNSRJ/cE334szq20BZFaD3M1W4ehyiiDpx7CZIHBrxeFwWSBELtEFS/FwrDskTEJZn
IF1NOoWO7Fy4hCV45w/7PyTBiF/lFbQ/zidrpbdmJCaom3aOewvt078uZaBWyjfJ+ZggS9A9AS/q
b0Pu4iSQ/sotdTdL1+HvjrevWq5JpAR0BSyJZ3Au4jGKc/ONJXC+i11NzojCS/0OjVIq7XAqmfcA
HoJwNvXU24Pq66S23mY+I6T64DFSgvamgWKjwFA62Zay3aE4puV92XXEGOMreVUyBv9TaXeqNE0I
TrRPYiXsF7sOrcTqUfmzLxynfHfBGOGsWdxUaJVaLxK9zsdlMAI1dkuCJCQ2jzri4a4xpjol8dCF
IAcSNNl9Lo4zqjeuMyyWdG1PE+2npjZgsV0pe1Qe+NX4WEx3MmDX/r3LjiYK8yp16DByQ4OmQzvv
9wXWGUu9E/hv5pw+dgTBh7NL4lIyj0piXfNqjo6/n8wvMNh8xP5wRzmeMij0H2MLS4D9E8msiSaO
QC9uWuOPVEj6C0mTuhKgD4PjDEPKXY5wGh2VGgIVKvhIinl4QsKPP4hMQZLN7Tj+QT5iE1nzcQHy
2ZQxvonj1htM6+Tesq1kJ3/W9FZyIK1vHr5Tsd3JbZTP78sVM7Oo7zHoBizIYDWzbhkl5O9uY8cH
cDIWEJrk/h7u7/H1VBmPZ1c5vTgvkee5bVOaRlHQClActKepMODv0lPvyMnbKF1c/RY5Ydb5Cv1V
OCL72gxqVquFofm7BpVjTdDNd8ZJ2x4woRxPhLhMeq8eGgD7bSs3z7vCUmvr/YfKq+bvNgRRxxOz
PpcB/pqjS9osCMMEHGPWac/R2ohGb6OboJi9fajX6hmoCnvw2iT7YBF9AxDJz5JdR5VRmoH++fgt
8Pt4O9lWl/FcC4ml1pXi0XMHm1llmJqe69iYKJQKRkgpf5yDk3FtIbz3xnPa2IksL7K+eCejoHau
LVVaRcwjOVIHBgAsCCNclKj4Rj3bazDFdCf4zZF1MZ+iFgh+2I5QZSh6XA6y9uJN6LSJMXPvDGas
V0+HOhkRW4wCW/Qv5fkP55SGx0hcvaVHew7OQmBXS2O2SMO3oWdem9TBoXmswAu9ivOF0oxJL4R5
odIhNwFMgNFkMCMbwgesRq+fTfGNRHHSk0KFGhGAD1FZJLrYuEtbxzDbiiiaRv7pu/8n2LQr3cn+
WgUBUQXCOJ6lNfc7xDozmL4bOw8KnL5aOsOgghwKeCQS2c+uYZfCyuFRCo3nVWqtBOoQhCEA1dYN
hjPnI19sYlXUalDfjCt2QCOJxbKSM8OIP+iv9LilaqWIJsAylmZqYSvlZSFRIVxjj6coUESVumlq
cc58Pzsh23QUHK/1g3WQquok3n0h0jKet/vXFigCGm2YUsWcicW3m6Uii0YTV0xFPRh9PLNHmofi
/v8Em0ftwvozETCLDASYIKYVr/Zp7ngy6TFeXiMitfPUSZhlykS35A5D+SsQWdff3fQtAlBiLeTX
RyAFvWNbmct4HMI2S8BgnaIv0IPUXrl83dlNwmP6qA8BzgmaN6nQX9JTaWNdvLsx+BG4JgEjydPD
bMEqKsRX5Zd9ugdYF6OjSfRG+rEl3vLAz/ZDm9uUbCyrcDBc6jC3Qq0uGuZq3PR5deLkN5xseGYn
6wr/D/DFsIzS9PDZ9CDqzsMp0o1ayerJh8U3MvTwUyJ6T96Hv6IPxvxkz3G80mahQzTchmh0vpC6
YyO39VkZuxJkPNCOFwCyshaGkt2iQi0W4oj2F/ObLyJieU2NMCFeg+xxXf39YUEFCPF+Kovdiwtj
pIj0xfZiHmxh/vdtVs/47BrZ94LMVgxsdm0kCB5AZapOOD0TLgWDHrNNv4lv7fRQWU7AmQ+BSItJ
2JZnVBoj+1GDCQU7LfU0R6J26W4fdEbhoB/cywMermdCD4dHn/FqSdOUNxhF5GhLsqiaLBf+ORO2
2GEBpPvVvLo6FVkZnV3W1WOpez8hkxxd/cWOU30P5pA/teaRugtzOgUoTKA/JKNbOYph5Z/GIjw+
G53V1HBaJmM11ZnbaU6u661O34j1Y8ftqbdq77il+/hxUAsb0zkv7Wrh1Hwi8PYXpmCXO4X5kiO4
vK4ZmRbTAG4Mpy3TUxu1BCZuOwJFxZRSlkkue6apGO6RaDEQzDKeEefqftr14Eo4knFMtJ0XBixp
Nt6gDbiXfFwzWxvPwXdy+/F9OwCziKt0fIw42+Z3Gx7CiiWBpuUn2INEsDZyP9bxa0sXHN9RRpYZ
xRdE2E4dkeZ3TGv1OKpa8YFZO/l4m6M76mI+Pe/L1NqVsqfTs3HtlCFeVgJCoI106KQgGnxz8Tnq
fDGwUaO4o16XuhVO4QmBZ3pKzrN8PLBp/C9dj15JTy24M4IIBpZfLySwQX7wDa59+h/ZPlNeXMZ8
Z9jqLMwBakjQq9oTNMdeGcsrP96RRXZnO+YOnEhT8WVBdPFPMMlOLumgtojgg9Zbn/P32z4/mTGt
TgYl/XiB6zuM6HIWWBu6Q8CkWnbZQ9KodSwrIsBVjYWIP4tUULIg1VnAnnlvffnybsUllCWYq+XW
IEQPvougX5/bMR/rHhOfMcEnDe1NlY1SmPo3n43KDxfPOIuamGrErkMFO14cm0FNNkkRsSmNquPq
8RX5/y/6o536neFiH30bKtRDAJlT4wLtAKqLJHllETIksczIyucv2EFW0NmF0FC94Uh13H7+NBRU
E0sk/3d0Hy4o5/2tDtC08CPhbgAkgzH8YXk35QRxtWzj/4dkXZb0EthG5+oH12o26gXxLROT+MdU
yosXuA4t2JVDwNTJ+Z2NUY8f0s1/xzKCj3LYYsalj1ML5Gy8zpC0BBzrkz+zstL+qPEFUQ+MjbFD
hB9sUUPI4DZ9O+J7QfqwYmytNHW+srzpN41yGj/h7REGoqLBv4qqr1UMWOwdzVR7mwKI/tUAhNYh
HYhX37HmLHxZ076TXnakq8M3tGCvITxqPGfZ4Q1wZJyyqC9i+kQRvBosup/xVur8gYc2kL+wBKwx
NDcbNLosnrtVQJKeU6zH4lzieiRcv6xPyCO2XbcH36toyf+cI4fimC1c0Lnn7rDPPgmNHHwH/h1j
K7E9argJhSHypNL7/bdMj2nMCWSwF1V03WutEvG1AmKn6swdXct+JAiYT/ITZ8Hvv/tJt0ChXWxk
A2anXLwgCJ4M34OULhAeeodUclTnIlk5qPdY3RAd9lUFJ6sOwWiYKLuMFL2lsn0Hu1jXjkJ7PogY
lh9DogxiMaCCeJjIhhCqAJKy+FKEv0JJlsLq4u/BO+hJXjkFFM+yzvPpEMx8VbJIeVx3kyPoV8L5
UxA1Dtz1qiKA7bsFPKYuoxqt2IsvjrGFSy7uVy71orvCOzMOY8HR5pdHtQ7+6bW3qtybkMwz4AEs
NGpunXJYGyPCiBlDYQ+k6eJvALdqNC6HgCHN9r7F/tht4z3nrNOXWY3e5UOcKsRKiqHYB9+WAhPN
uQ5B7BBC8cCwY0OuNHmIBcjzvpjIUP1SRiQ7x/HCe/i8VRKZwyeqXLUHphSqKTo5ffXBGUPR3VCs
ooAItpBCTm80B64kj1ennlpJUeMP2AFHs0wPV+/DunCBbOmS7nFI9djqA9lCee+Fq2fEE4WELAWF
tTSmOwdu8ORuQpi4l2O2XibGPeP5fMXXzGcNRNxvaME/JYb1KU5Fet101bFR4Ga6GcFhKmPXkiLp
I77CmjVq3DTFiSwVF5HgCrsemTFYKCOjl6ITQuiGnQhaYndz9gm+/BmjNOW1rCED3TXgpFx8o14x
bwouJyy6Sx9/joixe9Cg/mn+Ltb1t5x2m/OSTHrRt9h7dX4tgjIpkaWQC081Owi+LVyovQ8e/dLi
4DQYFYN+zyNF7XFujivStq6k2o6RjfuEMJiqMsVasC2klTqmXrOaC5aGVjKY9qXKiATTzWgGBV3G
OMEojhn4sXi6MXLdlLZv5GA5lENlkf2DPVWE8xwwDBw+ilPx2vh4zzL4d4NXnZpi67D+dYCn+gaU
Q3mdFsKRahhcURHynKB5x2nlVHlttK0Y5sbZDMb7IkIkiKa3JZoVjR3S9Q9OdO5toTcFIRVUnrIV
LfYbzdEI/IHBBLjLgkWNiZp4koiTms9R99QhBu7H/VabhmykOS2z/6nBlTuqDH1VOqw/3kXQNC0M
wJCD6yPj/+vPoX3Gd2B4/fCYwfD4WvXKrYBgFrM21mmLgLEj84vG8MsssjAQVjOoD55NZMAHenGL
lpOIDWWRkv+wi27tDtyco/zvkhdJu+MIjkN3aKrB08ZTTwL8BYY5Nk/XHuEAgt+Vf8zSS5r7REJO
d+7YK5F2tHg4yQis6hIHiJX4b6ADKKpmeMQFGyDQKEWi6hHQqUrgypSnOk9Ezz1xesJ8stcqaqzp
lKus7kVCFonkrp3lbrj/oCBvLak8tgk7atWjikZoiR+Tp5Z/yVMZLh5+ke166vV+QboQnKefhOAa
DBOQDd84/W7YLpolJR+N2NfG8svp61o/jUdbcZcE7mYwKKNQFyZJcuEmF8HPMVotKGto4WZwJBw9
r5J5H2zqNbJRkMT0NGPM9TfBzssJ4DiXr1TYFbCsr+/rEVrO4YRKJwj3iTsJAmv5j8nnmRmRONlv
T6hxy9vjWOZuHFTlO4jPR4EJ0egeH6wWErGQsYG9/fyChqiwClNQV075m3rRM9wG/I5ldXxlZoja
tm64czU8BLApPlGCqVl31LvzLBQ1J/i6FO8l3yDXdQGAjpCX57OD9yl4+DTC2QR4tSZBYqVCkHBj
eY75SViO5cAnzYGNXo/2o0Wq4jzh/QbzynM+tJ8tUzjJz9MJwToRB6oGTZs03VAD8/f9rxPjTJYV
Ob0zWj8ymZcq4H6BtBSUgJVtchY8pUp9sAeIam8nMQqpvCnraV3qAQ+PcUlV85BdUoUjrsngAXym
o9CamyIndeTD6wbmWsX8FbOeI/yNzNW2CH/FGz0oRJM3lx86yNuu03YfPIMb6uXICtcDvNJFH7y6
2D1UuGQwzyk0Us6OsGOyZSZu7vwSdKZ+Nw+11dEFoAPu8xRgp/A1HWg3cJol9WeUYNjz92B1Yt9v
DBBvjFSE8HVqyUTJDVfUt+KValFYfBh24jl9fvDMGd5DTz7XGfzL4Ae4Xjl3F2SF/6cZJIQo7oXq
AclmcrEdMAHw+aNh2/bQFA41YXKFn7/vxTe8v/HLx2ASDWHKnaTqMWyegPR/HKmUiqlW41kWdUiM
rzweHHMkbyLOAzIQ8K6GMs1q3xcmAk6dkFlrVFPMHe3jPduloI6k6Rg0LS137PNESFEoVVoMLora
F1+VS+kdqICMcOGHKp0gpIh7lkd1w9nHQyqOsDl8JDAMEJuMA6BmSTEQgs8Jnnwf45XLAtgXRKvw
LNsaI2VsVpXCnmpX24uOdC/G7DwqkQ2pGKoWNPRL4RsorRhj4xHxkiZH3WyTbEjdtWtJnHyietCj
EZKzWiwsA5zBG8PlCTwIbcvcp1NBjrz9+Hdwkh+rCV6r7VcifskCwsMUPNUlaKqnrsaEGAq0ZEl7
mcJ4Ofryyq/Go8ennF/ZfxLZblM4sCHWcgy4LsGzxShSBSNMxqmwhDjLs95+brMkOZ3+oPUV/q8k
T/dKsAhUBGgWYT5N6h+VlfmsP1gtqICtfYKGTxofoPVWZXu6GOzuD0sKQL4tkgfhWiIgv4IOZ0Ek
RtKh0K0M1Sh85qyx21Rf5QeheIVIRcte3DTxKja9JTw2v/oONhVCUl5wmvtnW7oJB776RkuQQMZf
oR+XxTO8TFhqDUqgPfkeRFUrCgY8ZXlksix+Ox72W+woD7g0fC6EzV0SrsOUTSdeohyrv+hqBSiH
6mZyDOJCPa4/FySAz6CUyRr5y3wlcuN/rSXyZ4U0mW1cB1zJL8+YKPymm43qjNARlA5oslTHvMPU
d4ya6OFzrU6Vb8IrEXRqVQP3FBdTffkv6JJ4itCU1SLFrYn/JG1FCUcjUuNQU+OSkok0gPTQCYz1
0PnqegR5tb487k2UEIBnPm3zTlscSzcokxu4mbJD/RlqTwvzIQ+Wli/0wzkz0GEJEHgDIZcChu09
6QMh4jgzWCaA0i+w8QQQxAtUvk0G3uraK7bX2uLCsFoa2KupqRQy64Th+xMY8k3YWaexX87ZrGY9
YK6FZPP7cIpR4eJBqIy0rZVaVVFTFhP+yeEQ3Wjku2+3AM/xucwGkLToI8mGy3PJAu3RlMuC0qAP
uMRz6A0HnJrE8NCAVp0LQhHdy43cPd2d+XUxm+mIfKDXhxhsOzA53+Yylrr9u1WgZXQNlzQJ6SYS
gjte4WQca39NiyzUpTq3NjXD2I+N5p8NeHmOA7P4+kio6vGt+IkXb/cctbmrJNhI8Q8jyYVyKKvi
J3lJrR/C2P8IDYRMxy0OZN/3Or0Rn6ervBnjuiOvBCyvloM9+mwOC57fEuu2uDoM28wYC0jB16DM
ZCxHHrVnFnUwWvOB/Wynm/DJH+6SQzvLKZ8YpO/YkrkELTmoL1/HVicqqAFxdWXjStUCPeuVmRIg
DbdDq/kIMotSQGr7iDNP+qALbjGPfEbC6gqxWH+xqmcw0wtPHTe/XkX77mSQNhjE/vx+Ex21Q08O
JC5EsUgmHgvq/CgpPNqxuchEfvgl5HKUp2JqlfnUvPlURBPzqfd+cL7ju23qnCT318eOMiKS95Ec
0trrwEMrLX92VtoNVAl5d9HUOZHuFOG4pyKs7k4ny26RoKBdXzsOtgsiD6noxevf5DCHjS7BBLPs
rwihmlIiSSl6ifBATHzplhWWgC3nOu5zQ5rYtULYtKhlsNPR3vLcNsL2U3jSicnSE+ZsMV3QVwag
pJBfVOhpPXg9Obq1/2H6iuKu99INOQ1DCBAWW9UFC6eiz2SoTkshm9PYNX3n06CBm/Fi8HHJ8Uq0
+kD1mfcO43DHPHcRhkDZa7y30KEhHjFot3hd5KSjO1InrE4BTBQoHLHvt0VHAsLpcWy2U2X9OIRh
I7+4FnokrOljW+S/FkWPU0h/Oq72haobwmUKF5SUpojjHcaP3rHXjTn6WwpiQiQMD82t4utW+Eo0
KlQeazE0GknTOdYAdoRGG+6iiVpB3ueCInba1QWRM6p/4Nnlk0DB81/4pNRb7leYxf23fhn8ALMG
LGNevfm205C8VOdgM/jM7sujgwYMOGGed/Q5zH6EeHLlSImWo30tj9nztVotj0Q1pFIYg6JOD7cY
tC9dfcgv9JDp7zGSVQqSbbSeTZ3+plBM2X1BPhPlCiUSX+0MmrjIoZ/BrQ+uu8u+1zMcHd7YPTMd
O1h7UUvEaIb6QHwcU5iIV6SBemSzob9kfV94qN5Rahxsc/ly2x31UkI8W6x8w36Vg6bJ4eW0FnTM
jOBKO5nOoMJXcf8golDhO3pU3U9iUI8qhH32EOlN5PISOhedg8NBrtxHTKzcHwhEm5o55+DWSH0a
3WWbEXQnZaozf/CIpXPG7GpWy3WccqlMqJe90KeEHhOS1cXHhIAo9GiPFnP42n51oiva2LeOGPOu
dfSce9mO93U6Ukgp/vcosFRIyGi+yGdGRa+mODnNY9bSSY8cT5LCQSzn0FTMlsy92WPbvxJeK+yL
0Vn777+4n2g111dfcN3Te9VlNZg6Uq6P/aDBnNXIIk1aaO7uT7UggbU9S3xLMl/xwMa3nPCTHEPr
03p7LkYYr7v2kzDraJjXuuJekM5UCt5YP8Hx+75mS8j+feXknZ/k/OWM1JwjItwpPfwZfm+4J7/4
fuY5nCTqp6AXAVC62EgGb2at8GmirmVl2IlEAZt5pNm5ioHQx6hBKw4pcqqGQSXuPVZL7fyGM1Os
rSyjUpsPbhOVyJUqumiAG3eWdX4nBMqqsad0dVuLWE8hHEPvMD0pOMVDfRBVVK7bRnzC1/dodSpF
67aJemn5eiduqvwMm3gEG63a1MTM6IwyyQ+BMONAxGABbBKutjbfsyqnQQLfcA9wn3yLfX9QgtwR
9w77cb5YfB8iciu5H1csbCuCWFS6JwbDKaQTSPHy80rcKFOB5ltTXtHhVwFiFLVXjcKlLiJ4JoVJ
n2Prg+QzP5C/YAKY4Um4XCkB6nagSeHUlR/Ple+4NAZzFKmaKDVc192XDkkTpQInkN2IdPrbBzVC
TzcSONh+LlIYSqVjAxYBENKBmC97UWtlCVhxYlhha93mFl80xE6r5wY6Icx2wqzOfrrm5L56eetq
q5yA6mchiZ5vyvnHMwoSQLidrYP3YFalcfHjGUyWNVzbh2VKef+X3WEmeTBkMSbo4f1Opnk/805/
0Z1hbLX4cFIh0QylIYptC8FoWzVXC43WX29hExnrkxUdqG9wTqi92SPtk0nEwqy+UZLMGZN5h16b
biYQE43ElSCavO5ofroVg7haMzHbL3NOC8sb3ujcj2VUDBhGeJynGajKD3k4WZ8+F+uLDL35SPvg
ucabMMAEsKB7arEMy7lJ+9TgvUXiNUcqEhSaY1QjI0KE17dDXNK5ERGvo7H0IeF+I5UM+9LsSLdS
OFWFcQ2cnyero7LRoBYAD6JnoHtgVRyAlYbEv3C9PpXn07oGVBhOeQDgXFK+A5TlkJQ+ZEmwnRQt
/mgCOtwqgCk4xyx1yeUCdinLqEDNmX5Goe7ZWO4PYj5DOOCx3ab04LQ1+bdYmGFfOX2Do3D8+bD0
XuPUpmKUO015g/SFQ2IC4coF/LHbm35SvtIhkJCTLEtiexl73+Y3ylOX+w73l7APuJ/XzHR2P828
I8q4VR54ZWEgnoo1J+FuBZKao1a8BTPgsQk+Nd//DpJn3Ri6Ou7IJeODhjTWny0MptV0n5OdS1qu
WELQvfcE3wj9H84JngivHmRfdb+6detCYW4dlX55N2xS1Q1qbAmeb+mbtGS0ATYDPzwUwIMMf4My
dgazdJkqCvai7qDOS40lYoMwAGhwjOFp5HhvsNNHa18JpUivS5lDZFupBdxGVG8hvP9EMi6hirAu
4p3JsydIDa2PiW0pyFu42GCLa26Oc/B3muN6T8iY6BuxSMz0PwFhOWHhCeHb/wijZg5BI1JM3ouU
cWl4qNUbicnwJ76Hd1r5rrt/O/Ih6lW6w/UZSp7QTTdlEezcizjH6TCJ14kSHfNRIIdJ/MNWDQcN
eBBvQpL0ckSqIxdej2M7VI/EfMExXRoWYlPq2P24GvFY3NyjNihXjXL0v61bzTvj9lDr+hLvkROd
FSJEEXTx9SaqgdGWuVdiIxqMEqZLe3QHMCYAInElnyNgQZQeECxtO1KXQVbFob3M2yPsf7D6qwIC
oz2msMK/H9z4jEu3/JGLjg7wOdg21+2Ys2fSslMUm+PaDtrnQ33rtsausnMDFXATs06S8OkoI5G9
19O7EkR4oz7AiHzWE/Ix7VyIM2uWWaACYXIymIuryODTP85lB0Yyje7m3qI1/+oXoj8fAiXF6Y71
50g9Lj7/MfVeoPR/qRfIpC1SRY7n5JSbiaRIL76OzbgQePbZqbRk3BpRy6KmCC5K8Nng7h5PlAe5
s7tpN1rpbjPQnmSaQ0bVRQLb4V6peEqSx1RNeSa/Wl+QkjqimjPQN1QTbzwQ9sOOn/HRm8kiPh7Z
qc/fpld6Cq9QkUi6QsJIXampJuVMnQS6cb/f1GU0JBlAydkCQtxsxYL48iNhEIntLc+aSUzCm0kn
7VZapLUksgaSc+vCbubQwSUfZZb7JnQiNRgYsVmyjizA3PIrceb0kRX+XSxS5tQc/A14dUC2hF/0
dbfoWVx3idCDaKk+UVbVwpS2PLHE9iPExvL5SAtNB1SpeX6Ui8tsrDUcSdJIgFoRnhYsfgn0geEH
r4oxquqCepGiWGbdxJAsJ9VuZ5c7lK2Igfz3d6XLw1SKDxQqpsFj3B39zkvhsGS7HnVI0BNViWf5
NQ6jG9siYM8StXznoNiMi4fGocFcAAXNSZKEqwmOQnn1r8+eVk38pf4KfzI4yyEDUmbki5N43q1N
i8ih1mdGu5Jo+KuiWaXzFu7I6vkW1nvfidFwDq96JeS7hIt+cGPggbwUv7orstACr4mqvo1vzl5I
vKFoV9lpl9MMVJ8I9Dv/E/3s1EUApkSMLtVI0ANtGFJ9q40BqnN39wE+tkwuCsrFIyZDtznYErMM
B/0vQ4/POvM1/x35QhA91MT66WqejM9pdH20wicQKh/IhpGOAJl/Z0Q7iB2/oyzXEnOB7Z/bekEQ
rRCc6gD9dC6Apyf5JyPOBbU69Tgzkpm5Enawh3WmNRbqjHAA38w7iEAIY+tkjDtjhiT71XMrcJWK
Z91GtNr4+4Yt+g/A8EZPM0S9Fu3bmedhgtXz9JRYtXpmXqkmehZLcECr37ADBu6WAAx4/8dW4lWq
90SRSbd/XPldqNfgTrII4XoHMSwHxCEu+eNIfXX28hblybyewB+ILzqmRR6/nbyLYNsmC7zPzt42
9ZIulDhKfKE6y/fyh12gpAwu3qEQu0XQJ2YtIgYqExWxggWm9RwLaU716JGA3LxiQUrsHUgieKWY
76ox1zsJmzpKSdVU//oSGJ+RJTSlPybkyGOWdDft4FUUvJo5u4a2iEQrIaf5x6MvTwxkun95OzSY
N572+tgU8+4vrCQqDpU1NTtRGLClwVOy3xRJtIdim5/kHhtwD1GFal4Y/rmiN4aaOoCNMY7eKBAp
YiBm4IbpzDSa0wX1p1Og8YrQwc6zGc8kMOt5dfkaIyB07hGtkGHUPAH95d16RUjhq9I23wex3gId
7CvUOalOig3BO/sSJ6cH/PKjxD+SSSSqLIy59vOC0aVYaqm64PZj4QITxSA5qz1aN70Y7tdcSIu+
ui+J8/b/BIF6tnXR0FnCh3iE44SDTr0cRnMZyncsNTnO44vJMyH7ASNViLx6ZDb+1r9Fj+5E1wO0
t4coyMxuYX0/yfrt4A8IofDast9WL8sSyVA7qHeCkyz7K4XIzc60qShCIJtO9v03vQa8+JEsIPZW
fYEUlQH/SGmUzLTO9Swm4W0q74MC9GX0Cuw0ECc8ZFiOesrUuCOPSiy9ViKrf6NdIQ3xtAhzMEz5
KE/h+tpEmxIVTpu//Cr/FEJDuntm3yxY+gVJ+W6pfuBIxfZErJS1NWJlIRaPdUJDyN1x2Ic+F6jb
6n275VuZl3DpngI3NDZeJJ5TbjQ4fiR9RLAo0KfZrUvkDN+QUfkDEvdg785WhjoCc68bBjhha00v
hcXpWavsfPjONrk4Iw+Krf7n3c44cG3sCxFRb2QAMlq8/97mIHWSxaC8JtHqSaug5EfDu9EOUb70
lNrim2W46MqxwBOEiHXey+/a4iWADBrhsfuOg5C458XiwN1/rT6b2Ek8C/3p0e0Speb6JXvIQ2HK
N5VsCKcNg5NrABBMMbGWJ7r2lbdqUH1bNbiloI3B3YOVZSFCjSDmGZ+LCIWMiMuo787EOG+6w+gL
wWdjnNvmsoLLvJc/70vqjMZYeIetKm2mwRNg7f7VRRavOhfdDnbrkuPbasR9QATJAPONH0Lwp9LM
BQ/12VGfoBvlMA8kl2iBxGBUAe8bC7BSI8vVGcu34gpeZ58c695wq7yPiFGbyexMGKB6jcD129Or
6MkDPCwX9Ba5uTSeDto1m0MJjct/9gBw0xLgHwArpeMgA3mqGNjRXwswCCjZwoWQ9NWInBAMhNdg
PsrIF4QJmNyNV+bM9itBlgIRD3Nn4h0Lka1GGNk3GMl3PevlsmeN3p1ydBtvoXeWCemxGYU2320O
ro6HWVBDEaLvaA/w2oTly19rZhc48GMlLADFrvqVDklSkTjOmKLwJ2gloeLA/eFR6/3fEEt3KEJ7
yTnFoqWRiFoJ5IOgd6LkeGBGZA+XWKPEQEbQGCL9P1F3uVwJ81bAr1qgS371N2L2kaP0PUsFdEJF
lB1RngbzIiPfNFQspl9HCT3UWp5BoYsvz1df3XVOCTfVNTsGFLu4sBDj4JjbnrcGH6rzYqK2PtsR
9V8bSh4kJQzFV4gpGmwLNGDbnXFGleWorkVx3QOSvZf+4a7mu7swohzIVbRecW3SKCobb2l/Stkj
gEvYg9HptS4sNNIdm27kvXoGVJzsUL4FzltVzs0N3l4nu55YESWVNTM4TrkbMeZWi5xZwiiZpc+7
MgIpNUc4L2L1FZfqipmk0cj8nlfsPzG8vS61Cp5tpaewi0Sao6LZSzeoASel8jCmTigL+Dl9bXuc
N0dC0G0YGqim62JNPcMPNbPq8QE7hKP1e1Hnyu1xbo1nW1SPEVf0WVwhe/jB7tR99gZfLKIq+95P
FeY6Uq8rXmz++a6pOCN0Y59s/ZRrWaYEvvwEsICMptVFyR1AECX+Q0dlxBItrt4czUeSStJhmXa5
KN3iy+ItJC3TV4wS35F0D3s0cB5TjldIVA3blkQ0t8S5bSnZRhG/LK6OoIXcgrMEv4/Uz+Oi9R9J
02dM9Qy/CJqJHTfkWny9Iy3sRvfx+hcHSpbD6o7hZRo8APefmpmBZuCutQSKnh/5xTAIk/ZOpSNk
3tMWorxiuacacncsRUzx2muE6ojvdYupsMJjC9SRZ4TllQB/VEwoW4hdQ/NoH/Uaf7Li2DA+Cp1M
iZjHpfDLh+MncB8q8MR2vysSPpX0Uu6EJndmbuWy/hcCn5aqRgwjKjVuAOgBXKzkurWo+9AnHeFl
buxQHens7y/mqikmrwGPV4us3gZ4T5uxHYsTxMeOEf4EYCrWpa10DFgwYvJkPE9BM8RDU0jVAOL8
MGnKeSebtiynmjNYZxUgBKyEB4VYODSeKgQxIG5JEcWHhPwba+j0uC9uUYzAsb09MiRdOGu+Vqz8
caE43aXXUFi33YUkTwwppjKA8MS3aNXAtc9WGZ8qAN1YXn3rzyvV9BiLDzKNmPfWTjWFUQqnMQk1
zl8TeRncSLR9N6fQKrmE+pjpsc0KAsgo9WeitEKGuD9mcd7jKM5KQxEgzK4ctE2j9YwB7OCYSS97
/wTTqKcxdsn6IzfJOGsgjmd3EKAdTQSfRS4nxn29ZCGTDHZnJEswq8RRXtmxv4NbgFoDDrI4zGKh
kwcAvHRyjA/u4eawsPMedFpMiw+4gRHJVTMYCOpw+ONumQUl0MCzT6EAWgUaqSuIb3MlQg1AMQr9
+XHQV3QVQ+MFEOQHEK2Qkw+rLJuWAfPQyHQJ20IufJfAeHJGywq0GRAFvUMD5RHUmLexKtc4M3ou
12aQ/sibYuuEVzJVkaqxu2Orkfv2dE96o1JltW/8PnVHPLeQ6H0wt/ZovmETXlWgRZ7VjoH70X9T
eGkgcRkONme5V0I/hqdXImNAkORpvtLebj4ZMkmHvnjQxoBoMYSXz4iRYF7whB6c2Zlmz6MNfGhF
xHe3hyEnAW007mBYoAskJzHRsWrXFSJIylapUnNTja18FCYMXebTtxpZVw1PJnQ2PRQapCM1eFCK
t/aklkb6yFTee0nd/r8y19l7Uz2TucuVL//nG66cUlDrPuivqwmj/Y6oZQ+sPr1NSI0PkQqPJil4
u4fgonTUXySTxoHZksBtFSeJ7deTgEdsXi9vFGfqrqipWyOkjiLuVshAHJSAerwAFBqvMqg3ac+C
tJB7AeET+Ddfbn863woGweEFSTIU9zm5cHaW3dXGBaUctZjlfroPsHIF7VFd/fX9kItO2CBJFg+I
WD0fyR3zbu0+XkOUaz6zAYRW3EWZZjRRcGw9TCqGwnOt5eKJmGrU7DbktdxiNXvG2CRvxK+zU8OR
C6qRFm9pMRsVjzj/qAPqZw4AKhM16wAlSMuaVZTtlr2WNCnR2RpbHGPX42oiQjIwaDjnIeVra+J0
b/0Cfhhvjw+8D9IaN6iWyQ43X82gis+K4oaISum12ZFL0OIwfKflUQRXx0qtqs3DyatWNcrNfaLa
C2K+wdmoSglgR64BwMNzaQXh+rBjaoXV6Vpj8Y6GOJw+QjdktTvHW/LdVEWqX5jiHBw2CZwC/bDg
Jx/U+TlOtDochl/CaInVwyyYL8IshVX4fYxOEPb/6UWEgX1dxDmWex8NX9MGxrMn1p/POyAehFFJ
7ntK6F5YPk7fjHHNq8Yra8NWWDtJtX12ckHdgRfvRX5sO7o3+/EsNez3k0SRLGP3UJadH8J1AKZU
iE7eIImFT/e7VbC5cIH/O0AUx7FMNtDjbX9tSAvi+pVzNaPNzKQAgqqbc/G46evsNwQ6BUu1PrIo
0WF0W+BJNB4U4EAXeEwYj98bqM9BTGO0My6PkCNBQU+Qcdm0Qi3Goq3lY1i8QLpmiN6/BrziYMTV
jo0nf8cIjGsyUtjtKQaCGV0NWhTAs7SszSJIG0dEHZVWuBTeCzR8RssHRq9mrIDVKZQW4lpHGAZc
GAMt2n3hxsdaUxoNLD0LDW+9PUIhCxVMtnrljHpgwZj/OhSWveSaLP6EQWq+MxSBe7/7q8gzne2Z
xoZqcxbz3/mYcVyu3w7y4mC8ifGvTlqRdh62kNPXyYEjwTjiNVsAcB5JhVXD48MMIyeVtctA+369
ZPDUjBi8YLtU4ingvdAXKp9aFA4v9E9p61g3SJ+v85cC07H2Z5hshIRTEPARFfm54Sb00+5w1NJq
uCvkvVI51OhnTosGXxnYiEwFw6zsHRKyHSOE3ICjPMd/KIZgAByDcBfdgRPycrPHLGOZNiBwcPoC
koUsSNvB9AiOViMNLVJVtRBR3id/E06vOWKHbhe0BOH/NgPK7CVWrEzL7khS+xPo9E+DFuHoYw/S
KaTp9uZ2WUeGnYkNownhE1fJjgPRe9D5vNcS6GA0L5ZlHS6af5KOUWkqIt/k0qmqqDUHMA88JUpq
aL2CnaajbbA6Df6BUmti/KC22TzCD03XAlWZyMHX0oIWxy6xVF1Cy+REZGnvHdNoiLgSehKgCuVj
U0Dhn056z4gLu3aJE1hymb+ZuiBLwt9QwmongiYfaBOljshMYAhuPPlqzStqBlaa5svjKmeLgzoZ
QjFnFJd4anpC2/AoKxacR/YS/swUMsrnw07EfIpaBOoTBnQn8j3gJDAFy26X2//GSSdkQIeMlGru
Azd17YsybXKavLTeNVO+rPcVF+EjIrOU7QWojOpaWT09nL5qHhVt9MWEREBHc+8+k2f/C6JZrI6M
txbd0A/jRi5j28EPm0ORXilxjmcSmUSrM8ukDJqFhKVsjIpmUmXzg2djHUFdOINV40X644x14CLz
4J2bO+kaz8KUfAuvmAUPkxtfVhvaR4/fdiFTOJ91uqZQ4a2NNedJervLNxdvshzk4cZP4QbM7FFI
ReNl/eiR2p/ysV1PA1hFSgtUE0scOK9DphLzs2zUI8UDbv72fuuZBDE5YCP1PG9ckp78UR9FmJCG
KbK+TRXYdPQbAh0O85sVG2KRLwKGjSPITxO8QqavS1Xs2D5Xi8yoj00bC0waWA9cFkEf/TZ2r8j5
39GJb7oudUOcALDL8xPCDz3rL/inkYoLQR7IwOdAX1XI7ty8EtNTnqQCrhboOAw6LxPL15MF4Alg
QMRls7UJps7T2UZvCf3mV0W6CDo8StyFP1qCufW7kI1XM1ZTMSCvBa92dSHZaWLA8IclK7ZoNtWf
ig8xvzvNidJTi+yReFiH6Ml8mf5EH0WSCl9PD+LB8vhZrMz75R7hiS+2Cq7EQPYB2T9XmBK2eIKV
5rXnfXVKpnsTa5CP45UJ+RSZ2VR3xqPqWl09z2ZN6nEgkXfbUdiHYLzm15jGjrcDKRvX0kaamzuc
x2fODlO2cU4ysb7QU8UgHPCCBwZRiDto6+8abVQ1vLMP2s1kByAHQorz7t26hQ6X0iJxM8aldcuN
xjapAkzzUS7ozcIlEuyCv3MXrgn9x+d3WlafgA/2KMA93y6LPBFhXf6Shq/uP+Gy3S54oFJWNaQY
oETF2JPHC0fciQHImr9QT69JkPfBpUvnD1X3mqeaGvPxKDsW2RVQGvJxANoUlFJjTReKGhXpYdsW
A6nJTcv5O41FHEelaliZzz9EGzRr74flxqiDyyTbrsID75dFq9bqoRhYfn18ogGRl/mWD3ORKPIt
msajrOCWxJqnCIbeBkmuLF6yQ7joUDXR7hXPdh4IN9Le0+ZoXbGT7r3kGrWTHlTACxTOXOu0ZDjM
vlLUEuy9MJB9CWoOP58xPJsnTy1pkZp5NIG6biyOfp8xkkjnAI+7+LVJYWzRRJj3I5Kn75Vc7xwI
gzN/8iBd7nfI1MaQIFm4ndccVeLEXVMw6z5SoZwua61VcPXaZvhfR5VKRtdHOUtfIT/a9z3OfnlD
ztY4ZV4VY12i0AuM8h7wGmrL5p+fsuBUTtF3GRmdfjmhpwK3y6T84+k1Rg55RkC7xkRkK4PaQ4Gl
Alzr2HTQIEE7oOuov9vD153hdvmYZAbUCrOGfgRPAIdHykmkANrka4DBJ0cBg7g5wp6sg7N88KDD
GFW4TWJZr61bc5pwIYEz76HYN1dmjUMMnASX8ZAFsla1jKM0G7BFKTiJ0oJWbemkxdA9onrFtrjT
S5SQMYSjNjDv6/tafoFYLNMkhsSk+rCsDZ+TDk0yz/ql6FXHIDByUjBiZkMzbHXizDlnis0Wu/tM
zkXjtwF1wJZAkSvGWkgmvn5jxVoo/WT2D9N65/iC/ja024uFWL3exKpROhkhVgXkUrS2tW/x+7FR
mTQWurTCOs8CveVjLvptkaWNKetQad3ixjC70mXEhEgni0KdCqRTLn22eSdMMe2niOf2BL9CF+Fw
1f+5cBXzzIQPNfWR1jWALbn9NzFsOwLGoalN4sZIzjtCvMK0FqVwdqkyukN5M6N9HXTmoyf+kZSu
ZD1D4g3BqfyWL6NUAzT2BKq9CgRDFkWEnNzPbD5ckgCKY5g5P5chbD+PwUOfpvwq79BaUQ4K7c5/
0S/dkA4jKEHP96NhfKepKrw6d+2lrEN7TBnM3mrZzE/8waIggFZ0LwguiK+AnA+YYv0RQi7tAvCr
qPfLzJaP5SqZs2thPlBYO4SEQaoIKouHmbaFyNRoMH1DHccAAeWzZ9VAFFlQqXZEeB5CZwoPfLq/
yjrvBCLGTbDIM4CgL5Gyrd5acxwg58ZRSkRJ+86EEh1MEzCGUYLbr07Kh82/D5APXAWP1ZRzI/WJ
/bjQiU2loNMEjE9cB1hQ4uB3HbLn5Rr8X+ZuqOskuyDUh0wPqPHnQ6sfVdQunHczy3n3NUTrWEdW
7FE94i3B1lzFolRQJKkki5/5+cvCUcIvtyGXqbQpg4nrL9xJEzInpwCfPdT3s8F8ENH8Hkxh30jB
iVv75ogg+Mk721euXGdoMWHDoY4rmEEu1S46jD4KEZ/KZoV9oW20HzDtUgr5MK3LIHmYKSxak9yL
wHvP4O1Wv70S+Lf/uJOcuKrk+4GjWik5JxbP0/8B5x7FuWsMXPQs9A5/geXYZq2WuGwtkoWA0AYX
LVIK3sNeriWWLGr8qSXz89RsuelzsB/J892zRJHNEJS9J+k48B9gO/ltQ+LMJicSp82caBklRR3o
JXrXa1pGZV+aFu+/LteLnbjj3EiAYTmHPd5j1yibSDE7RKTAdWiBmdxr3jwd/CdksUDS9vXdtjaP
W92oiLp7F42guN3VCINjB72V8Jyz9u0FM6FiLyXThMXvbHkX2Mq/cufLr1Z2fZzAoaYQVw5Pw8Q1
n7lV8W/62Jw5AyMUgRExazmkqCDzbsUbKxKhFXuiiXviHIXy25vTL6qtOn0Woo1xeXQegA3bgUde
5aQT/08VYA3VJjSn2dAXCYLueg1SKFl8h+dtv7BwyQtBz7Os/vfc7+ztC6DDGbwU387HoI4pwRtA
+6fY1/NcC5Mo7sGvkldDzm2laYSo0uG21DCVK/anuzgvX7ePjhtoABXSceTNt9NR+VSMlcnXLB7d
t6PFCwE5u8ayGcwNXIF5k/ywKC4FVyg70tLR/Qyz1mKpo1BOsrIF4T50OA0RgWvAjZE1LEU7MdIT
02mV0f7xnTIb5sKsgtMibP20E95iN1MWXttJGAjVJ3MonTAk8aAE/eCZdmG4z7+kc07eIzu4bScg
0ilDWiHwPxECoIGiaMRLqHxx2nlJ2Tt1nf3JM3ejukYxNB2w3O+bmX0W7e/7JL5VsNhGw1VH8B4L
9OEXuIZTazc8mhUCRJmBgpO5p3aBefw53H+k1gaa3wHGmDMfyBAjZ9+DioEyTspqyZu/066JGc3Z
iq+ccnIKfBTrZakMVnThPZaeqmdrXiE/+B9qtGYP1S3LhPJ4jBkCN1++4YFwTMhDISgQcNzDxe8W
3XuYLD9aWyWF1Sglk39KrYv/t4M0DDJHRr2hjmYPjUv7TLyRxcUjY0Gn4Jm6Ryy5VdLXSIvbFeb/
Jp/rq0Vf1Sjz8x57Le73G5MZZvp2fAjglqHAk5JE81yGWcfLJaXbBxK9nA4vcfvrhOF1LXlkUnxj
Qfavo+4dZQ3IqLsC676TduhW5RVBaEOB+pPSfmwSmus4APGppb3kZ5Mm8s50CDZ6aokmjE8xEObO
TwnFc32UTCiiXoCrYuu7rDKD9L0usAzoxFakVZi9RAogw9uUBlGQdadRk4C97V1K+fwi7+rh6j1J
ojEpyXVKkta9YIPhNpVT+mLEb5+LB1V0CWS6NH4Z0kPN0ea/HqoWQz9YvMPtQ53cKK1/80T7xUVl
ROXAGO2IJgVGuvejtYtSI5V3vx4Hl+XH4la34m8k2vNwlp4Ny1ctI+dUZ3D4QCSl9JWZ9nKS7AzO
aouy+UV6oN7oOeiDnQMd2HCAHdFVKuH1CEH6R89a8tPbrtsDKMgIyWYrxvE2a9dBmrWOwPjA0eFc
fzDYETABpek6JO9HLeuvx39sqPl/4hc6a8Ig8I+c4p0WyUkV5purWPrY+Itmiz5/NJ/dJhCCMyfo
iIdfHxz8IQNijxy1SUHgrfAzLVrisCh/BC64+fIjtDtYNZAiiH2WeR+lIKzdfYRtmGzT2r4mzNRk
Al4SZMCq7K3ZiBAprFw8jJHykQvz9XcpHbwMYH3ab/g1fFkcT32OOi93mBGszMCrFOhaTM8F8Gl8
Yxhl8ae95YBMpTkvm5M2tQrSb/VICQuoEHNP4rzrVwKNOz4R9L8ogE1rI16UFhPLOPn81sfMLpTt
bxsh5EzDMdPvdQUQXp6HQXOc34Vt6gztw0KGb98zHDP8qE0i8bKkocMR7oEki1MEKo18dxZx50rq
E8kG4k2rCuA6Fl9lM0/WsyJBTJ9AD5v6A0zW530hrnXZ/uzvhIWco6kA0MWSubJ2tTByJkUHJDmr
ovJwBfVlUFv5jcosl59pBudlozEWbs/lTrmC+BO3UzrjIyYoOXvYE7Opyg/C9eeGCKZuM+TJIbgi
30vXMcnvPudKtCt0V+LAy4jpIsqrsyj6mTpf/ydwKmzCpAFxe/3iauUjPBd9r5ZjWtu4X0cpat5P
zrYLBKb/puGjs5fnlwlP/4XrI2kv5eZmRajifpjqTmBpzUtOLwdBAE9kpVpFk7guPa8N8nGqh22X
lUi2HbFOEfs+vLWvk8EyarQ96Lqx4n+t9D1PJSwjLwdmV4bhXn92wMBwxl5LP4SVOtfWeEbz7QsK
6052Z2bcDWQyH/oi+iQwiotbqp4I8x2e3G8hXuN6H/5GhWa2L/xdRUbK/QBIjYhzvcrsKZi9UgFh
5Why770TnoXDD0V6CGQ/PXS30I7xV6BWINOLE5CWuoRq4E7Pn77JmgEQt7a1lXZ0TtNX0mtuvZLC
riORtNwrbATCZSX7mEb1391F4wiLIpQwW8C3gAV60qYMca0nxvine2xTC/cj9VNONeaVzoE/hQvc
JXt/BA2mBySnaiWMh1Y267WxKdQiWz9tk+qy6jHzBfEmmbyX1DLgp0+emDSFz2K2InFyOBUBW5RN
dQKCRrcv69RN6bjPfZtMRfBRkQMPezOY329bZr5HZzDZFOxE5CyoslhwxNIVXiWdy88vJYEn30uT
6QKZo4A2SIiIyo1xQnoGxc2OUwI1e9tF3cRXS9brmeo2DusBXp2e0sIi9UaDRF9+uGKGIAGD1ezc
i7u4wbSSgM4tdaMGMzZmhmrMnUNHQZTmpu9xBc9hjV0FFjZgSM0rf7hdNal3K4gEWjNSNHk1yynd
Cyod6gWCnQ9Gud00d2OJS+DuwHu9fTWZqCsw03MLi8spUFoyTnKOsw4ImZCbVHsdibeVH5Mmeh4f
FN+rDCUM14l/YPrrOlckY29wtcCGiV76zJ34OatbEHxd0NJcohuPY5cbx0OZZH9fKYOif9lA1Mv3
e+RJro3xoz85T07njzUOoob7IYepVfERX4HCV9B5cPWNc3R4/YBpqawWbdW4QZ3B52veezotz4jY
iAlJrBxlSo3BlylbwO1H6W0Ogs1ozm/XvLh5hFyqR69gd9xqskOP6rl4KSPPhTT6q4kEwux8evFd
xRwu6XMHtLl4ax7ZUtDjA18JdojZzqC2YKZmeoqdN2vNM4C0jQSHI91yPJye92MIQuv3XihiG/qJ
ECTE9R76H8/uAiem+3OHR9io8xl0kUh8oyZEHdYsLziiEm+tRxjFp0pxXhioY4LdzYfCnH657WXg
w0/mIU/drcsWSKCSuUo4xuwDaB2+OIfqZSx1EoXfaBjNNxkfFUArzJSKwjD7YOWhRRCVZZWpliDv
hcbPaz+Sjv7bLsgMBIbE33fatKsGQ97vWiYpH6pHUm87o5fvvo2R+rXHorePbK3Kk05OviWW8LE6
3q3vZ7K3SXC8tm9xCkG13l3j6PYKFyenD36o2GW+ksi8h08WDz1UzyzupZitvKUFkczFgcDp1KIZ
/a3QEU3FGzb9wdPysWR0jPmDh9UU2rTQJ65A4urCKm9DnmyBgGqHn/fDWK8ubRn/g1NgiAc4gwJO
MBINCrEel5jYkNuf8G97U1uUUooK1HSE6VFzml2YZwRSiNExbpI+a48D9AZvQ5ASdVglqCnFgkBg
KhJ8pxW8zt/s9ZCd4rN8p2s5XRZTaQOUnofHBdmCW7+OZuyIw3VKb++l9s9iiyT+hzjCWIoKpoIl
E3hjEepErK35S2jppx8VPazMv9B6ATddAAaWQiAj/Ibd/tAbWlJ3ogxRQI0v5yn64bYntyxUN51J
9jLC+T/s6XW/nYjToJvjlEOGZYg/FeOZEHqJtud4qAz7Sdn8gXj27wMvQ3RRXALSkZptzvpaITYS
zM85qG5mHMGnKWP6tfA1nNOG1+6UaLh024uDIUxHWODWNUYilPK68qSmehqpgd5CC3m4L3vwwPLq
wMLR6Jz8pB0TMAIywno4DmY5ZUEODsyHEuX8z1mjvfT2ue6Fc4VS2J2IX6iN5SWkIN7tJv9+o5ed
OkDjAIxgxJ60oLs0w+YgsUq6Q4sCJI9kRSANjAG7sXiCOKqNNrzrMFLPDUPsU+GlHIdARsprEoak
Zn3+U5UeZncgUaTccsWzcEd6XGdwYcQnSwsn29G0/0M3dFvNqmp3P+iXYlaEY2agNqnG6H3btIr3
OM4PIXpxeiPvUX/X66ysfxMlkIHfZCrGIh7L3LeCFM66hLXxG2ejgKSZ/76TNs02zqzZdiXkUGbP
b/8tcxW0OfEKlIg2ih9Qdo2cio61taJpAIXp//S2zWup/DeGDM1XMO7gnt7kJxu1M0ST1Ss3WceL
idTnK48X4KiqP/YL1STD/UG3tnn0c8JfmkYdqVhGew8AZ6swTeqnWpq5kGzUFm0C4MZ6WoLye5yJ
JnWn0U0SucGiht8viNsUUwTAVoYHQx62Hx1cfL6EBbg/vZ6Y1o7TBZ/xIp6fxZ4+41PHFvSYjMAf
HdTGZRNdeMAIGVCck245BFaJJxxgrgEddAxj8gB5RCsEJTrZcT9NqtHRqNB3VYAhStyzSxDfJwU/
3jZabjLPz0EpHUjG6lCZbbFJUlkWfKPpwGl/cn/LRWXj/t2Hi4Kzqz6JweRhwI0d7HwH36aIQpCP
tGpnpAXJ5tr5S5+YpbF9QTnUmXbNDHORlvVGHcwlNgzLyev6xgQWOsjI0HWpdJ/CdnSPz/ZNgADU
0pFNmB/8xtd29kCC4QLsEthGV1mhvP5CYL6Yt9unhJe6UaEIq6zfuRlwveaTLNHXHoCsmUidJWhT
iidCWt0IL8LUbfTSlMwDNYJK8uKWlVZIDmGlwkLoOhQYsFT7Q3xCw+Kg53LWTfXn1WxWwX+bclTO
u8VdxV/ws6GsAukDD4I0QKoXrzgipsXGD0btCBeBiiICSQCQpTFaSwBPn5KUC/Z8ATMtE4Y/3B6E
R9SZBj00QFAIPLWpue1BTrL2tHMV/vXzp+mNOr1/f5HObE/VoOP/3we8ECwFYNvdgsLUk+du9bgz
XPzhvQJyEKsnro+ZUEnwpUGBrO6ZFNi5JGFKVf0N+FFmniyZfCghDNNvDD7eDFlxTa58XxfdCplN
EUzkt2+rRKssK5dGyxJfXvMTAf0AJWSZ+jkKXdgqYuGGnvWyUrxb3vu7JsNjdsWV4nSEiEnkyncf
kBHtcNl5aot6orn5nEc7cz4fZn64hhTarcMj84eOgAGKdAOujDAunSQHhRQG7+8F9HIwlPWVhX7W
KMJ2pCRG9opI9KI737V1vHkqyeIYLOnt6mWc0Sb6AfbtU3v1p2ecpXV7P144MqCnY/9zvHLaCSoA
gyfjcMYGC76jvPeSXf8Tm/RrMQRM1nb/2pgrcihXAHHakvDI1qA2MBhZcPiG3rNGlAY/ljS5foAt
pOhoS3FCDEN7cQLKIlZ9Q+yPz/xQbjjRyz7q0vdq9Sj7c7LuDJYFuBtRh98buwJ+wGnUIovazRXo
gNgKRR1eSFUV3BXK+pQzB6jZ+NwctizUXdiI3Z1rB054T+bpSuUzjaU3yyWlrU/lg9ZPmp7ABGIB
U1VSIVybUx3WdAZGLfaXFQ01oS8DIIagj3saiis20qe4tXN0mgsXedNK2bGfu5tPvvhM+oadhDjo
/QSwb1w5kkP6iNjhcgL6wYaaSId4M0Vo/JBtPGposmwfd6+eXNdNnbAvhCuXEwEwQyiohVUG0RX0
rBYqd2dfFtc1LVNPqMWOCygD+DbJCVjLvp8kt/bzhCJFxikuKmalEi85LpLYuKF4+p9oKSuCWpdS
OpvDr4Mnx/RxXKBtI/VOtLnIfdpUqmjuM1oj2cUksBNSuaAPiSo+2hR5bRZEbXuJDBaqjjEQvwL0
/Y+fKQkxdJHmZ4Pc/ZWsgO3HwUUyJGIOaIg8SolDRAgNKUfezNnshaMpYJERh/IWAZOIezlh/3RO
h0BKfti0XkDaMuR2HK4Xgzm9nkY5aqPFMjsqupkCNFz8NbMq31TglVlVbjAlVxJ3TSliJXctQ9Lw
0NBQQrTOeVQAm7imnK7BudowSibJEF6cpBWDgr+Hb0a7w/FD9W2uFkFK0reP22nwRWt8frDRGon5
8jvAs0yDw7WC/B6a0NNTNfe8pp5SgJIdHj/7Kh0ZBS93aTTSF319aHeji6bBsxmyUatDe6UY175R
WXIAmUJyXSjzx5jH7++IaylNmrtajao1eSUmAQ0SCxQq+f+G1Zx/ZCa8iFKzDsz7c8+mM5gtV5Z/
u1HCNOo4DeXwwmWo6f5fBoaIxAIULcKEy8/XASejTg1jbM/ZvKiTwrKmGQUsZXrA2JAr0wtlQjG3
jabUYVFGek/KLpcR998J0w1So6DcA007jIcggEm3qPyKTUvnAJhJvECfeWQptYxNOTgwxhhztlP3
56HWFIaBcmsrgpZhA7QSax53dld/s2uSiRdg98+CZJJfSNhqgtUVZoO/rLX3gbkKIHI6KeksOzRh
a/ci7DEYLNw+NMIxasWEhVv/dEV3vFrlxOdptmkKbEbF7oEJ2imB/Unq8LUB6w7gVWe2wktMslF7
DivdRhqqVw06FxQ8a8Bj1iIKjpfdCcMFOvKurYuajtt+8sbOuwvYng3JGe2ND6kZYS1VwW3ZGZgc
WQBlBa5qvSpryVJ0ZvknytixWsR16w0N/hSYIDV3x2AgQz+KH7Om8M/H/5wQm+OLaJs/M6Mp0YYj
eYjOyGD+z6jEncQf9y4AAiC2XiqeQdGQ9IYh/3862aAjnQlnjGMLkHy3fWNBnC/O0QBuA5qb5p2A
mYr7rngyDIoZTMSV+MaCSdotW9JROY3iE/2UOWkH5OV6OcRJFiSaLaQeqkVZWSSs7CZfoLUL2+SX
e9nuWOsjySS/ooAa1YhHfAwPxE4gb6s7qVzuZoiXDJNLUqnKsBV8oi3iv4Wu5WtRCMeBOJY0XIkv
gbM+jQaf2coTkeCG3IbJAWD1yJtI+CWkY8GWDTzW1V+Pqxd71yRsTz0wtsYPF9wskKvHv0cV6siZ
Z0OFqDmFPkGX8r4CcR4/pLNT3u+nQhqHV6aSmKLAoDFVP+sXy6jSZv6U7REQ7dAryfQM3vJxwWQt
wBHz7p+UZiS2LUHPqUn8p8ozO6Wf6NwZw0xejd4XRjIwdrRpDuqpnW8HJGig18v5xjNZk1Pae03o
+HJf7IujnEK5RGWO1MwW5roY5VhPAdF421O0Ctwtm+Ffbf004nagyvTxuV3TgLs0sMFdxpJaSS9T
9t1ecR2JIRRvMD6sC0x0TLYMkfoFSUH5o2B1pP+bpORbFW1R6WDM6ZY3kV06jcIcge18QbEeXgA0
TrlKfXAUiWwGekYY0FkYW8aq3hi7tya9gHsUUKlpoD9hJkjpDVqIx+8pSDWQ1/kUu+NAeWJY9B/V
rk2IT9RmrBK7oMFjIi+NnZODXtKoQUlHi5E4HSBFhp7FLbSwsYXIt0HSeAAwJXU+44qgvjEsuNm9
mxQHJ6fL/s/a6UPK0Ai0roUAl0EHVbFijoiCHDsg07p+UC8qer2Ih5r2cEMGmQ1VLoH4N9jkWwFq
KxRNUp6ozk6zS1YnOMCMGZOPtRzQ0GLy9P/wPaJc5sTsBWyAWmGzQ0I5FOHZ1Az5maIHnNM1Ra/K
wRIH878n4+lNqjEH7yQi7egpiILdvXgOqlLzNmwOpo7gCoy17swWRrY3v65YvSw+PKPGwMWTmUvt
5OCxDZb96BtTTSmqtFctdG8IHlYpUTOnJvvBTQ1n1RFJTY+QtQh62wsSjCytAFcDXy2tdDKoqULi
449AcrkNv3RD/g9ehlG0RgaLjqVKBWpvtgQt7U4J/LyX91diapbcikXD9zYTSXDiOH2ViwswvQ7g
JXZADEowHUH1GO2qtjR60q8cr9G6IXF5R99VZ8I/vQI/ClnLJwsgoHbB95IED7GNsGN39SCdHlMJ
w/pBCZ/JhNuYaNbnZwJpOMdPlUDjri2GGMxfglKeR2z9qG1Zq54YIf5rzyxUTMqYHCSst7Q750/2
V6tjH3Z0g5WSKR2A74sDJpcit1lbIXfUYSmpdgnKeaoCNZGixU1bZFg6OBLrvbZqJn9xcXt6e4LZ
MsfFFnpbS+xreUNx9uHk7XYJt7aFKUxU8cKsmkoQqfm2DKrPYUn75cdsTebsDWI2f0ooqbGtvIN0
m2aXiwmWx9fNdOS+fMhuv8STJ4HHXKJ2gTFIeU6Gjq7tsXrJ+3TqTkVzYx9qX0QtOzJ4ZpTIpTON
NbXCsLRahCVDvaa0IRUjv3CQvP3oFwx90Lh0UYOzahFF91GLmMp+n7DRgMZUYLcCF5XY8V3blV8y
VyZKSAJLtUNiXc6Qm0+W/HBbWRwwV0mYhRqFpOx5y9B8gmqU5UNr0+HGhxdPSdhTG++MaylNEcr9
d7HivF3C4xry+0C4Md2WdEYBgA0xOl9RkhHzDTMNeQ7W7ebSLxcByQD0KoZav6qwZufPeonOOTAz
R4d/DOKG6djuOZPkZII1kVtWMr2EIDqWvwCoO5xW3Xkrasl0Qw9t/ndsEVY586XHygAUYhZcGwOB
KKhpJk7y4pJiAjejKE6BfOWhAmNg0Xjnpq7hbCx+cOM/oXIRSueONkJVggEaJvqxik9vDyWwpvj8
0Kx44B+LaprBFpuetRrPrODTEeKr4cDl4ED+Ww1UcLRhRh0kJoBawuabRaBaKBJgNEkYjoNJLm5b
/4kXOSCAIMxCvgA1oJIdhjFPPxSUgkpfBRXMiq1OWNxnBtDE8eI6SygweDE9RiqPPcGyEW+LFv2d
vCbeJVG3nS+vv2pfWZvQgQCcU7XHtv/HJRWzm2ZZ+7OPrV84wAbRIXYYLio3Tih+WLvrcviJGEsT
pcAbsc8ri0E=
`protect end_protected
