`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EGHLcWi3oQtKBVeyS/bZCRr3OYfPcrdtC0KHQ2AsZmjWoi9CdCNNY3cE15kSIumg4ALV16bOWKWr
7XGsS04MvQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fYcCDngAeK/JOFXbMkXqqFwPr7qQUYY0MWIJ22ywbQDW35Nzr+5II2J8GzSlalC1CiUx/o3uJNTJ
jpI7LLWoHbofY3sNggOskQFqS/CzjzvHRwXi348NxbTFu+p+QZDdnGcnxwJc6/GW7ptaTf31+Ya4
TcZkO200LaZWlQ3g6FA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kND4OAADRploGtSlemwskZdynrLC4ZZdHi617phpJDe4yIPOwCttQ/+fx65oAOiiPuh6MbOIm6MI
7owhyW+ufSZ9kHOrT2D8NEvYPRuv9olz8T/K6cTJILue5I0MiS/BQIk0S3dUyEwpQ+W8pnEU5hgi
8qPM8wO8rGfcoBOHTI7J1lMDsILj7n/hUophAyrZriEWPbUQGD/ZnP3YFs0SQkS9ggg/sJ8bug9X
SiGxi7z/9g6Gn4deuVBXUZOhdw3IbuDKMYTViXd232BECJFfF6Sttsufr79UuKP24o0RE+G/mC4E
9nxBnsIqjl3D/oJYHlLA+3xriBbML1I8/Uphfw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GD+GRv0V0tiaJnIdZQVmniXxhvkm6lqrIFKK6IdOc4JZ64Gl5XOkP4Aw3lIAKC276DfiPCc6xZxt
KVgVPgxZJfDy0HseTdG1yiZ64EqCGIHFiZ9e65faV7S0+fq/CfOEg1ZU+VVbVQEpo/cvk3Ld5WmJ
sO+kF2K4tL07d5Fz6D0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fpoD7fjN44iYsJ3yWP7aXkKvCMFJXWCMk2ErTGcPw2S1Ua4I5TKv+hie7SO/J9KtvOkegmr94d6J
gSf0D9UMXcxp1vIKBa1ukuJSmLQxcqdmhPnEfIaeG5tkInCRoZiWoJJ2+R+1zg2bmEf7iZYibZ1K
q/DAXPj2N3x7a0lH6sVn4ygag+o7+q/jH0Zcyp5OvWQi9LEKljgBPe+hct999CmbGq62TOUPv6CE
uLOeJngp23e2DsFlHwgbBHs4sOm4vvMKve48jaLG02+Hc4463Dhr8odshY070zH1Cqu7jIBHKAHn
jiove1Mge0hMje9BeXLCD5v2AdhIRMiC6kkzug==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12256)
`protect data_block
hZVagWPVbOOe+8Z/Yn3o8J0KP3+08R/tgUIlDEEijqzwW7lB4YCVrpJ0LSEwIn5/5fiATt9wbnwz
LIUj3sHIXd0LV0sLZl0aTNEXp689kIheLlYF752ZGFwuL1qFjS482aS0lZfWJhAZydPhFED2s6S/
Hf195uBRRs3Zz1nRp3NSgYweW0dkR64anXfNC7PRIMN95xm75k3uGY52YQYThgWnzZr/mw2odgbi
uNMY2+geRkuUesZB5Cs2sC6s/48mHzdnSwbBbXwo1076N6CfA+LCMBYXDmgfTqhP8He5NVXr0Oz6
AO2AcAwHerb6wbFrL9e2PLR/NmLOW4BxMoAHR5ti0FOrG/yDENQKEQc/lQkt0vVYgdIHelgcwNHc
CMfZpm5yiedjia2HkjLYvVI73YwzBpF92ZQ/HS1yXqWCBHMxzfVmaRuw1jD+eMKRlzzlNYe2nxEG
mMgwtKhc5F2tj4ob1TE+PmKtLNr2wf6Lezaah0wgSpNxFtx0Ss+Pyq0+uuspAJvku18iRFchEggn
di5uv1tUV4neW8Yj1+QYvSKVvkQZKdjRYuPL3uw+x28vfJgBbQHPcy2K/LQyTd/KT7V6J6JCr3YS
neszSQ7MGbS6Rx01MfEbbTjMbFEurZ1tMlb5KCPPhzcDXg+60S2AQmtTTaahp6j2ykUFUUWwCUYj
ocQKhBIGcBCI5kxeNj1kG46k/+kcIN9HpUjaUAIezxSzxJYhrInZ1dXzFQVKl9pSoxB7RcbRgdP4
1hRgqcZAKWvCEQNU+VLeAtR3yLS8nZ7MTLTf6b1k4P3IM8Ua3gfbFW6ZsBumTuJFaBC3tBTyuBdD
AEg3uJptfTP6Kv28fYTSs9qZcOUoHQh1zyXMbcCyfT90hoc0KaHdZdhCkoitdn6cYuADn2CYKxHn
RXq5c9dr8Fr04vCISpeXjlyk165Hsg2N1+9ohEeZyHVzr7/tjfAiiEwwtaOnWPorxN/UT/9WWXh4
ZuJcqDQzX2mohHO9uPcCgPDK2jqTNdVkD986vICqs5KuR5xX5Y/bG9OGlBoSEK2YufXaS/Vumxly
SPRnF12aI1BZLsmS4SIrLWSdSkzo+6XF3H8sXJJQhL4EWHQTNg+fWcXe3BSnssh+/tF5pmc9vIOF
GITpBiH/cewGEWZ23XnfFFgrJ5LWmHxuIdu21eIBLkKSbeaF/CmPw2RivYSrrM6P914wdo1weZLu
GcvWVpfNrJ+jWNezhE49i9Szi+MoHV9jGMp8iLtbRpTBRYq3/S2Us/rqIwP8O1d7A4EHDyYVI2Yd
157xIm5gLXV3CEdcuS20+31XbB2ELdcdA1EjPQGPl10Pbqbz9+aT+RgiK07n5A5s8yFMf68YWatK
APaeWiVlg/AQjORZeWsB6nzBYNMcXadLzhBpbcI9drhQdOsHGXTyl4FZ0hguRnbrW4GAZq7GROiv
dYhZaLpzQt2toX7WHjgRaUkTxMqfQz2goWXCDf8rSEM8p5RERIUmqGi5Pe3XINuJN2af+wSHZRq3
dKnWmZQKBPWbt2yOXhkJ6BzuBtBDF5IkSnRAUjtrCsWZWf+T5uNhPengEXjhJ01jFSCf/KS3DogW
vAneFx/i8mnG/9Fw+XAjMD9YmhTMBI0NfVKy9IBPgNqYk+ENaEnQjbWKRvlAfXWd/whOE8WeqbM6
7tNMVBU7lHEBxlA/CUaJqY30mr7NinmOb5rJezdOJ9bpyFoi3G7JpaO/r1Otcy1U1SlfwMTB3nnF
qLN2iIphoK76vIl4KEDA0ATLDqElZNcUr+PHXWMFUQxMUkaQ3UKwhnG7fo1s6WvKbzDEWmx/JpqP
3IKjVpL/yaYJIAUBXe7FliJvMc+dyOL5f0J/6C+5pIWdkezbcWUByid3eloa2PCZCZelS+sn2n9n
AVQXpljSPGx/Asgk5vlYbY3TYzXGGVrVYAPdhSXjoEPGAQElAAPQOpp3e9t04/LI6OQytKIsaiSV
SgqGkF47OfANylEQc+aO8pVOJi4Go5ZvYYMDKRXJ/NOyCw4lRFKMX3sdbGNBceaSqzbAry0uisTm
vrfIb+sYq2wpWA11R/vCBykH+oiTpdDLCd5KUqf5SGJ6sQcaFmITVWlP3xpQC5gucljbFk+arWZW
SWTo5zXyYdp+Q/8VupaFNuy1us2T9X3gKtwSEmZxRvNIMoiUhCOpc6l82hmSdUfxPOPQmaaFq/xi
0bgh2fikrSMZlBEudoFIjwtkGM5xhBCrxkJsEFkgB8v9rGA/KqhuVSSbB7IMaqmM9dmEq1AXOiXh
z4evB9VPUG4egOuAZo4ecWmDXZ3Bq4z1AcolK478CljP4ML5cKZ3FG/pTvfIsZEL2bTJVyQ8CQ5x
IcS8MD1KSz6484nukq6bFbUy/lTdjvJyZGI9nO+tqIY6P2WFujDPmTqZ9DnYtW9VxjmrflJqwN+K
BPV/op8MYwf2BvYZyniScWRq7mJLU0Zvvl5ztHxXSJrAFbjf6HV0sovbJOSlt49AIbOnRsdpSYem
AhczRtvX5AgPRdC9I1gWiG5fNFKNU5tBv0yjwYh+grFWh08viAZrXZhAcAxKBe/9WL6DhsgR5wSQ
dbqRvYGCY9PEuIOal/1fywqRkQzJhtEcYPi0+8JKPlZqiii9SJ/SExU2j8YprfcfAu9EWcgzvfoK
4dUs3FLlrlyPa4RDrkI0OgxwcYnvqrQKcXafveflL9cMm0rKIOgQqIFQp9psDDdFMo0W3nR8WxHI
3AmZoVbpOT9IYVnyUJJ/KhBkQk1IKEz20fq8y33vqhw6r2syenLesZwFW/w1pLFxys3Euwpz3vpk
iggen5cD4JimA31jwKC3FWK/UyaZBIn3WgBW0JbS8tw9jykAmXm2UEYSP5mTXWFgY5iK1GubiorO
LPH/6JzSLggN/u9P9NaWZsHaXSkzbp3LjM6pfTBwECg6rcet+MbOnu0Q4VAmqvo2GEbUV1Q3/x4h
3mQFikjFtujxhm/fxk9Bv31IAMQOtK7jd3Bg3n39KP96HDx1K2L/RUggf+HFXokAiJKzBAa9rLme
Iej4bZpr684Jydpki2pQwuLLGNBwz97Dtu1Bo+OZbq6Aili521eS3C7q7Idh6uD/4bxX/A9VeJH0
25OioR3cdL9i7hlTCo/PQ/XdvGZnNvrPBSQ9qAQLkiHSlt3lR8GyF4af2EF8vhQJZQUiS0L3HJLI
CksssfFCOeuDfopnVAY/JZlwrxoE/1xFYSWau75kkF4m+GRvU6DdWo47ptzK5wzAJ6PpKEs2gu0I
sFy7TNF0K3QDO9CByPFyMWierDy88RCDHbwvDF3hywhwSq5KEZgLBjp5jfMIbEOyBBuwq48zgi10
PfnRQotz4r0kw7JiqQtKiE5ywObB07L1K+nPuBNK615i8EdsjwvZrdFGJJ2f2o/u3E3qZGPpDGJg
gkPmhWtZs5Vp+ubTzaKS/DKSLsCRuDpRHy2oIr7I4iOWb7RY66FVVhhFcCwOaAx4WJx0YLwn/CiR
v2EQIvbpt3S0LoIaYtIHYCkGwAxEzIOiHfGK6uDk+747X3VORZYI15H5jLPK13qP6wMjvJC18eda
m+i24vyhOdPDaan3+rQWm7reO1tuaP6u+vHe4ie4lHVihiSwCEEbBrBWOQV7UGFppN9EdodJg28/
u3CiC8kRIbjYCtibs+JGeZPL9Icnpj9CDcDVJyAmFxoB/+ZkeBb9e6xfNxC0agJo8jXiUB2DChmR
HN59yI3OMtKW6D/PyPBHb4JED1xrKq7JQkuTH+THRN4HljScoSjo6xElDS67tTzAANA8Lxq5eRxH
vPniJm5wcRg5wJm8UoCuzh1Opc/2Kido/ilPWigM0pzl6YG4CISZSseO8IxCYBhj+8GbejRS4BCo
gpsRp4HPDlIuak2WbLez96vG44U+i+wA7h6GC5Uv09jXL2a0CN9tWtNntznGHBpPSt/sOvrx/Cgn
SDnbtMSdEzE9Hj+9ULstvkZgEUk3CsIBrLohh2Rpz+a8bJs3KOjlJnU+rJ827xAZh5uiT3A1xhQD
WMLaF+7fxVBlA7i99nASR068o4vaQ9Ynky2qsJL7ZL4gR8hTqhcOv96TnECz46/ex6TCtmDIsBnk
dF6r9SOEtLFUrfZPTmLmMbSnbrSH6JNXH1ApTWS/M7sc6RYwSo9K+LbZK3OBsj+wdMoHxP67wR4s
o3KD1ilhHlKK/735G8H6kWinaX7iXnkVn48Wt/lJE7dtTN5ClPXmt4qNXGvr25e7JXbXCiYP0RY4
dJGammpM+F2Oz3w7D6UTXxZQm3aCL1hoC6XbVTvGserb1TNmn6Jdglc3Qt9TuHw6+MYUSwGVPc0R
7542XVwvbPt2AXpuZ/fC7bqakG3Ax7Wju+exeTaSCzRlab32zvbnF8jDtmezZ1udKmzum08S2JX5
bzMZDI6yrzLIOfkOpgUJ2eDx0WdDRPbcfr5k/F/nbUgj+MhJJF68R1NNGMe1JrFqsmPcH9gRRq62
nVBAvimHOm50VikmVNKPCgz1EaSpthqUdwfZb0w2ElRGy57RCzKaodXhmtu+cAFD64XKhlvNmKti
tIQhcyxlOpMUSDO2z2sseOdOPfEUp/aGlw57DXt9sGFMcHR0Vdt/5GhzrGETe2MbXHdwwFoiQkys
go3929u81rB6Ef941GKmP5ZYCO+YNNqRZttCMvM71aqihlD90I7KiCC4KXBCpb2lEa1geDutEFVM
YPzcbs8gK731DskiAaJAgSRNnPBp0izG0Fj+EEk5pgzRm+9RVs/4DFpUlm4PQeGZvi1tyESqVxWQ
jQ1XRLtrtFmRHrHs17nDkmB/jD3Aglkut5xdThw9Ew0fOQljdoWmTXBGfOMXOyzmD/8CWrxoWb3M
9YRh+YFhps00vqAbU2hg0qumqYV0RXHIzqZwQlU+bf5zZkq2eXyHobMifUDB6BNAi5Yfu6qXUFUM
24a4WMSzKLa/pq6Z95cCr2K6sZmfy34rAIZQpB7D37k9B+j1IoOX0qTX7GjRvVysJudM8O5/blIV
nyS4d+f6pEkdsfKmtwTuu4+UaXP20DSsWGBNoLLSKWyUv9Q/5AiNjSN/XBzKZ3oMfMDvRMQGxJAi
eV7dDF339Mg1QX8ImM1n2gl1qDTR4nD4m1Txtntc/KIkJ1l8w2PnNn2moR5jeHY4tlrDDVMaacwa
uElqqjsPLAUM56n8YWfiIMpBqbiOAJAGug9OoCSah1V4At9WLJlXG3+BLKR4QVjao9udhj5i+aA9
obnduAN16QEsLzOPzcOpY3RBcfgxcalfmnKHy3d6pN0Z9yCmd6LJpz0fFTz3dDfxPHt1h/pqtKvc
zR/iGMKzFNouciYgLPPS49bgrvpqgMSj9oOlrH9vQqa7XIcGtSmn3OS0VU73Fwf+AevWWmD32MFi
/S57GgmiAQ4gsgrdLQzHAUYRav78fpJBeeJ/PQZFMSEV8Y/Hugdsg0jnMGaw6cPmtrvw8Sk63C0n
0VqO3Pz4l0NWtGpia8ZpRYbcCO0oSEdeJS0IrOYUueG/sXHwqObDtlrSUHqQnAB/uru3GuhILyAf
TCp90WTsWNDdmdV/+Lz44AYSI5eHM2G98RqXcD/qso5CiMIMn/xGF26DD0DxXm2jQMDmniNE7THT
qI+n6R7jEwh/VXWi57TwmLTKCGgdcf3PvDf4dgbX7JFULcXkd432rgiJ6zVg5MOPUWLbraud9I8w
zji58PiNgRMQBDfQfKnljRqb3o4ONQvHwL2pt6O8KZUg8lSjUlSpbdcuQsxznqnlzHBuA8BJHOXS
yi9/DO1LaAYgbhvtJn/eP0/faXcr5lAaKmPyZ85nn9cqcoCn+2IJ9THKJT+fq0HrntPO4+4Ogjt2
3HVdxAw601gPnooMgGd69YYe14j3WuzirlgCbCoYqkipfCWWwRj7LGv2rO6x2a5pnZRpU2EImJ7u
VHvNmk5Xb/2/dWDZ047h1KHg2sYLOUUPADLNzmBZUVgGi2ILad/rsj5hF3w5TOSY/T2Te1Mcphbf
/OesOzw1rqa/cmEdl1hO9As193M6TcFM3JvP3OwANeO1mKqnzzQNwNCUA1gj8PO/ohqgrmQ2QpBw
Mm1fzkrss3HNPHYKwoxI9LF3GQBf1eeHXznpq7oDjBttO7W8pOANh5NmOQp9y46lAbNU0TrormA8
s0kTRkoheu01nHno7JejgpfSrtS9SmY2evl7jQcb9kuUsuVG+Ovx7vVI7+1NGEzOS1ffTXa4p7T+
ktAR6rSCrHYvDmjPFYucrMwDyOuMZsv7ik04JPFavvf3M/UtEh/BPKJ+BiUOqKAgqeUIe4N54Ebp
iCEvrgoS3l8ur4XTwYy63r7kcGBkCvyPOKSSQF9s9Pc2CZD03zN/YcpFyZ05hqosGDNg/WI9xPRP
3kyr8YT9VIe/8w+Ni4aENQV9UYXdDnc9ZJCkoDGhQL/PQ4za7636WUO4t22aBqCcSLZRiSBQ4k71
qMk/Mpq/S6SYpnS855gc0tISqmloZT712tCYyoYvTpUBzbleOr/7CSR2hds7nniTRQAgB8xaHLxE
+/A6TCfn5SaUxGECosFhxGY3C1pzGarzvKvEgARtaqyKolhxzIg6A1Z1tv3R+RbC1a0pzBfuAi7j
DBlDyckH+Qj6ahdsUErwVFMUf5clkgUxHuu4kFcfTT1VPyF/BvS3G2lKZElPQyUugOKmBx2gMPTF
awQvtGGb6Bw3B6B7F2GDaa1nL/g2SN+a6qxXIqeOE4O/nbxNxRmmDUs27E0lNggGNMZhw0Aj39en
OT1f31yLZqsMh+Kf2TH6SEuLue3qf0g3vZ5B93BIED/kBdQF8Pq20gaD1CztZe3SflXd1d3X4+04
wgPwIjAiNgNbUUOGVRWicpN87AAlIclaQCU0lUby4h0X7/rD3s62kTisF2WVLZY73b0zQDucyw0q
smRodUnGDVsklC1d8h77Gp4YM3t+xXVEZytqbtSKJLhRBzl9lIirB05iowT89RrT7S4YA4gPsu9j
82kTyZRIp4SLjR8h/pMKXD+ozy9pB54b5MnWoEU7JNZphlHrfnPFYGRUV0XcMUux0XHnbUM4jwFk
OgMxdxc3gRKx4BQnalj4mskZqgserBht+PEi7rBxMt+kGfX6f+oDKUxNyrmIlkAHrQBz0LtNfxiu
WPlq4nN+9e4wVu04H0l/duXQYV1K7eQlmmFunM7JCf+lN0z0SOW8+EKlAgnGkvO0EShzQX9iInKB
6k7gMsoNma1aEe7VrfT2xYvj/nHSQzYVRA5aMunbM9hxubRSf8aZjKiOpcPFNXv6fkBUj3q0cJAo
KRsYHWP+JBea+LBjbgtFqmnnXPhP8OS95XhT7vJHEycdVsdBBwlUVLnaRAwx8V6EHxnh8/ZEQSJ4
XiH1ScjDyjgFvWSgSZxcpwKY92Yg6HMGulCuIQC06U7cL+aJtQgF/M7/gqMD1w2UHpZEHnuah1o2
zAXKN9AqRzJ3pvqdL6vb0BK/ni4xFBjYz0qvTIf5S8labsMqxo2+RJFFEqTkPqlRNXdlYtUN5S1r
8PEF4F8kJ07FRlnWBgDwmQK4YPqpBcWqmEHvO9Z5HS+EIuGhuzygGp9E85BWh/+WHFWJT4ffrD8b
hFA6KgIld8rEQcUpVD9AwIx+WmApUXIEEvWSvkKNC784ELoyqtSm57z0WYVeLjlBBL44/45acUPO
w4TfanvyzvgQB7Rsv0q7siiGxbNvXNNViVFjQd4laLj6ZKm8K8o04io6cXz4C4ThPy8/ULOtVTi0
3qYqnpn177y3bYAxkrGeEgeevwF+4hJ+8CuAfjYtS5Ftvru9V9X5qzQaCnt87JKpn1FFAkpjQ6+W
H1/JEsNEeN46OBTa30USMkq9wHpBAKICkKar0kkANQxmQxWsjToIDXbxPgYZmmhFE5MjxMrss6SL
/rN+U8BKD3C3r+4joQ8cqhWNzpZpm6fSjmPT1JnYMOTvgpZkN7p/HHJ7VfE0rZLQbw56glfnNQ7j
nHmS6Hja5HuxURh9WNlwg2o6EsqkVwpAXmWwLYXDmpm44r2O4/+3kSaxh/CxyjTD+pzRtFeOXMhc
/A1b1Pklq5jfdvzAZYYa/RnhH/9IyeMPtwqLRw+T7+6IrYIR2PpHiEJDDfgq6LD9kuj3hSnRs18q
W2lnU34hgj2gHj4461hj2koHdM5c/7XzL/nSbWg1KTeBQqzhrsGhIwygW8tQkiCdg59ejUGWA3q5
0SkMILLq0edt8A2hRvUt2eNQbbGwyoqEneLjzIUD1ofvRyb5Aserp3lcD7hmENk2f8Q1eduKTI63
B6wWcuesU+p2ASwF1dc9HNUbSfPUJFCyWYgdy1zasvI6JJdn2v9SRnpVsXJIGKQPpIaKscTj6XHI
l+diWLc974I+VaXllWMxB1mu4LBhTKP5ZQKe2TX69EJrMA65siUgO3y4RVwAD/0L4bAckefz8mUF
5qy7yHadtPj6c4A8c6gzOoePRmdv37/TlcYhxlulBqRgAHpZjERsyhrfVg9S7cJ5fQGVGFaXeaAs
9lxTP4d3hD17H7zDWk5VRkhFU1ABBtnyeydvysy2vZtHs51r/vUySvjE4EkF0R72I2GGLT2oYzCq
vnKMgX0McRg2vv6J3ACKkZPH4ErBULpGg1AYhW555nR8w9SnRTALgEGM8QNwb88zZjQCsQWOApql
xhTW9Rng5VW9Nws9jjJypdDaHZojxEPwoMjNJpcYi0HYKOC0LoRnSFyFps+yMW7yQ2I5p22JidNp
2JNmTMvo0Z5YBVUnT2VLaxx8ueWtwAAXB3Gb3ONNeb0s8tLC+FTmCDW3fMpGar7A1XR3c2jObSnf
vhBpB6XzVe1cohE0cUnLP7JDcY+ITp0x0qVyA/nQW2rUd8NkjhBWX83AfjuxJZQaPfc5Ps3zaoha
WzSCGsxxkB6lulm4iCuCgyKre0i7JRLiLGraI9oHD7zSn+Wfih9piS9cZf51Of4QoktloiLhfziM
hjw4MsjOIEGlLnTCC0WdWFGC8VoiH7Txn5nuDKJ2HP/O87PoLuaxSe+REc8bX6kcF/4dY7JP5Elo
u2xjwkmO6be1aZekWnFC8mTSGDXfri3Kl6FAy/tsrrgV4s/HOH47e1jc/TzQqO/+UXFS/Y1F4hmR
8+wUnoj4Ivnw0mScc6DjnMQ3PvjV/QECe92I3TAV93bm1u557ZVJBfI8CVJVzhp4wzAzsAsZY0jr
oT+lm4F+oNFk3By5y/HGesrBtQqm+8n5Kl460TgRSDe5TbsAJZ5jd8KCu6OUTd+BC+H7+dyzs6A6
nXUQybGFByf0qCx0t6tIPa/fJpykgP1JLZ6AX5ZU8qXk+LVAdzScb+jrJ8MV/I5PCPpPyH1EOiDs
o+45JMcdTDCEGJqFxcB/HYORkz2WM++5bJ8zkV91WjEx6RbN9/5yqKM8hBEc5Mq1jlxdIknrRNJX
PY76wSThUEgq4bo5wjFXCXLEh8N1qJX+lFMfNhonLwfO60/sn8ELWxvOEcVkez/H1rX/Wr4Rw1jz
ggF8shwHkzM+3QyGioR7rieYQy5PBOSBqk2ZErLjaw5HptCioMjGwVp68q+aAH43fEeKOIO3vbvf
YG4wFwrcyYxYmg5VnOhhSes4go0Bm8CsZWv1AV1wJ/A76OCd23At8/dWBG8yPXVDGGxy58W3LebH
d6CJDT+wxG1xhW0J3oqx+hxy55bJNKl8COOK+YgXSEJ1IQcVmmcOamJZ0CuOJkMIaTfOCYl4MYjA
63QZIm3kv6eEF69TFjKcmatGZTaCqGgdeg6QF32m+StM1PpqU7+8BqriA9bF21FH3CJRk6yOMUn0
kwsjIO+7/R5RPzmUhaX9bL1H7EVdVPh9p5/HM02JiFpbjHr7ipbV3+v80RMfh5/JTlhAKX+Nz036
JhW0NvLOd8/Hky1sUVtZujzF4Td2IqU+89hQE4/71rsd8XhDkLSb6QgkXa24IZHIRGpHdOEBm1o4
i3LtRe+vFGfjO3Hsz+gzzJl92fl7fnHH8ola0U3ZmQfhLbhZgKQ4wtPHs7dYAB+TNpDjaKMtPIfE
73BwslTz50Adkc3gZaQz3mU6c2y7+lBpvosLrvKdOVQ/N4IOPHmF32OJ9ZftbWyIayQ7RlJtCV97
pF4npC2kMJ6gJ7S6LyiXRjnGrG6vRCIum+Tul7Ylb6zIiQl6VBdJF3yL5TGpep82JZTRs66xgDHD
w9Wob/sMGPBPlQoAbIzsTgNotU4wCrQP29v5rZl+0IS+1epjl3MI8C69e2h2zhTmKvmeTOdmsDBn
UFY7gDUCX7EZWxes9JGw/G2dH7sf3iw19cOpOhLpuIYE6E+GRM2ka4XE4YRAWv6kx4B2fdKIHWKQ
YdQFXG4yClgScidxYegk8+uEadcb6DKAl9b2ZZ75Vl+LV+pxkfafcydbC1r5ZsWtsHGDxCe5lWs2
3Xvu1/Lvh6aOwMiHep3jlP+u+Lcpl0KTFbUnZzpFGV5aN3d1I1WcCrXjqLidbSQmN3vQe7It+Meg
2zPD/eNJFlJe0LvxR6ARJ82CPpYwVqM7H//yy2etu1KsKsEGE88wfYJGEH8P6kC4b7NVgu++KmHl
7L+TqaMT+wXUo1QKn/gJA/UVOgHTWmAcvQvPWkWG4mvMlMk2I6PLMP8poQ7q7WlPDHv7j6m3CTB5
A24F3pemSpCOK8aKcU7CNyTlB/5VXEMtl0hBZnp1UXYlADdo0XCpmtMF+8fyfkg/snnVJAHVA13e
YJ+besl/2UTh7mG3rexeG/GPdCmjUGWgMrHDQtb/il0p20HMituImIgBk64KnQA0SyQLRITliiXA
L4hgDqJkZL6a8bUnPyCyR7ykn3s0G4T/0barEVonVEcw82hf//hDhbcDmt4031GRcQookqO/zppQ
MhmyOT5s1DBFeeen1i5RKz0E7cWBaKJVfn3gi2zdN85M+HrrllMu42o+Sn2ENIYPwyMP2lL58ImC
s5nctDdhq8Sbti7lsmRcIYxfNmk6RiDFD3U65W5RK0O0DYY3Pm+jpyr70EBgSlRmY1SsxkmE1sgp
g3MREJRwI5NLg2/Uj6PAUSvG+HgZNJzRxutERWCC5SRmlvD4YmRbGQzlMjs/m4Gy4vZc0ZlUGxMc
s7Eop1/wQUJkQUH1c++9ldbmsKLos3YqifpKDYYS3H7d2qTskFj2vmXfNTjARTcubRjBIiBiWUeM
vxkB1u2Vv+lfoMWrVBlKx17QtsU30Nmd/xvQ43lr9Sj5i1w8+yGQu1gLESfYqexwz5Tt8/g2actg
Q1zOcdjBJQF51XTTSsuLxGQqnBMcc5rmcBQ7w1tEoNOGSIZCQbI4BRyIlTKpMrCalS9o61j6Flcz
eCdac+qTGJx0XqtZ89Qo5SLWKADYnO8l6hxyeuCzZu0ENFV9MqPpwC7pUljWZFZGqB5T/fjtHIPe
AKuybL4kSIHXnhvBOP2IqrhabDnes/StAHwMBcyvDmIT9KPhogYMIPvMjtoYXtoVxOd6SfDvtrUR
k2EaqrJpj3ycaWFmHrTfpMSRu+SiGbKlAf4xR1pDM9tLwZc+lWoSueVngViuaMWDbR1Zu3S71JAE
olij5PnCUov0x/0yXCwElBuVlV2Zk1E7gADizxULa4yBm8O3mLIBFfMogvfL0b1q5wcOo2R3QkAB
Y3T9fmG/+3oTMlGL7YlcH58cMJMIFeuI4YRIz/uTiIuD1dRdAso4hywosQ4LznZzHdB5vTKurECQ
9/htVpYFvh6VY/6rk9TDePXliuQwBBDbkeHb9cS0IkiaMr/X7pn8ARg+7rTmAI4+xu+cmqwToMBl
u0rBqisrCsFJezjbo+Ik4zSYcWBrkb+jGOp87kBZPLMxsP5aUiOnFaDA7jfooBVIp2IcEpZayXoL
uR2vVnYqO7etwmHQ49RFkT65/d1YhYxH7AiGJSyWg23hZnnXz3qX/VP2LTeIK9eJTxvRsRTP2EzJ
ryoS/3OIr6Ri0K8w3biqpywzgSEFFIXiMwIGoOdX0d11/08D9Ow0yYSJfILkuKVVemgIJMI+EY3C
gPnn7xV08OyJr2GHqzdVxn7KQg8MwQ+wg3JxODwc7xSpeKFNd9XOk/4Ej63Xaq17sdmUBYP2vpk/
2L44HUm8/PQ9rpV/bVEzvjCUAvS/4cpTndR56tp5X4fqb/4q10LgAaLHMAQ6cgVcvDCOGh5b1QQz
E/DhS4KmKxIczbjDZlTDCl95aCOeqO3t4rIqJw3gTgValYqt56Io6ul1Y3hj/M58yTrh2wlu7fDA
QeSpRQReTylXv6Jy313RbeKkSTLC/6PCRzirNcVVNueWGDA0bAkZRsSuZ8bdTn97ZMPSgcM9zLfE
GUlE1gCL6/3sMVMBth7Jto9SvLmxfQx0FP7kwTAvAUeDwOFiNJsLa5Qzf211vXlILRBKO988GxP5
Gbfo6lcvXJQe0BKBxJbxNM+S74okj8vzT7FsPinWxDMbtCOFiXkXJUupAojH4a0xHlJ06p8JxquB
Mv+c4YPBiiNjrg8/TOucN7Iuhq3+ve//yMQrqW2CaW6ghY2kOjw9/MNkao3jchF8zK87Vx00v1u2
dD4wgbUOtuf/+2t1v9r3akNfIl2qOT9XJ+6hdVGHrZCnzmN4jbLDyrnt5+RIsuMffC1ws//a8EE6
0YM49jBiNoiuoFP5ebbC0db6hnPmra4cjQVCpXTewBgNbYSFYFaGgWwZt12bwF5s5jAlWHix9+Il
TaBXUZMqAD1scxjFISSwFsIgnrslnM9H/9r2KPWyGFBmO6oTPrCTqoEYFrSRSr2FddBpxx5knbdw
D2lUCST8t4hAgCk7MjWD3KAEwGUV4+RsXhy1jTknYAG/FOw9f+3Poio4UHRErT5mtci9wWAvkZ/r
8fpttsykRml1EOUBnpoekKd2YjXvTfqyrq/Z9b8MlzyQyjtVAF1FuJu5G+uBKeSeV+82l5vC1bxl
zjCvxC5WUscjudabLbjBPsYFdk7PicA37fI0pYRkgzVejRybxsC/0BYlvOKuqErAWTpbOl/2QgcP
3Mt9KdSzGnYkBtJWCZSdAl2Pn/SzkHi5EXiccU8tuj3SRDBjpGEYl6u3N1GvMUyslQSleyDDnoZU
iT84eJ2m2+URvgcWdjcEXuQ7wkq8DjH47Tt5fLdc1Qu7t2uPiy5b+5cXmkqqZmzA1VrKQKCnb3uG
SYIoDR+z0Xvi6aw4X9YZ8GcastptmOfLPay6PEeOWzRxAUMxb14ezjM1SXhy1PaOoR2hTsxygLgF
9Y8jnjJvI6nQV/Ox8WP9fG6dKX0fwHlmuVnUcqpgrLcVSWSCeZPHZbEqnKY9tPlRak3AfPiUzlb0
aH/n9ikIhDGeHcg9NI84IfrPvvvBwCk2JwFX/U77MGYRYKB3i8ItCPLISc7h85tyZxxjUuLuiOBF
QgQs5DXIcCz83tiztLgp0iubNL2Ukd0RkwT8wSz7oXaifTRt8xpkqeFrI+sIs6lZoxwIBsQkpOSL
fDss3b5UO1IuYjwO99YIJJEFlfIJbXo9jBxx/aC5ImCKALBp8JgCtvAY3Qn6AVOwXG9UfJSLY6qy
IjrEF9dnvUbJvZE6pJ/cTj/HBX8+ug6kOeCwZJDaVljMz75sMuh6M5fhfCpp0v2Z77kGVZ24Dxn9
PPdJjtm3itV/Ei6UC0qWBBC6LzDNh4Pkjb7YEmHxJNV7IWGwNoTYDpOJai46b/2hAe6b2UXL7gkV
izIY9aI2fAIrbySdsJs1S+gZZ5aP7ltC5U72ateTJiFZA+8eTu4FrVk25uTcx29+rpJZIFvR0eH1
IxJYfcoYgVQY67er1CxKHhsatK2cZdA8lXyCgQqIYgHXtLCVHYunRjPNLMxxugOGQ6lg1XvNy8ub
/eo908qbdYeK3G816kSuOEXtd3AONlD2tM1ClOo6+JvBBoKtN6jDwZ+E9kmTC3r7E/71AAJebAGW
VlH7R/yh+DuzyVccjJ300RsyBoUgi8xUMIgUIkhqJUZOIqz+aJf/zrqXk5k+CrkY0dcGlXuMlEyq
9Pg8Vrjuye6whz4YLiUaMNe19GxQVdGxvzyFv+nQhLjNr4aeCIgc4bWGPQZ1wrwB6rWtMh7er9kz
CNL1d36a29ZmsM+e8Ohm8T+bGDws50LZ4YE/M7tiSh52b0yEHoMecjxROqogD5TR6OjNVg2w+5QK
tfmp+fo28WPoBNXYjwuZZnD7EBONva/J7Hox64clxe9Kflr4fwtBbHCfvqQXweVNYVRpl6cCCMpf
bze6Y96VmiNjKM3NwbZF7U1MEe6z55IFojIXoP4+FaUTuW+vyEP/ftqVgWFKi1O7+EvefS3uCCh9
NrYO1w4NGHX96ZggvTCBR1Bh+oyhjZcFRulUBtZxfAPUrquxEPS8LEmWab6gWgPUth93XLa1ksI5
cyoBac9M+uDTIAp4Dw7A8+ZYNd2P38Vypt2zjAEJzo3bsnjKRNISETb/jcQ3/QCBjxQfLx7Fi+7s
agX4iGMRawD1xr4iUnsqqeM7aiusuGybRxOgwCdPubY/aLBoLTLMOXk6RvkqFWawUpw5YuvFug4k
6CMaY1Db2foj2Xyhgn3+xh2v/Bz6Bn7syMLMC4qFBHEERUEaFHuuw5QPBDNU3nowEh94IAJSoUXb
I66x+N+0hfr7/m07g+R7k01ID7sezg3of1e4EJhU4bn3xAJj1UysC9Q1obSiLRquHGvcD+eSvKwN
/nGjYn3B7/mF4Y6TA51FKzHLf4362G0iQH9e4rya6Bh0LqpzIaie2QtYOn9UZvZtexvrmiakj/83
sEUuYvORUt2IHBps7PJTzmWBuV5MbS3GXhGtV7ZjqCtBxa27qg3qBlbDSo2FACFDiajaKo6zSjLv
PNCVowaBgYbAnDvgPZOPH09WGRYfL8jZYNrg3zW9p+nqxlMSxSeAg8uFY0JYw51CUZZrTjIW73am
M7+ouuAd5ZJ8wJO7PS/wzCITG2kCwcvaQsov5rI9jTNfzKLPGpAicOARz2CkOsuzDhEmefoWyaf7
zOAXd31ifJpCR2ZbvTnZ8Ra0PrrDZr0WuGibHMEfC1+u6Hp8lnMRBs15wquykqBDD/RK7tWCNrjI
WbkbhjSNikj6TgnECiBPhRGzHUO/peNxtqNo6OUZIxv/pcO2yMCvjqhqiBDNTgRCbVw/d7/Ut6Y0
6n0duJqh1jUwXRWUGm6WLywnxy1B7FdeWg5fFR6G+IDK/JXyXM5Q6D/uOXLRQvh19xNRnhKEaWq7
3misuFptsXYareZMz9FD6boVwVEW+HaYUyTKaX/f+y671CXToVXf9kzkbvhZQFG7AVdBvu4DMRd3
tTCl/HapfCIkpY9Rsqgop1zSERtaOEZuSDrHPxlGLmdI8EBLFURgE7/1Vux6fzDG9ZN9B8l5wPlq
d61UYcjWfHe6AeWE9tal+bIUKoGBITjQkTR1GvNd/F3JvkZ4PUp0YFX0NbBs77EzYZTf9Ujp9en0
ywV1gYfSEShxoVEHYLf5SRfLFahkZc7mXuNvwADHNpAUto3P5/471hzXdBDVBF0/aNsnxEH8gXxk
PU7VfAgns118U3nSnEYlp2lVpjQqJdfA4cXu91X2Dj0h5EnWs3kc9Y8TmgYjR+8vetFD2Rd0O+Qt
rh069nPGGOoFGPgAXQQLga4hjCQhUAnw+jsyFyb1G9rembaxFjaaDlUTYy/EgqZYeMHalsh3NEYd
NRP2ey70Fkaos+9MftQKz2uwaLZxB9AhguZzk6wo2sbl/LKz5UvUDme+A1jkuT6CaiYrW09/TIrB
NWzR7cvxZzsPkNVInTMX/xDIbgk8jnTCBiyO5Xf2oSETvx+q0waQeoiCcjOrX/BLg8ulv9iSg9zy
1F7tNC2IgxHQ/CdqOsZUwy5Qz9WyR8HZBm1B2DQXNqI0II/5P1cwASQTW6YSPMEql5JKhcktClOJ
li6Oo46qBvwZzQr17QA+uvOMEcy5mkSJqhdaGcNgFv2RIzJBI9Mt8sqacs4Kl9p5CRRG5CwRrJ6i
p9kJZ5b2A/kOmyTqpTqiUV5UGcPvQ4FcJA/eOF9zxQ9DKqQEOH25p1erhvGMkpAlLZ07sW5Du+Sy
inskM79DdMRI8evYr22rVxVgycOJnwEVcX5OQDRpcgBc38cwCWGXGZZbIE+UpD44r3KnWoXxsP4V
yQd1ziiUzeFFsUQxJytBmjQjxgo26DdP4MgafFwSz2vqjNxb7r0IaC8rLZ0Rm496dc2RSzPWQ0QC
bNiHXLi0jwILzU9tEZMnEuEGErhravOnqrJgSt3cZQecZ5wVIk3AKaMAi0j0OjWbuA3982a9vvUi
ZQWkqLwWw0FpyskfOSLQl00SQcZxdvmtjIQMI2rJyfJWfbqA//9xBwCMccjVyIvjU8tXadtylbIi
hQ==
`protect end_protected
