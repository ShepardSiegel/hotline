`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ut6eNwSNS73oTxEgoRGt7N9JFdYfxSWYmAF0gqo9x+NDfPEZw4M2q/TdykiHRR9xyC301M4DetsW
slTlxDXOCw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DHlw5NxMAYaQNptcVLJkS/Ef464AnPcq44mpu/FIPwGnWv64GVZ68lTN6zJ1gNxI5rrRoAyC5dNT
SuAye1zAK9V+Y8of4uvAj349kO7EBkBRQw6rSDDEhQaxdRn+BHIJmqp+L43TPr1Iptri7nFVNbEb
CVspY18nd38LcE2ih2w=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ViPqio9JLRBhz4R/qB/ldlh1cp9uH55ptbhZD8LOGOZ+xJI5ezF9EZ/Y9i713J4PYIWKxjmWVY8s
fwSJ57bMPvnhcuI2vIIs1kjxfWtl9Z2bEqzFATRhP5HuXWlZuzWcqK9o4zLfeH1KIu/aDAB0ZlIv
YgawTajFMIR1WW7V/WJH9czVgEAJnXJdNA8+Q36YcG32KIZtINK7eBS8ITqWUVmcVP8ssrIDe0PJ
FvN6QXBq4sXAnOASasdpvrY36QIE5TVHakhbqIETLJR/TmE2k6L/utZe9SnPf7Ic1SJCsQsqozI+
ZOq9oWa/xkMOYFn8mDpcbLW9yc0Yfy53lNgLKQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
V5Oo4U2mZRZdVmh4BCW1+HPDM7Lo7/c8t6CdKO238mXYXaEwvGjuwdt2FLN/8NCja1CrVlTR0sx/
Cnq1/kJ1vSKXlEcVU8LoUebHHhjxU1hnC/vZ7oE5mZf10insyqXZIRU9gv0sSp9pdQyQtyc1UR/J
ssnnF92RPeliFXd/2OM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KucqbCj0U+ugMzfkCcSQvbcXUgY5dvaceyopbbW5QNTmbdpDahsnBA/YwEYsubJeG81GwD5EZ0pD
FxlsmcSzuwd5HITqj3VJcf2AhrnJLQvsDEo8PaIjzX43vSrHm/Wmep+X2WVequtie/7xduVJyPcr
tEKmfSptSYMBQvy2cRjbrnmZmKWpOzMnSUOybxZK3Qzz7unAxea4j5//a2cBdkDl60KNyewqewlW
JPZ1Om7Ks10jolxg/ULofM71bXg9vnXDccD2RleiyyQGV7ICF1d+QQfkgGUQGqoNVETze1JH+LED
GIzvJUIBemGtzb6XVleCfNDvfTEq91suMyvZ+w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17184)
`protect data_block
1ppByAutUHD4fGKO6nJvqP47aPbJDnEbfX/zN9GA9NffTbZcndlLdwioGGHrknn8XJjU+RjfaWbB
SgRUZutsPmvoNIxxZabEVBQFDPyJ4LGRnGAIqoc3PfpGFJHfIOJ6xBhVYdZKzqUlo4VAG42caXmL
JSvMYLbiPFe6g1fq2Lmgvnvl7i2XVVDQM1I4T74dJLdj3HIlQKsHJqWWSpsLxvNBwe3+nEklWzAp
awHXJBhwiaXLP1h3MMO4+qdIxCAEfZhfpp3hDj8f0UYCxUS44XC4MWngHUBQUwuCR7dQngQdIHoV
xH0adbBLagOwQtJ+DmWDQCxe/kkhseYoNg7HlkO3QRUfRTlmBnPeCMqNWVk7kNUJULnDK83EYecJ
btdvICQGj3wpZAZGLw6/esmi1lWbB7E3GJ1KjEN3r3NzfFbTOtbuo4FoyRqafJu9Yk7l4eq+uBhd
VMGtQ3LXBU5IgUCXrgMJyM9ql7iakDKruKRfsnvgBumNTwhe5g6G6nmjF/cqpdGaq89FeKhUwlLt
8GFgfR2uYrE0jIVuAsozefIMcnn6k0onbzSm5V2JYHr+2hf2xP13WEqhCV2A1zr/acYpyHc5z9Tm
u5qm5jU57PuRTeG/jAWgdQneWTOB9Mzi4pOKfhf1SJ5eE+Rxr3bRCoFpgxcCgZA8JqhHTbovd4e/
mI+iRQ/UpmRaGHS0gPcNfCwiP7/mWJbK4b0y+ZchnLtA30xNnubdgYrDZHZcQKTtB38gioHThI1Q
Khs2KsPQ3BMOOyCffQqzPWvgrUFQwpLuOq+XcuuNYJeeKaQfjIsaqiARe9nsMrX0NL4SqKEtMWXE
j23XrF5BRyZ6pl75tt5RTdX76dhPRqxo2ifchC8FcUenJgX0wK6VwtNNkQETpNu2lz+s09sjHCX4
+DDnUEiP6OkzReXJBPDnDHjL3RwMxYZBt8O9Cu4oEQznHE7gYTs2fjUBwc1ET7w7+VR3Sp061Wt0
r4iUpHrYVWhrdGHNn8L28PxXux7wEInykii/d8SU8HI85kQOVvo9SnC6HI092A3l41hZYFDDUj7u
jG+qpDjpeAX36zJIcv/G3PTKOptvOxR9KlE99iInZ+YE7r7UmLnYx6Y6CBRlRF4BjdZVmVr0ZS1e
7I8Ba9E+tEbBqTPHxLoEXE7jKXng1exfpnvvuTqaP3RIV5YmV06pvgC+XqNnL0Ndjj+rfARIXAbl
6Svs9GJqdaJeoyt8F2i+hCiUWsL2pT0mN/WMjwLfI7KxP4xoLrg8urcDsObZa/zk9fgvox+1odl4
qFh/uxNbuaetFMfx+ydyeKvRMNVNZ9o8Nclf/olKTU9ioQuuqt6Hy3zHLKjVziAxCj8NlE4LSsB7
5K0IYZSeRZsE5bRkiMGHwmG9f1tCc3Pw9Q8BFjfP+OVYwr+Tmx2NMDW9Z7zClrUsLFyLm0LyPTfb
LxgCAdoQzf9C/y+p+C85lWW3ITJqkzwRVoqS7e636rnk4b4v3Whx6rYzgvhUzy6Au188wSpdWL73
dK3Eju9wxmXPS2PQ6IFgtJktnVoLj3N5iTawCEIiYqUQPOAqlPJZCrOMzbxONvvg8jO4/qy17OCV
XxzU6iDDQim+8gAJBjWs7wWSc+A+KpfCVAPWTLxbxsHAqTrKU+x/BGJ76JdJIqe/KgdpumH8BED2
aHvOhEmHVPrRa0N3Y1NPy9ChSZY98yfAbMChMuEtt6U1XbFdroO7dMPkx8RYtZA3thXFmZKeHw6R
3Wobs/iQT8Zj7BpcwlpoYq3vWf9oQ1j6w/aGUqHA3NiARDi9GAMNdMOx2gxRgik/ECHfqBTVts84
c3l/KAI9cmlWrP6QeYImM85C9F7aXu21IB2yiWDfH+fG0rGTggPwwGgE2677L4rQHxy8w8ppg1sz
geq55wt8EpkJfCunv1fqu360EZjRZCA24BV4H20lv359dpJfz6DxXLtb9o/8MFA3YQlaDAMBanDq
8Y5gmaauuQebkaoh0jrXFb6tWIBL57HOYF+uinL4BxNyEgHzCYjA9nXWAO2x3EXagDPz9uGBU9Nc
nVG58DAWm1BbPy32LOpz70hz/YPXvCs094GEdXOVa8n2fnxiMSAYg0/8p5o8zfSRuHuHEAQ5yR0Q
uPgWJJ3ztIOHmlkj2fDDry0fHMukuAfLYbga/qWpmbw+3xYedykkKJ7qPmwKXKH+xsOZTz3TfiqU
JvATC57mOlhkauifO2Frm3mJEUN8Cf5aTFTqNjQ0W2PXmLBqD3HA7mp4e9n4cyG8GKTPztHbZhLi
ZVq+pwni1FiovtOjqc05OIfm7Rp0jte3oDTpEIzmDVqswzaIbHshXTUgDHqhSqXA3HaaOs8uM79W
Co9bJL/psikfC3PZ4QFP+0q6L4SSjdVZzLRIAVx50Dti1RPGJh1npWa4Psxp7X9YRaCm+04G7IuS
ISFs9qPOLcX8UwThFHu/puHydGBhhlS4fd2NaLgEnspFRNvqPFeT6toWKgjhIlUwADB2hK0G/5yC
/b0RsofDH3iw3/9BtVUN2/l1agQY2EIqcnY40j81CNoGotu+0GSGL+P00e1nluKEDdhqGiJ9M8ij
nsXLZVvCZobKgDb2rsN1tBzxdPcetqhOBY6qaKR0e8OyaNzeem1LJKLLCkKT1ekKHHA1HR0uUkw/
X4o5ZHFCyaZkjxhApb1iE9oEZ0Fi/QmNscJLEwtoWQjVMjTp7pb+/6N/4g8MyrPmc3bvOZebOVDo
DAcDxjcWDd/bZNocdtZ/fXfm6E1bbSCM/cMSNsylbTDMrm0ErBEiZqmsHG8L1lgpe5guqawlX6Tn
SacPAQf4/FQ/CgIRut4FNE7KZ0ic/5HFYxLdOI2i50dwVAg2peIyXaXcxwsvL87qJkP0iXuymC44
BcDG9+iTf3adUamaUiJnHO+++oxhrecP7dBpzpgfyWEgmJ7CpAq7aNPa8bAC3EF8xjJ8ZgQ0aCh9
wqzZgl696qvK+H7gWIctPUyQVCmpXTSigMNwaVdzZggrdCA09RUdrKJw6CpmOaMgPWez5hrCehxx
52RKee1/Wivv+hjNlThWvyBtp7GzttSweB0jLEqFJRkYvWjGPDoxQewhfO5MK7ANz9e9K5+TKhxI
xQyioN99xzG44ur4iiphmAF7QFhM8T88kgcTHQMdY5ERex3iT017nbl0ZW8LIjIomZnqvo3X6IVJ
nPLCE+LXXp+syOKYwXrMrVErStsdUDOVgSpJdUW8r+PQ56kpTGDvLzFN/E6Je8G54cuClZ5py40r
V2SzBLvHF5B/63M6bXRMV9ZSAxv+QTHhtRtHVj7PsvmA/1M2CL0VSSItsyKQCT6KDoMQzYK32ErR
gJtewgOJPxgRZLtHEuz3lZX8oRgUlfDoCUtaUhIZ8psO1Kvw0qW9GyXlsMp8sXQQsO5JbjvYT5eU
Rti8T/BTcpwue/bg5TfGCWngUV2z65jpT/0Zpwclwj5p0MLrTtkoYkS3XgfaoWKwQARBAofknN7T
2mGmlw5cDnDi8RmhAnK4W6FpCfOGdiZLCWQezp9qZJrtr/XuqMZzXiIrdyd1nm69ISnvCofcvvsj
3E3/X4af5VSd0ylsfQXdSDKAG74iD8iHBB/Tig+v7QlKG2TlgdXkIkNPLtgSZavSfKsyuHTGAkaO
YKSEfQ5LdeOJGOEOgVxJVlTvNc5L3u96RyN8O/iK8u+sULtBeCVZelVOhtSW4tcVaPfnbPL9QvYk
BMAzdmELDI0yxslnXsxx41YjDCd7BJRtStZL6uzAivSwiu1r0Zk11tBBVrhJB46iakleluviqjfL
NYczayol0MDeje02+d/MuzFCQIsXIKkooqCFYS+rHTNPXps3rc7+ik1bfF5Q/ff2ECNaZoBIzSfB
1rd2HslowaF772So1mZJI9y+7iFJoOM5epIVIq9qEzzkbR+oOP0vDGUaSQYvX/1BtWi+Ai3vYrBh
SpZON9gu+7oPMnDyQtvtTfreYyI3s+vRdCNKjx+7RVWzdMWIhGoRES2fKMso//Mre9GvN9l71jR/
vvpQvIQ9kDbW2NhFe/hicFKUtGXXYoa54DrM+Mwik2BH8i7ix15cK6998m3FdIez2npVelH4u0uN
BxhtdKCSQqHXmJI+5K/8sXmjj7Sksd7gBYb5Uxdd3Hu1WsRDBLuqAK7IRMqub0Xv46zFaqupFu44
TnBzgG1v0xtbrFadvWbe2RKB7viQTriUiG7LlPaRUfSi334iy3GnLV/PE8GHr86NJPTNIRqcSlBN
K/XmzhJc//MGEtXbZBAwWbA0BbsvH/KCQFZ0pZDRWzfzmW7NyBBxncSCb3ritCI8LMrIhOWj102Q
4268jQx2H19muWsVnY3DEa71DeJRMKQQiQ6OuywSYRUAZIRd0ZtRLUlvPfsIUwAhhwBZwGoJIeeo
1DM8O1EnLs/5nl014n5ITuB6B2IFiw9deLmu6GeaQN9Jm64sHxx31HHzLy0/uqG17yC87AM7g8w/
lJNeTCOKQU3uo6YbPOcI/E1tWpWvPnw4oDaqHK9PmNF6TkoyHuxaKymakH8jNXFjtAZ77GwgEPwn
9QcacbYyTa2B4nEtakCJrXh9lzsrwnR//poj3jSoRDLFVRdo4mjIW1vyzMPDTB0xp+f0nD6dZMsM
PmUN7CRcMpvC2AqCLuft7f05/7XGiOpeohDBfZfvGsQOse26T6/ODKt5Q/4QPGGvm5eaglOLNFYt
Un5w4HrRiOR8/UEnxjR3o4a9l+SyfEiy2+4tUXdcOt+qMo1sNm33ysPW6x6KiwzMhv4iZRnrr7qn
g+gt07sAYLOMEHbKo4fLjPU40BWEruMYBCy5mFryuKZoxJ1tS4GwIgWUorYe+ObYzKRc2WTogiS5
557sy5EQEfF1MeRXql1Njom4dj572kqHIbGY7UB/Kl2nQJBzVFBiEWX1FyvO7GMSKTbUeKPXm3A+
qQH3KNGfNjybeh3LDcWSrxOlMsr6r+HNhqmXFhZ0NGasiRkvtWwt3emOIjW6pUUOYWKKLI4+RM5D
SUnmVxG8ZZWmYEsXTjxw+0ugDLx1wH4B3QBuaeLGHdgzGs3nuSrT5QRDOb5bIeXvKaIFR07dI85X
LTdBpi0fvYZN1A1iZ3VylqggSdb8RyGHgR625S6oKhw/VrwDnV3ly23DwfF5CxABObL7LsyKaCRZ
NAH/RUcyZSljipsKcBqPu4rT9YhR8Ee0lVDDnTwlfOdoMtzHYvGQlTlvUGcctdE/g51nQ6CWVrVf
Zp9P7HtkAq1T4Nyf+xcbzlPC8tH4uB0noGWFlV+eEX5z7jogzxH5EFZmdkhd0pVSomtHlVyfsKn1
jQo7s3mwJ9PGTCy4+2Qsv+s+7vakvWfHkqeVuAKlvWlqYenWz/GG4dYA9mUi1PuEodb1Cepa8JnY
Z48Jn+TiGlZ40EhIvuagSfKGxXiKuA/83DgV2r6dEd8TteClSPcGCNFvaRfR9VuUQblSXdNJYn10
W6mX43Pl0CDKlckg+3lujjpFnXv5nx5Nk/I9vHmKgPVWEdXCotM7WNiGzH/8cVh7hywGy8eoTQGK
4Zsn7yK8rndim7d6lg32//TbXAH7CquXu2qR/46rB3ILdhaUf5tJ8NNb88u9BL/93sNY+L4wTY30
BVPpzfuDFLm+50vm28zQn5pCMqLVyCUi1db8z0VyEnHHCLTuk0a8EOtWIVCGiuqK5XZvaJeS7y5P
Y0e+jhoN5JrlsM0Uxf79VHUhKsPn5sRo3/MgVnqcpz3wi5phKUfvkWMZ4NhyIV9fm7nvtScyq1BN
GUKceY80GOaCiIBQx8FljtSRt9Si/Cpa40FIm9t59dHym8AFxz1caFEesPqwX+5FTzY77gAIy0G1
w9nTb3NynzD2F2yoBbHy9m908HBi2ifP+2JAjTRCk/XZnon1hnBtyV3AWpqrvrGZEWJ+d6955Q/l
YcIErm3e5yCLgA0/wEGAqOGDCKoVVN2r97GhsJOL3gPbg9OBWMZ7z3CW5A126YuFK8Y6xY7rDowM
G5j0avqDDLbNlBelbvXyiaggMMUJEsf5bk5Mam5/5JY92dE8ip/fmY8x3w6kTx/0fhqY4acUly5K
6vD61tt+VNqThW6biKoVWY1bZSEXFBf9as3EQPldaihQrmIf2l1zFtyEggfjscPTt8TU78YPngs6
0S05Qqoh2QCrwadtkQKusqzIM/Q9Da3EAiRnJHJma9H9uyN8DBOHNBBQTEfUte3WKV0ll7kiI9t9
0g/z6ZkqN1icrybI3Q+0uTPYDq0FTJcteHaUReaG4cCGx1+2dSS4y5tJceLRRiRxdOh7rsVqU1Nw
LXSBP5Tqv/XRHWaGvW4JkIghSX796iMSPqhxRwfllYI9xcY7PVouc06tWvFWQXxtWgmW7ryQNiyK
6Hf4vn+8lr0/EFaCqRmUgEm7CQj5ykee/Vg4G9Ihyp9lmcFeM2ADgFDstxxIrbzDGpmrAQZsIsRA
ZcmoZhpqXSkHTV4GGEHSkSfDxF+JqfP3D5m2rthXp9KAQAxWTpttV1Arg4x6Rts58f7iIiggBSUR
q1hRClAXudvifwpSK1dJFh0p41vSX2pouPa48Jd/s6dFa3s1puMEYcF1ej7TSkgwzn28AEIpKUmF
CUy9eFpV5hrukyDFKUgCpMQmvX80naIwHwgTi2FJ3LysxVAF83FBEZno/p0EQp2Y+zSkqL6pm7EJ
2kBK+zKNzqqEDAsF5h1CYnbMiNIk2KU7aet2HuKA8ZvUFMSpKm0VR0iw2KOeeaptcRhp/jZRJ2n1
tv5aQk0DvhpWnZ3U1KMRtN5sU5YTerV0qREwE5lEppEme7giJDe9fgWhLsMDxKOzMfoZrfOLCXgQ
isdVWakZRAliQm63qg3J29sFjNk9mddaGqubD8vGIcee+6jeq2SrrX9YJHI4Ipow8qiBJ1/ewk3/
Ok9sc58o8aY3kijAYLVYCJAbTTSbZenOFRXIciiblDjqsdg50ZivTcPq1zpuCWLxwpSI2PRsW0tQ
pSYnSufwRN2Eh85wxJvFbob0g6VXRVJvlAHiDBmnMjkbgqtkJ/yvXHJQLHdc4PMqloG3SFe/d6FC
8hZY0ERWftX2Jz/YG5+qbfTslbwcWCcOLyyC3VXXpMa668yMMCQoxTLjZJWYPRq8UNwjqNQiOOW0
1D+GX0UQeWSbSQNNxKRMNs806p8sD3UGDSm+DwfMlwg333xfM7yQi+LU09WlJL2Kj080v2srPeJB
k+XZ3U7NDdskV9oV0mknqPLILu8EKd22sCvkb08ZMQ8rT6odMqt6fvpjw1rjHmT+4Ekhh/8l6ht8
Uj1znfVz8a04ZxwxxktFlETibf8QJVZsQ7n69NWhTQ4DE4y6XyWKfOeLWMt/nfpBT+j2zXs+Psb8
NH6Tv81PK3gb/5508mCu0nE5wJRgnjzTKDK62cAyGrO25cW6r1NkJOj8mbzNcMnx8UU72FtYAQoq
F7RsZBT3QvVSGjk0NAdr0m1bA3ZmZsW+vAE5HGWmV58IelhOFVN1NiRvBnnEV6wB9pWJBiII1uWO
S3kKQNEYbJBdfJy8mnR+kDw9IoyKHZHvuOrjlhUNg2hB8/JbTcdRRTYNIi+3eByHlZbXsUdbAJWu
qfv2I1HRkVDyvE396E3mK9aQtmH27pEwEU88bMcDKIPb2Ubfe8hR+3DKiKfBmyD2S2PZwjF0oWlj
Pw1yQo/CteM887nLh4XitxiRcuEX150y12ZNITyroxBItxz2gk7jQ1OR7zEXpiQo+vQ1VhX5fSnL
YXaz5XOHzUjXHZ4dlYlmmLYHx9PKhbzT4i8Dwr5RTSbMp7uVItmY3EpW6IoaAFGMyYM2wDgAlScr
g6ORspo4Y+NmghJO7GLiEYhyy0ke2z7gABpcsdFMjoXfRX6HxV8f7Fp0MXYkDz5Aa/AEQ/BqsORF
X3CNWFnmaxN1BAiWHZkdBNUlShRpkpmAuBQeimQcvKv9g4iLhUu/bPGpvpIHJcF09E5GTupXecj5
vAf5QCmhTtxa5nBcGKF8jLx67EED8AsC2IQB0pEBdtUreaUXtnV3XF1Ial6tHl0q8jfuV6sm4V1E
hif1BUy0gjFCX+wtyUlbvoPO0w/lUkRSJ2rC2yRWb9T997oM+xHHLIXFVpPrH1Mdvq3twlndqT6N
pHdQdKMacK/NKNEIqVYKx8MK+ej0f6srut1f07zoKNOcD70wTZFVV6xhZA51usjwmWwXUEj5YBsZ
tcierl+RJP+T6XCTsPWP3h+VbB59I/MMAoJ8kCJIkW6joKMobli3h3s9AVI/EIbimzQQcsYPh/qi
GzeJV07iYToD7OXqDHIMbyaLjoG7geSJ6qS4wJsakFzhRlKvmIVe/sITy9GzBftljPT/sfBNBlYg
B0u1vXt4+9X5qKqxOF6UqiSXVZpcWEA+w27qlqAs+hJg0KYk+i02UrwK3Km8RXN5yBQKgD/0OSc4
iOfnTn7djXZDosU5dSBrWKKZ0ESWOYqcXhq/aHGZ9hABEHcU3d2hIvZrSKh7nZwst7R/igW96V1G
KD7C/5WFvWHhi24YfFXPR3YydCpHVu6TeOwQG4k5tQynVI7YbQTJBLaOH8KxF6u8ODNBTnVKTWmT
Ckdb7slXz5VLXSNpbnADbj2nx8Pf42cwraJKXBtVvs4oOxgGV1Rkd7G++SSSvqkskf8mkbT34s3I
MTWvFpMWr9sbLgDYm2IpjYFvKW/9I2qjXvvbZl6wHSR6yInrrjVweEVQesMxfx/ClOtPzpaVBed5
zdPogo1uJphFoPxQC8mlg03AA3vkJtjedDpPLwdX9j4YMNCMQE9DTSTz+X57fpiq/w4ltzhehL7q
YeSdahDtqC0U3BAT3ATkzRAQuVu0or4c2G/Hposeq15G9p9NDZCPIoj/RYq2knMGJYxSUbeebCIg
ak1Eb99x2qEHrKkJrMosAsnvKgdDv9T1CS0BJVk3huEFrvainbf4TmP9Tn4pn+k2ghe2N2p+vs4A
Gbw1YvVYP1MiQ1sRaGVHMrMGtddGC8XbXaahjA0BaYXwyGeZT2dcd5oQ91czNOmGNpojH8fGfO+s
lhyH+z6vfJSKRryiWK46Bhg4Ttzz+4iH3E4f3USKhoMC/XqpIt5aoY/A0zKsfMFPdvn0A/4Gi9F1
MF6u/CJU+6RUtuEAfHWlPsTQHxdJ46Y3+7a/gWAceH0/kIZVoOFkFD6mZBhS5CE5qS5uUPOzqLPp
HxcOVI646NAlhBMCRiVrw3ZsXFn3ZHJrbd/K3/mgaN1oH5leX+paVQUiHV2LKtfgADW4iR6M9wEW
9hTRpQw4ZV9ae546vAgE10RIkRlErNA7CVLKzhh/eJym0N449yEhf+d4WIF9eyxa63J4WFeO6EwW
IILBZHs1hc97e9WBbDbSdwxMjxAkXYsfdAntxUREQ7NjLBU5y+dFXzZEy5IecZ66qCqxM0wJ5JfQ
nYH2hgkZjHIn3alf0bMPD899zyrOy58Fv5CTRR+vXjRxIbkvfkTzgWHeBlDs0zBWDJn+OA0uZ5ZN
Arjh3wJ3N7kuVMkkaq5/xumW8okSHe2sQ+hfCIz1rly6YMrM6gFaNXCVvZ7cSoJ+R7JP6c8mgucb
NmXJERYAduvDmrKZFSVmECA3Ob887mLOLqqvkMWzWa30UmybYPQh7/9pXpbtvCRjUOm5AlSXiSvx
jZi+x+jbArKO7dM4j6doLE/eTHUDpGFXMMKh4ymGbYDVD044DO1YXo/SaAlPy2No+NDS7NbmFvgg
oc0K/NVkQLT7fuQILFBvnCidN4mVCkYpKtmVuU6aZUXaGa2t4//Z3JjtjWSzYb0YTVvq95Mh/MOD
TeBoDkLfpmW5HQ5v12Cp0s2CQmOLEFUblMJyzEFnNvPua2qACOHMpx1L5XQW/0c/HJQBoAjuJCJb
M0fzL6+DnY4ELp6Cjd7nDcdjA+QyxvPIzuOuTmdAQ8GS05krg0aPj/8sOmxsT+t6Il48WdrY2mIY
JT9Zo3PiFKGKh66Asbow0gzLJG8XkiMrn/+QMRWirz2wwHgxOOa5ryqF/ELfysXM55dERbxlzNiU
g7KTwoXNwZ4VjAVY4CX6a1L26QhFKxscfwTO5HUZ93MZWKxWLMg1yyWE6ghOg3RTuai7FaO9Is2z
cd1c6MpOTVTSZwoJzTiqT++0BRZBrfFUb58pekQdlCCywzZwMEAib/MhVbcBIOf8w/FokR8DvbZv
dnoCp7QZDvahEi8SsolmJWOL+lRt7DpFekq5lWoWaGqXz0nwj/pbMvnSwrtxQWVDL+D2bYGlyUhu
NB/yn9xnpUCZ4ADFNl73ZaV0P0rL59dMRiczbURCF+wx7C4Raf7xfvMuHmymOFWYARTpxEnloZhu
UG4MnYcEleZ8rMWnG4rkTa3hfKeKhSnnYdE/CbzYkvdPdEGHPKq+DPbnpn4ifqrEdGH4SqeEIsPQ
lRx8S5pLgCcQ5zLhC9mmKr2DO/fhywJgJcuL4miZZEbcslb91mvwFwtZE0dcFEff/JIuZLtsJH9V
ftHVwlksyNTtQfSkb1wPjuRYUJDXGIc/mfSD9cqLFpiN9oThCS/NRU1+lIX8A5zbp275YQyc+tfR
MN5NgWkVaFH73hiamTPUEB115UozRwpPizIx9o7d2z0v5Sr4CWzoftL25e1YFwlUhwU2NNRHYOTG
F3ulG6IhzDtulA9Mjan/eyS4fKjcU0FushofSGeeNPEzjVupbJ56FSFdypKqqAgEQP6uOZW49q2h
M+MQYhfX45sVoYk5cgyL3L5m4kdXKA3fowlhEiQNuxQzi5iSoo+aIZ9bOv1mX1GkwSizQ+e8AK5u
E2BP1Sc8t3q5gwTo9Oa8AqvnREpw4uzPFfHnBTlBPZ3zU2N2aBmOKYkARasVZiJvSNl+l4jNf/NS
sOK9QBFILzAxm7/4/8P/LBbiw5BIRV5Fk621wxbY3HLKdSHkVcaF4n2pb9IAVeHzzHEC5/EMyQE4
BikORN+IKGoaOxxViGpcMGGEGa7XCJYTokEgsamoZE79g2FJBvJDwBiftqWrrKSTFLFwvzJhdnTm
D2kFZu4pHqG/hzX6LnQx1spsCic9v4amLXH6+PCMNE74pIcvmS1i56pleSFMi6vcwYfBub9HlaCQ
/4pHtOZhz/9tsTFs5DTtX5yziryHOBQreKS1ThyhmlqwvpCimQTbZLJ0YZNf1T1+kNEGu5Xc4H64
VMDN6cHdR/y/36xSqw+rPGQ2nVVNEKqS908S8ePgcS8cLfbhQQZgW5ufEliAmBFZdB/bxRJaSfgT
V8VCqKKAlXZ208b861PvHImD42wN4XzluHBXP2gs5NcjLPRo5MjjvBl6te7goT5gdDlvhRuhfnEQ
c0Va9ehQkdfT0yGdaSRCgf8Clmf/Pv5wZH8jnBynJiJoR7i/SlDI4akOfceRayLWO5W5wPisrhuD
sHJ675aYpkAHpZZetIexR61AC8I55gdtvpqD7Ra3lb96LIv6BI3IoJlwGbbu5I6y5g93ybcTtomq
sHxDOh2v2qcO2wTm9MiiVLY0eHgReiQEL4mxlRbxHq7OsWKGu3VzCp82MOeOxAmGBoUhj2Y/AgCV
u7phRg8uIirlp8SFVUudhXUp33WoarMSOn1IuCgbyNWJ6U52fh4H9VlC1Nd+uT0jvTr2aOyBgZwL
vdBVKcbgpwDyJcSh28z4AtVN6r/rNnCBZujkxI3eENJvhHiiBlt6XvFGCwA6Dkhg/FhfHqBWxDdy
U5QNIHeBNFIA0KeyJaITJf5NrS1z3H/zkpOR6yZ0UOWin1lmSVbE/4e5D2bZvTxqdB/oX80W8I0J
0ko7UxkCmwjnHm/QhpVUdzmAkcaC0xZdAgeInZWqYuK+gc799G7Y7JrmEvVs/r/yU/bVkLMS40t5
KHr8W8OmxU7FLOTB1APsXzBKMTJUqNS1RGMxU8KoGm+TSlAo18FJGrg64hsuX6Zir4XKLC0Cs8BA
VJFFDrKHbGAymdlloUgu2TAMR47dP58Vp0RrKbbP//5ObpysFHLTcUNhDihpn5JzndHcDztsOoHW
GDsLAkCgeVRTSpeZDDOVrzfukbX/GSOplr7lTQf0Y/LYox3850DdbWojOzoZD4pV/L8QVmfM6NWO
NlRT1hovY0OvtnqYNuDa9eiz3GtRkqNSRQxcMuJqsPRm4PSgjJqbVHQz7Lr0MYQDjngOxBPTvucj
0dkFPPgAOrLkvPg+oovFwh28E61C+VGBgenKJ1RzKCivcQqO/EVjXHV2KomTf1B+CV+m+4qGNJf8
RMJSvq8cymFJy8vPtoNgrRg7Xeu0WL3c2fEyZfGYOQ4cs4pskKBTP3D2j4V1H1AUu7LrLwvwZwSt
UCuigqb+s0vgmFiPRunVrKm65NzQ5/TKIzfYpMwSRfpvTdnxy5OHwxH0ZNF1GnS7ncsvDMkgwmio
WPBqRkFQVINdbB3eft9pb5IwfOWVZbbEeLQIuEgrR71SnzvHeI7ko9XGcxy2FUt78pyGyJgOzEYq
G3ufwX+ejBp7+MNJX9bonDvfyrCZXrtvL7XHTXDZ75Nq91sNFEubodVlf8BBgP1BScF1XjYWV0ZK
kvXoC10LHbF4X3fklE74Mwt8OgeRPUSI3/ONigxHt9caLja+grq5OD57uViaXoW61NGLxf8OKiMd
PlGi8grludvZY9Gt5zrszJ0NQpj8ewHqt8tL1fP31tRo3diO2Bk8AO+LDzvV1k94QNKFLBZcnbe/
RogBlGIu5Q/GNNg+/zaPqzfnvSqrvVvJf+GFAkA/7BrO88HG5UDqVWpMaNPcaK22/0A7CZTA9zF4
BAMci9pOVutJ6/wwHl1xq7jHQ98pwiRUR0ye+72rekQ/Pd/B/tkIG0AhUcmY2NzEacbPTz/5rL6U
/3GJX4h31RSVWzi0NnDanRSVzEP/exStycf0JCJ/PPq0iI7tGZxtgxjjAIKLJFi+8Kw5a2jGQnsB
iSQter+TUzEJd+Ux9VVakUAPlB+uVPxLjiFNej4Y8KaorJIkVaKEMXgmUTM/MwHbxDbX8+sQNu64
Juq6NphsunZAv/sk7p/841IeHECTSELXd+Zu86uUZQmIpKIfjPAxvXaev1XNmKtEnGGkCIduNT5N
MY4TKFgFI5aUVk+txKTKDkARgebxej5hcYntVnPZy6g7vTByYGWH4D6DbcF1O+pwutHoqCf/9XWp
nD3Exn2jkyuV+m6tElp5UvyqtS00v400Gh0h6vr/+cyJYfr1sMxeueH4l510vz623pTRf4tNwQt6
kbfZBqnklfDQRRYKpWy8YyS55prrivShDyr60mLYbyAjj/gcGxnorDKKknW3tYT6vMMaGzU7eRuz
Q662ag2kC+0SFlzeqXv6ONSa2x/LyD+pyaQnpeHCiziX76HNkj9qWTaVFjN8k9E38MvkOx0ma1ce
vR9J8MD8tWFlhpy0qdmHmyD+IgkUXDv26rG0Fs9EjNHM01cPrH9eDae0ljEy0uALm2Itf/OvuPPZ
lNywpFaxOX9U2W2mISGqrwS8Igh+rVS4iZJwAfLD7lMW2LKoDiZhzC4ozD7qeRO4fkdeU7yffxSx
ST8isLSEg/a7HVwWpb8gFSM3JwaETLksFpx+r1VSk2ij+4tt/rRDVUOo/BFcdToq2dpK75eKnueJ
SueqJ25q9v2nx8GHefB94nrEVTmLi4PoiGG6sE24rWMm2HSn2o92wNM0WmNXbW54zTw5CHiW8xgJ
BnHliIdCciqa3OgaK4zYt/hBuzPmCA5g9MEpHTeX468JHca3D7d+B6RODUQad02vgBUxYaninJKC
BfaVQqZMTpPQfjro95AnAPQd80d0eQmT+Q/Y0exoQPLOFPvt8iHlACjrkiPJsYJhnsXkLi9u1Qei
UNmHnwEZfZIOv38IODXdGZRvN0NMogm9q4FjQh7dLSxLkZwh4Fv4/5KtM3oLd9x8qiyJ9/eEdwc6
l5rU0zE1SIDsaH1+TQYZXp7+eHOsIa8LDydrqSzY4m3K+VTl7shC6AGe+loROOWKzQErHGH4WSkV
s5ovTV6MbWFMBFLfpDCJd3qEJW+01U5zfejDcvA1eCbNnl7BPHc/pNCc3OenA9UTDL+Ud2gg2vjd
2JWHdV67RuMMH/1nhNzAkkGrfRoAUR8on5hRsZ7q3Ncm+ohBhFQhiG45pF59zZv88VBalo07KrFi
NB9VisMaRXULqNcoOTFAXyUlYTI0QEmAOhjSdfx3n3D/6i0B6oWuJgiIX2+qGEAGfKudwzrG1Vox
r7rdNV6vlDkaRofoJyibE+Qrm2Yn78Vt8ps+ulbOs5RAhMwEzacckgDC1B6Fg3iNAJJsFWe1+10p
bbVo/+o56uVGPlfEnINhMunZmTjlW64OqPJGLjgfGFdmfZOPO0i7tzuwUxUkiRormqST0ZJTstGU
aTFi3dgd1zvlcd6yBeNO3jpO9yHP9bOjudfSwgCvqnlwvNiq3+kYWu6xTlYWiT3h/Dtu1IR5W3yi
N6tGqn3NIxB29GKYM6ZD/8ALq0Hxj/lyjpLbjbawQOEk5/FhwMGuCbewrCVKT0Q3TbrL0wdyNJQh
lJIgQo7T7sLk6pQ0c33JXRpQPMzCUK7l8FTZswkmSU0cfV2Va0r+69iPqsBBB3oq+i0+WbOBPE7K
jA2l2tIzr9x3j1JYOGoGBaBKznAghWgrd5eHlHSEdRDU42GQ0oBzFWsGbOii8H+4EWc4sxTieHS7
nabC/OA/62BGeJ6sGEJfRT4BnC0jRt01NYeI132zygMtRR/s/SuM0F3g5HS3XL5eqbmCnTHQQ19k
PMSaRiRFUj0BrJ7kCFLXamgHJtKgFf0VOvY4A0PaPGv83HduA13jbAJAIpNaCIBGCfN3M9rzmKRa
DKO0bL63hCnQl2LkrqG58SbaIeTdvEyv1J4mICVoINoVuAgqbeMXbPW9CkES16NR6196VrTf5zK1
v6gNWEc8ymliFtbmixhSAqx9+PI7PmD0UtsG+M/4x+mhpqXKloar6G7XZiIMsHgDt1mYWeh3B3MJ
j71ITM4IwCKUktn24CQHE/rwn/UoVMYcbPt/ndEHyuqiKZ6njb7/kN6lhH8dtj7OlGmYjTWQ6MN5
6T59aBqoLqArxx0cS1S9aIqIeUK77RhJSm3OxamI4/7rZ/Ix0XXMWpwI/Lb7KH2jWyHKfe2HDY6L
OaK+zsFeHwaD1KqTlFyLGw6LkKy2IdJHl9tg+8YJ5sosDA6Tc5EpmENGSasRguujetvsXOGyecL1
QbrkgyGd5VYWUzp3mKKo+jD/GUcwP2c+r4L7rDMHbgqImkWJ8y/EyFvsKBz5fb0WPQ7q2555pcQJ
kzXeU8EZjU+6knnCrGz1dlvIw4GM7Vj0CJvKxIiLpX7u6KKEV9+8s4gpT6Qru/633o9sR2b1nP9s
Q4nXbFaq6p7pgoE9z50oNzTCZvW8q8HaQ+PAKrfdEsKur4/2sSX/cGXI7CgAOQA+FXjU5dMjOGuR
30L9TuG89U6dnGTrqiPgcdv65573zbs925czkhdYLK+p528Ew5sXXCYdTLv8XPN0YAvjANEgjiEA
U0+5wEpZhqLtaZDyahXZaSnM+sRrJ+fjFdbMTfcylbz5X1qRocNtZyJdFGs4Dh4CZIPIWqC8Jj6G
oMR7S7kkfemzlijXs+YmwCzW9QFpDZrmD8kVuXRe1xREGeK6Slznt15QuJNVCUs65HeQYfmZMRdN
qczIM4Pn7LSen3oQonwOJLQadk8sZ+0Svx0YndildFdgB98HqibLNk6kP/XVYpb1MxWU4nnxWhOC
RL2V/kGDoG8w2O9cAYRlVXoNln2LdUqmPe8VEm0kWybEz42yAOXp9Y8T1kyxbZvTtjK2kNJF3Mzs
xLNG9bFzDITtlbKEocwrMFZ4wBUaLoxV33ZWYbnZVs9aRY0vAuCxKUqj+IPQW5SKl3mdxt5amxzI
qRERkjk19JDW+V5Vjfzsv+3XxoyzMyn5TVnj9Evr2MZkjkg+yoczM3P7PcUa38auUye5K10geLHb
CeKo44yz6k0tqjmf8s7g9M1szLuLoQyj1qJk9UWfJEywYlzOeB/li+aNaQRwNnN2EFcJKKsSuD+M
mMCrkOsEp+gL5d9Oos6UlZ2LTNQI9o+b+oLRctjbfhNDmFpJBsOSv+122FExlxVrJCntOkRxxqDF
L9qycq9+XzKUe7JaIkJp3pq3iC6YXeXbxuPalTaAsXK3xlFAfqnlE4CFNG863d+YoqcFV4+PN79g
l9MR9pNnj5SjJvWiAS+JixOl2tH+4qrqmUbaSoj0Ln9sOPvvRIgL5eJkELxgYFnjUd2hN0sOFaZV
cIz5ylFxcmOueLiyQwadiDVQLaDPA0BcOfjb+Vv6KWGwvO/0MLl2WB3JXkh0+JDDHlZ5guhPdkhc
Fh+GlI/IU2jeKU2/zgyFINoAghOZPLyq19cW12EjOn/SS7QMA5X64D0fg9vaNuaQ3lP/sv0gxH5w
vx/iURV9AI90YhSixdk84NTAXcq8UP0j0s5ov3kFeHodQtzM/HPMR2L6VN3yigPeWXrMLq6B546v
CPWRDF+/X5s6IBL+KxQfWK8X+jCLhvZ4gnc0BTTwBzgCI/4JZAt8KJuLMTC0QJSKGUylCpoX6jCZ
jUih/AYuOlnYTKWnzQwkqjQzi0WCwyZg7TFGNP1PAF8vXO3NLn7LZxkL7zH/kjOVyOgqas2Tov77
k6W+W1+iXbc14u7YYD9+uhntwoY3yBMDMKAU2rG5OUQ7Pt9hnDFNPzCaX0ydbLRFQr4ARUIeULLp
C/ioYKvuZxNumH4JbHymX9CQTQ3XP9zgwpB+auV7vvNQIfBt/dtli6esAhLEFvply5j3bVcNB2gD
RwmY0tFrb7R3F2dC8mnXoyiQjtIiJgb3Sa5BZgYnYnJSFpMiTqiQGrSW2J1cwqM2Cw0svOpNEYbg
Q2WF8Tvs8dXjkra1Fna1o3Vikl0c94xgrQ0i4bgeNm+7jDWeG3lWvpS+Bln1DSfra8TFR5eiYzZp
Q70ZCXd+Hk3b7whC5X7Mb1LG4G7z+Gxdv/7+ltTJqf+3AoZoa2oSYjgf/SvesuWeZaon/akMD7KD
ncmM3hI7X0nsY0A4+8ZxYq+N1HTw5CF/QUMoqUmxjE4L8D23HGri4ALfH56t6lLj4qKMrQlqMXtT
PzShidcUr5W9R70w/NWrqSjKsXTMm20AIjOVGIJ+/i3iEQ5vwGra6n6oF7Fn82TlzdVpjwnAfE0u
1Uv1GXa1sNYCU24LfVzMIPKohJOTeuXvCx6EVkeQHoQpApv4E6qLKbNN3LWnd8I1Or6XB/SVtqGz
EyzsWrkEeN+jifNBNdKp7/x3YDFYor2q3kH3+MHPoH0ojfp/h3TSHvPA51JvrGOiO/KKi+ysSV9x
il36paHYfzUJ6gVkTfyhUG0h4pbtyyMMgt+O3UbkSxhDXlvtjTM2HTm9F2Yvdz3DYJtKOrH09Khr
ytNef3rHGexN2FsuzbsEddNLHiTexPdMfVYicgz/DCO24+Lr8Si6fcvykme8cJ0DkpiGdLG5C1vc
AcbhNkQqYQ/iK8sHav6zWvTlLOknw88HfRYnc+Nwq/cHg7A/9A3FrXGfTaVZEwKFqReZG0vGNZrT
088qrpsxnczpXSQe74B9g+oGFznOwSdP3i/x+h0GZBMaPWrdlYZo6dLJdGQchneZB/2MnMbml4rs
boaZnP6d52HjtDXyoMapzTHx/MB+jbRoeLwTigNZHKQBWaV+rXRpKs7fTK2iHl5oIbwlxLsneXqO
3LkMmkitvFkhSSGpfZ9dhiQfd91YKXu0p8wEIpB5E9OmWwAy/n4ctgU0n4dRqUwP1dcSIMysicFX
bi5yar/79jZ83appm3JZ6gO5T4XEeaKn0yZTsdN+Vj8OlPp9v7nYJnrN2I3gE6uO86X5PGdqL5Qi
qpQpiPOT+fXEdgG/euE2flENc9h/RFaqbGfINtKS9LSejUNHpek3eB7A1YQL4udYLrGIAh1gz7Cn
OFAAwoqeesg5ZfNkO5uv3W746WTWxsUi+wtMKERuK91bLlhvHTRH7marodw7jYDw/D721EzE5ZsX
eu+z1YrjKEJwMRNp1ElW7981QZnv5B0j1o4n0HqJwpz+6+SFf7ZbbU86AlK2eB2soq9NfpcBnmm8
n/GMnC+/Hq5g2TBzDwL4EXXxOTMRjsIJSakQKs3yN8oAZyB/mirQ+/PMhWYb6Cet/UKCDgaidtKx
yqQqGgowr0XVhx2U8ayVZKYSUhdPMieVX88LwLx3aNVfhWsD7KAEJq9O8+ZvOkS7hPJoygrk0CDd
ou/2r35qsZld5knbObHNJDNs23cmO3d1zGJV9rb4CgyA0Zj+iKKuss888RMV9/mnEh5eaHzZMRIO
3IUOq5vVOa8lXxjrB1d4efz6BxDvf8KUIv2QuYxW4tP7Es1BmR0mRbT3KtGYJJhjpnJab8SUosCX
AuTxLb+bi+t5z41fUxVUdJqSBkrO6e+O7e3h4Yz+W5fwLso5knnuB6pMRNSsiFlVVCCrNZqCY24U
N3FQ1UtnaLYf4BGw1rW+XcRQJEfqOH70Gh3oH9SwOJLGiU6mO09Qw1oIpam+snVN8LUDUvu4pnJA
59wiCeq875alI9OTm8JUDAg6kvyKWAH6jxmRRro91jB6rYxP8aFV63LqZoCAdV/QgxmDB6QnffP/
/7yK9YMn0PQwVNRRWrKm46vUQw6s7pswaFAIWAtAGgA1rxSVc0IXS8Ne4JDk1fOhe7xioYv+yqrU
NwIngIG8GOQPX7nW0F5fOHNtNp005ukJPv1/hvR243WyPP4JiwO4TUWWwxU7A5YdUTpOTJMhXEgc
fj51mBjxdYNPG3kU6FuaBB1Z16WpyL3GecShwiH6OK/SsRVf8ZYx0z4BfY/66iMW/gERDq/z3ftv
TAARWaipMHeB3DNzBoyWEneJmv8Apktee45Nh0BV+KFW/58t3QWVurtB6AqJlIhgVCPsi7QcIsIh
eIr5dGcctwGhn7QPlGxBazLUdfD1zCpvhem4xIPrt8F4JEYU/DqgyqBobnMcu5DlSW5xo85SSuY0
zZvAzK4MGWKZwN6uxqB/D+0gHJFM2/rxmPbWCFGR5RQpVST+tsIJ+rJ356b87HpLdUDy0498+l1L
5lyyBY3tKnE1IJvMeiIbUgfyq5/WlPC2K3nwcFnJP895GKiTbhWcXzv1ZbjiPZhCB9xgN2pjFFyL
sTBfUeuxw7YU9Sq1v9QKcFQT146hzMMEPL/ePF+PIUE/KY956n1cMKXjrVT6B6nLQH5FoHmGJSQ7
xEM6alGQ2gGglwKEZZiFUtfGdqFxKeYbVbZ1cXxkNmqL/VHG0zMt/5ZHMMxzWZAP0luVpeUC+x+r
XpGteXDbpzC2i82hBt4dayjr+zlc3/P8Oi0c8Wva9fjFuP7ehgDMvox8ZA0jVjj4AKKv3h1GdTaP
NTKx9fiYh2d70dGrMSMb5fVkctDC7yTZGmRC5BfvYUn7Tbrfawq1lNKPwIqU+ca40RiQCyqHB2ik
Jfr7RIaUycTKZMW2JkD6Z92VULF2tdhCMfLlj09Zb3AI6nstBCIF6OralbgiecA6Qqao0ZkkFMTE
PxP+/0m2nP2PWykz6mMGo7xmmOQxpT416BR8WyGzcP1v+/l4V++AAinfNM14ij+U1SJwSrXLNwjw
/1S85ZqBCQHgBClPzIH1iSbBxWHHHJK5QZZpc5m1LxYi6DyYmubXo2n4fT/en1B9Btft/1GVQKt3
zt449FJBlIaJuMPiolPVNTNe5gh4ERjGliPFuVwChUIXc0C+K7XbzRr54tME9gsnda4ik3E18BvG
tYBi7DRruue1vwbnYUzlmpR+bpgaGz64qDAm26jy7356FWXpa/dy6xRFX6vm8CiA2TD+ZRhTw6YK
CPyPadqSRpky/fjx5+N/cPIrJoNCRO/KxalDGUcAyigDGEKpXr7KHwmdM2om09ROgdgwTCzvyac7
ymTQ3/2I2b8hz8UD1qQIx1U9wC1+yNRVZ61VtsMTVmpjkGnwy6P90fn7RgRrx40WXowz3cRS3N1I
4kfPn9aEc0a+AhVQBZ8DA+DnbZrOyIyid3MDCx3K5GwoTSSm8gFgkl9gKNH6nKoWlX4+XKPLwxXq
gBnI4SNYT+JukcVtI27C078F75tHOm3nFdnPb3T6CqdWL0xK0ckCQLMhXWA38T0go5AghYksSoEX
3acyGZ+phEgZnQ4/661OJxvY4abbYy1eAJc7ENV3G9TUsJPEjlWJhL6etW7ctFP2MOaXs+o3/PDA
a/lZb7n6PJ8Y22kpH0/oJaJiy5FQSjePtZjB2P5+BTYHZis0qwVHXIRzt0XMOqw1HhokGXCcvFMf
vlBoC9AyWJUDGlL8b0YCIWKnfcSPsXhwqVt7U5emvqqhi7HGJG9D7do+86JJ5fSZyjDDnpRqUt6F
1ad2r4ageQxdg2T75vwSJN5UukeFsHC5mYdHDdK8yD5+8z1wEkN+dQQcVH+M3fcKUtldFCORLNCJ
ejaZokbVpRr9lPqExrYw9EP+f2aMUpMI4UBroc0a1yZzEg+z+AksryECC2PWwKdx7JOR+YL2C9Ee
fZWPKhx7Do6AeunB5TM6IT4QMCpS2jy1KXZnZxgs0hOSsZ2c4mIaGzOA7M8XTN3OYb4AkacLVlzd
1kt+V3A0pC9Kxk0kkPF9+aO8Rq3RIloyMk1E7wuDDv1mXSPnGd8UnBhkGF6GUWa7EA0lKjl0gNAO
rrP9fjep4Pq1WJnzaZfxmDr3xQtBAuSQBss9XaqRa6tIi8Wrp/Y5rv7e5OdQPse0Okc49t3wU1ly
DUNDEib2J+4eCr+j8mzaYTczcWKCkfDP0UcdvWqCYu0yGADrBNzY6XCcaFn7O7acFOKkw+LN4htl
0uNFfZmtuppWfLop7WxXKhlA5y2zPs/W+mcN2O5ny/xwPOZJzwep6go5kPLqRaKnSpLJlgQkH0nu
GPGfjS2+AxYQUhgrc0ZS5FN6mY/CyLjOFDuTzk/JVM/OgFl1qVLuX1UEzgKJNAj2+EaAw+FTXKVF
2V1dT3YIYXGoLvqacVTX6wDMHEQRZjSiNunXiM+6BwaHf2AuCr4EQowGFjvlpRhPMJl2OSFJu6xa
dL4agkPdqZLle3jkAkIDBLlZQ9qc7VJxXBpQaiFdfYn9utIW10y/SvljlygEQ6f7S37h6QoJS3OG
FwjH5KLvi/jxM0lisbzOvx9495Gx6oZjC1XUVoyiAuxeFDtepzIqzQ7pjNeQZ5HRgbXLH+bQS6f6
jp/XkePuJCDoeWD/BmSne7kQSF/bTy9fQWRCl6//OLs3gpjWYZTlirqJfakYEgVTwlejzxr4ZQTj
187cu07M69V9xk4x2MLxfRO6wYjfJ2jh3wfS2VVXiR3AoBMSRY4d41OuYgHwXor0tBm5O3X3l1dJ
PxRUVaS0iZ+H3O/+qlcY65ctL2KdhgYuptB4h8aYY3KAhMprB8nqygOT83okFqdiE/MZfhruConM
HSmNmiuvhj2Pxciyr4cBjFWW2+tRBxdntz+HJ0F/azrtYW3b6qXv91VBFX6gwT3nlR3hOjMM5QEz
GSnf92lVWwkijkEzH6klz76oJeF2SVsCOZ6rE+fUo1407XHhQl1IE6UhZ4SUzK2nK57Lk9NFKPrH
P0bKfExp8CLlKJe2F5wNdneqGKIQ8VtlRO+C4IWxCCmjKhFpX6Za6kxzEgaGF/Egw0ROXEio9gug
pr2Cc9afByntm0otXvnEKaLYD3KlilbTqC7emoEHzopbqnzWEQIGzkI/1qVPKXeSvKQGJlTJxwcS
smcO4TcL52LAWEdEjLO2LV0QP+N+zk/sFPhZ2onOj2Q4X4dSIUwISNWgdXfhpYqPW0KplSxyQi3n
vKiQo8pmN1+8poV5hIVnP66ccYtqbTK90iNMR0HBJa9GsyAle80krFHeT7NV6mOmQzOsGH2b3KCs
htuQlXwY0GzndxIU/jbUtQpMqHYGv/eVL9iZPUl3Mi2rJirThBUO/1lL+iVVisOc/erf3a9mtyV+
Ho95RnLRtVhunAbAqv1PfOxgJ65TYhKPv5sOYJ70llCMEGIymcGVir73lTmbMTEMAEcNDiN6tPsw
3tzsCmPd1YcI9p+JD+OIXyt31jcwmTizmIZvPUDkQwUbkfF8TaEQnhIpGtDwcZyfadfOL3UDcehh
sM0jknE6JBuX/WM2LM4bTV9fD1oSxKYiYCL0nvS1v1RzPULmOg31r6r3AFgyK3qEtcJaJPGxVARL
Bx3YOtb9s/olxcvk9u5zJNTinV+J0dG8WLGjwWvbbj1AmaA9NauQKVgO6hVCsYYkwbn8mq+xUOVJ
RQ6EFjLGX4ryuedw9eklY8CkT6unRP2Y+i+LYFbiFR+vdMBUePeVl/f5TI8+gUzCu0p7W/TsYel4
ce0TLn/X/Uh8T09pbzd95vthoWN7GSUR1v9JzioJTpATZYVf14GFWb3GboNGdj5UqUt5B3cvhzLU
fnKYOOHW/uyMmcf58/kII76a5Gk97nR0256SIetLC94YPTteuFI/9Knwa/0zYStMlZWLwsIJ3MsJ
7MCLmVQxGl3BZOv1aG71tHeqG/gG8PaJhQOB9VJ0zZUg3kg3YWGT5HFnZa5sixiGGOT+7dzNFkLj
sjYgygDHDviQ619JFcNGXxncAynA7eog+/rLrf+V928UVczuEVjD3RPxYwWeSyYJm7rVCRU/R2Nc
aFqw0g/gvGAtZR1QauGYlHV++rBX/ATdYb53lP16GMomSOnkuUHopFGmz2U0LttUuIa5rmWkP6WC
Oeq3/lqLSAtKllDw3sL5qf5tFneEggwP8KHmNv4mv4gCMMu4+3bUlZTKkHtefPvIS+wZSrxvYOi/
UthKgR74r73cD+shxP5pUGIKD5pAqdeTI5JPCVgf6NzhuuftG4JRvt7xzb3OAh30ZSRxLK/Cp+1D
cRXj5LDPgehx2z1eAkvqiJYEsx8hPY3UhLbV
`protect end_protected
