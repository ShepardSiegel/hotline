`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gkm1VXzcryq0k1gCjFgLgw0bHiJ5667/UU15c0smLnOqY2p56TsPzYzXnMdTTf8d4sOzkR49aPsF
/jhPRIwwgA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Hb66hEZFcqnXQvs4NjvMQe7IbyRHyY6FfP0Kiai1iXGDECXhneGPHfrFSEIhk0m7LWLDq+o7F9eU
CQd6wHF1sGTmoD6FVH6BnyDnXRisLam2djN7LQIAKxdhveFvSC4OhGF7LxmeqF030z5E/GH05r1O
NNqbH+WyYaydTJyt/3Q=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YWDo5k7lWFSMp9Pv0SPj7gfJdd7sv+sLQarew3ScYELGMpgsWIKfGfyOXzjwCK1sgHES7UAlNlLd
S3z1in42BaSsvWekB8BFEi2KJ8nJMvNHPxnvPJWKgyzKrXtlccC6ilR0r7Rkz2SxQzvs3m8dpOGP
Ip9Gaz8P044lI9HMBY4msrkgeqNRbZDfRRjcpAWqYMyeSU08oYxn2y3DG3Qk0rEbKvSDh/enQ5vi
BU43pj80UwX14PO6uy8YikCcVQc9aDhRPGwD8g8RksuFr+b/eCGsv/W1MU8Kk3I+dOLOkgfYFRyB
yDcQUlAis32TVD1rMZHPxBRtAAAUryKjD21L+Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tqmp3Lreqed/VOii38eOvexqZZT8DLx7Z3WimN10X/tQV1xlINeajU6PF9uD4shSnqAvHOcZcpPr
Rl/R0t1VgCDmGeMeLbykG09ry0bPKkfXOqT2IX74Q0UNz8O43XxMmu+Ny1/0v3TRGeULdlKPhiW3
RfI7Xs4lJ4Edv5SHFvE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YQeL33el0CusZ3l0FOeTO2P31q4EZm82RwKt5pk739bSx3jDb6SQy2Mg/bkR0qeLmsvSrximGHr3
yc37TChBTViVg2EEAJgq9NZw6taJjOBye2nO6zLCgdv+lhlsGbUzzYJCEaJ2/hfHpOKGoL9PgYKx
m0B8/Lw5kCS5IEmoE2/Wo/HDu7/38fwFCmAty728mQfYJ0lqYajkGlPjK7UoPZKqVZiCmmEVgos9
KlUjkkmjtI7Dm1FutC71kPdbAsqfnmcUqfb98bTTgRNH0uuwWVK0axiHcixIgxV/MTwvYUDfMIMn
IHmUh/9ex7k7BujIyl6XZogKaRFkKEyudzK+WA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 78192)
`protect data_block
IULTl3URiXT4nekoetKzU72AgSf98k5qgADCuiFnOMHRD4EdeDPkbqNbrK7fJI826wiDRijBb1L1
TOmxkxGWBNoVRGUAuUyd+1hyEnfTdGUeEsbrbWj8XuGvgDn1jeV9IE00rZH8t9TjBask5eKnXnyb
6/ZmgXH+55QMkVRI9R0MTyL38BgkLzTio+c2SpvKaSUfwLHSzJszXh4OgaFeHdMLWKxFLpOmRi/6
Bq0/R5ZfGZp/CBjvrF1Z55Q/pGTls4aYCjf6enOpGccbVzEHrXMeHr1uEL4rvAEdkWcnWVYzj8Sx
BREHdeCghwqzP7DhMPt9Tk98AJFAxiywXhvzA+0mTghk9T/DHzNMuzvJVFgpj8fHlQEHrHeJvkOz
1R0T2/euty/Bf3FIpB2hyUaVv8ezqg+DMrc71rqMbidb37ss8f2+8rGiTZ4WIhrYwVqHGWKTuIjo
Ag6TgqlVai1RBfZ0k8egyzn/P6YhAlJnZeVtm02h6/ZVrzZRdQALctBQwhfYR3oqEEypefHggB5Y
sCDIoZZLBCgcWywkHgE28WRYimIcKOVlAr29HYAiwhvKHxOqQyZRYg24X32J+r2pBaGFge2BFVi6
Kz+leDOaqSLt/66vMxmfM9gpxPe1tGYMZk5hECzU624sXRd1PDiyy36CUFAkedb/2auvi5FljHt7
23m/hHfh6pm3Feb8j3E2QJ++YOE+8NgBT1Ayq4PIklstt7MVmkR9/npUkZr6abulXCnns63nNCuq
+AY+9OUx3DaijKVzna2E+KLpfotBZJAa5Lbf3f+8fhc1rTYMPdhbXACuPM8B/f8zvzRhFET3TPxB
3DPsQUydKUnDVsNoEbP0iHguVNTVkqkhAoUJgWnUb7i7NmiwojaPaxy0Oma/CeBzyQoz3RnB1HC/
nPZ5jUE0vLwc/R3DiVHdGltCeTmyuO5d8suJPFx4ksfPw3xFMwhY7v+GXfA4SBP3Sl/1/wKGk3g4
quuvKAuQnGXV5UcPbk/bc42WQQnPQHqw+Lcn2tOPQ+4idqIUSctlVcpnRKOtQ7JqLNYFTZCk/NFV
VGbDkk7YsP8OBbjDUzO2vr5Nt0lvYkNKX2T5RlwuN9si604zvPtsRl7P4Uc0NZU6F7JAedo7i2Hg
GOjvlTd+9EQCBDByABzUi2rx2UOFguF8xfAeigJp/1Eeq1Q31axJUUa3BmQ0LQTZxdbpgV8wPyWr
y32Ae1t8XOGBrzVBooC9WAqXWo316PClB49MGtcdKYpkA4/gd+lazSTjktY+wVwa676wEyI6B3xy
p98JCyvsl7uLxwkQerEEF3ueT3/r7oFZ1iT0Xs4J9Wd0Eo9wN8c1hbG76rP/7HLvKxcqvth+C+mU
0QCp9HUoi0L3j4u0XLqzHNpQ7umr8WU6OIoNeJChWxHDmJ80HMXLc4OE1+VlSCMNLJ7h3ije3Hd1
Fj+wbQ2gkhvFCes0m/aB3tGqxLmT7Ge9DZokQ0swIwyeb3CbbwAeEXnk2vk0NdopNrUTUexTH+Am
w7yNqaktfYgrZXdp62tx15fefSH/NjQXshrDCKVM3RpNnL/5K4YXrzUwiBDQD9eAKAU7qArr8ZIS
xuSUDFDCeTjoEZfB2cj92tvy2ICh1NZF4NOxd9UPqZ+88uHI6PzApG6Zpt06IcMnb0WJtFS3GS89
+e3zn/EUtHULdoHSnekxH24nBcqjRu/tJU8y48mw92R8Hm0zPJd0t54bKqkU+AB+9x+Q5dFBteub
bVTwLqAFTSD+01nbUgzcwaIjQfoSyKwuNo4MOUyIYuQyUxXYF9Dz6Cl2ICH9Y1tH31Ssi2XUdloF
GyQJFE/8Ohw9nujzwGLXPcuihaOk5qyzBXOSJUy6Ba0eNI1lbKixFXIecOho6oxCu5tGU3haw5H9
eCg/RKZKegLymRjnpkfCMRQ53KAH3IF6xr5fZKLtGkgMZjVuBY4f9q1+y5MxpMgVf2mV0M/wzg8R
OORfZdAxqyw6BSnT5MvFYdU3AYCMQkWM91/saIjI7U88HKb7F79UB1Ko6+gr2oZuj2USBnorKSu9
/EIidxFxPBNb3BKK9uS+7gfEgB3sLBcaScdX6ZAtCqc7L6EAcSzHDii+pxfY3W3+4TrK6tHpKFRk
f4c68orGkFmRDoBt+P4WV1BkYfBtkcisDHwF/4xH5CHi4v3mQvMFS17VMKhcYNKb2mfgZhkdrAdH
YwYpWbIjp2u16gG0oLs8164Q85Uwcv7VJw5h33+AXLByUGG7L37/CfljzGKUTEq8EFYRh/cADymj
WGXv8F74Tue7KVSimFr1hARrPN3dgEf291vezKPlqmgrC3XqNn0i8Hx8HBYldC8CpDsgwwleqkui
/Qy65sSLhgbJNEq7RiVtnrdDlLfZCxFpYZUOhvhbor75b3MR37irgfWa2wtwnTBX5TOz/QAS5bLp
HnKv1y/DHnQOyY3R6Usv5Dwte6vkQszfVjEzhNnkm4n1ZAR6WpBVXKQlRwmbIxf7TmuodNUxHwpY
+VNyAB8fxvCPcBojfo36U+/uRQnIjfFvhegaPi3V0SYaN89MSZVwmqp3VfS6ANXei9LZ1DrRgSP7
1m0y/u/lYRLcNzMWph0e79NfB2Mq1ttFtugQQv9u8pH73/4hvuznEnFMtN2yvrB477+QNA//rYPH
VKFCCu3AG5gjQEg0sgELxbzP9IG/F7mXo+gSXCTbyRQsBhcteXEXQVQeXXPGCCFfj4Xey/iJ1ver
EQ+qLdKMXzUSa5m6N/Nw0DoiU02xXpq5ktaO4ruZfd17rR3bA8af7gS2z5xGP6Il/d6Sohm/K0UM
uOknWAmKdwmISWFulrPwu708GScxQ0jVJH7mEAL2CQPRZmfVsnjIRNMz5g6bOXnv9Vq8y4UeQqRB
qlHGfzsczEG7vVXGVksUhr8byNJ0ck+a/eV87PS+tpbKuMq5ZTKNbMMcnTAxIviKEnz/T4V11nLN
ioA3Xsw0upXuhlYcR6/5rU/FWgT3KDJGOXKtIwKmYoGOjQQiNqLiwRi/rePXsVhSt+k8IUmjLm0c
KTo4ozyHQeb43SC4ErBuGvfXBpzKY3XNDmE5cVvFs/5EoJrcsWFGmxIeKyG+fasJNaKk5NVfXEPz
l84pBd9HD0ZhGt+eW9GnOfU4PgAkPHukmPsLp7uUcf41BqGjwqjSZ7YAGgT4dAcmzow/ZHCxPMZT
KWiD7en7QUtd1KxD+6JCJhbI2kfN4B5ssgvcvyuaHzfTL7BgyMf5kmr8kgaU+YYpuT7RqgAZ6TWK
3YJ2xeOYP4kO5PzdPVto2pPDx9HDXOBRYT6zXKoqYxCSrL76xFr8OQ9yjDspaPB0e57U0BOJiuDu
ZdahhWJ/UzzdsLVDDw+WFD5toBlHvrKlYehmA+NDnCA+CQL5FNeVDwW7V8WrzvdHy/AJNh0vIYux
xO0hcMlpAeLU1bpJQv7P1UuYBID7IeX/efzaBGSDXUPr2zuJECa/eCyr+jbq6fMxbL+hbrQUS8bZ
+kFXrvylAUGJu20IAzoVkot4hPw0tCLccKE3+RkrV7Z6/kpeIdSUcJcMR8864fcUfoL0/QUNi8dp
3CnsjlyAqyE6bPdhSepth9qc5ncZLZuEH+kwfKrdKNOnaATuKABX/6hLWVieiCGQhOM+/wNZV7Vn
cqg6v3HB4lBKc8hyIAd6N0L4jZCn6d7umPWcZMxZXhOnXECRaUV9LzxkBlaf6TCnVkR7ndwVfvzY
C8+q6JrVLyjXrs4ECbnBPtrEpgMmDpyPQrp6keyAAGJ5mmkWVYfYL5SRErg9onHtuKbE23+ed/kR
6us5oZm6RWyoItjUNYUKOCcENSRSlaRzz92Z970FgH74Ct/TkCtYJIMTm/lpf7mNga9aQ/hc8nrN
6U05vs8oIgMhmVJtzXof3PjYIRJtz4bssL3gGD6cYx6lV6ALmWeyxP/pLXLA3FLrUR/wg8DTeyTk
CzC2/cfvtKe00SGPnszWE9gb6/9a2quAaDkdPd24dx7c0/lKg+B6vBAmAQXcgnmsmE7JF5M49FAz
3HSE4yw6+0jK0o2MYFh1LoiWc49lcV9lKEQiX8iU7iOWBGRiQq5XXDNhaNMO/FggWmXhxaF/WaiV
/qrKZU6WmWKxotVd2/2q64Vcikd+m5PY2mhjjj9JfMSalckgOYuGU8QmH2UQpTA2PjHNZQjI847n
ztjqbPZyFwaVnMg0YfCxrWfDG7w018wN5wGr+/t0UbqZeg0jQcfUkjAmSjcfh7hbSL7cmm3GeITN
WLrT7NUij7FdUQpwvv+S2Nf34snSoplcv48JQssJzdqvGqsJvMiUQEc36kIgn1tXE97dh6Aiqq2h
9mmnL3+q6jAHqHfkdxRY3ms6Gq9g6JHwSOGubneTxZa1v4tbn2UpT+zITPlKQNifrYvSL3BNZZOn
BG7v5T7HQBWv0W59RjzamOeRI7VBgRG6zREN6aAvR8N62uja6tBaYf/cr2LwJjrGa+RoUrNOIlA/
uOOVs0EuhQjmJq0kmpZj1kF/15Y8sm6cT7VLW2hsZkO3Tu3OSDAYyOP2pofzUjbI5MultqDPnBC0
XupRbZgi9Of7PI9W7Kb+uq9WWzQ/iHGdqyfsrciVDKYLQz4cOX3ITTHeMGvZ+POEn/kF+WI6Shxh
wxS/kKRVRjqV9ByzHO0wo7xSbmjt0O2eVD0XZhgU2zsvSEFNUOYddD7iPTGS9lSSDGxKHLSvAYvw
oMwQsVOXhU1XcGHXD8D1l2ULK7oXnGbeWWQqU8tsgxlEXEoBtoKF+d1fICem4Mu0SegB7PK3bVTP
y4n/EWQ7r0rBeIJc2xrfjH71W/YcIhG7Zn0xEYbcrWhZW38ZYlXHvttNmL/HQRYpDdHU8/L7/Sbu
yH9LG74v7XgzeFBVewgo9ne0VDDmRfwnb/vqgLQxTUpOmAFSETxqCAd6yjbnJSmrJ0XMP67yOOMS
99ENystG4eAOf4V601UdNxI3tpVsRRXUblXRcHumKF1KOBixXtqVax0PMiPkKue+LvIMsO1CYQ3G
h1xUvEqxG7O+jcpL5mUnV0SuidrMpSAJo7UB6xkiiNdia6y3nHVuHOFrotje+bPELWWk43I+JJJw
tvbuqifcxvMlwm8vutI8CTNjdi43GCUQBVB5TFYHvO+GP94SpbjKbtKsSvYtD/LN6mlzVCsaT6r/
gCaoM4Ie6ydYUzwi+Ih5J2//D1RzP/uMIE5TTwKGxPMyx8YhB7O1QSthkkgdey/0uIC/t53n1HvF
Wqqv1oeeOJncj9yel4tI9cs8P5yBNDfU8C5oZ7r6YllxrUgnNt9kuXWBl+UpH52IShmKy214KOMF
FqYLXwtOiXpL7TxD2b23n+3G2YpFx2kUk31MXyuN1q1N+PtcGgg92DHnKoVPPpAS6D7JRysSGdEB
lwJpwYPiQlthdmmGY8g/OlVcR5/qhWA4b2R6cKp+jdkIU/LC3I2XZz6/qs8T+RGWswFqB7PKQQTP
jTG4saeuJdhELA4k7q2jEho6cAXzipvD/9KsIn2PUip+WV4O8tiQ69g3i0yin1UetdoUEbkmjDmQ
QpZe82MwNQnbEIH5u9Yag8obpsCq1/tbubUFQ3q+uVayay6kX+HSRlNz2JnX+YgpPZVcslJObc5l
7t/8A3vJmKM4FDFsEmE2cCrq6ccoa70KRUP3lhMloHOdSQFKH2wG42JMScJzPbLip3MJOFe3kGUC
4AkDzzE+LKBhZ/ZThbAGjoRFMPr9VCH28nCAQS2NOVGPbHVDcnir9cz5eQfepT5J9WL3Z3yTHzXt
yAFDJdTyda6MiiosCGau2PYoRJFF5X3NjpD42O9Irjv3mt61jr2kwSteyBlFi8HdT24f/Z2B6fjL
9mRSzX7SyLhjPcj4ctAPKR6BBmg4QXpTf946WmfNx7BWNWYRV1ZmKB0xDHMiF3q4/ypCEpbtY+y0
muu37xY6JbeggZcMwVC0FyTP4K1Oq2YTYbJtu/64jN0zgIkltEr7qSmLzHvlYKKMu2AsnQkQu55v
g5G9SgYlfbrDze5bxYFWG4G0mUWl2rrf3KQ4x/WtXDyGm05aCsa2lblvnG65OXqyXhApzZHs5dvB
POxt/fEqvFjvcKbLWLLoAYuDQNoRxgkqHQ3P8Lv4sd4Cuor8YbcGF2SpsWaBBffU2lbXYKhpvysN
018Im386xnQEpyJJc0okeDCCMgY+ZUrhDND+y6T0TduF0T3HhDUVdRsJgfOirRlsMEOjG18Abqq7
+kVxEBI/259iOa4kJLwcmW4pJnNDp25cqpQmVngtJjWmexa3PwGChnRkE+lew3+sLpwtuZx8MOGh
rTbncxkL84EdEtcbtPSiXQoDywRFqqfXCyGJ/fIFM8zWql69BJIamBUy14gyFoDOeB3ZV5CC5CUd
81Omb7rEs1RiMNKig4dty8Drgoe8kUjylwx9M9kRHSrVA673TSwryr57WeBz1AYcWfZqx6t60iU7
RDtz6oRQ9lx6PTlwPY9DphRe+L9UccLGIpLpeMtw9h4LsOEwuZ6wGfjdNxPA35bAQjIPf0dWJssm
Thvxbti6QGEcbOW+pE+BxCMdotKlQfX2tQs6T1umoM9rWJPlGbklA5hjZgrmkclBlDJ+qj/fpbW6
NFxbn86q8zSUWwtjTUV8b9bq9xAMK1oRMTC3NBMBnLHV7RdnIz5FVmh5IfDjfEjdjizKDLjmwOgU
DvhNXYycM114zNAIwi1lo9Bl8U+xsd/klKhjPh4w2P1ibehvW541EC/py3LSSBYSO4R3C/BxdJM2
kL9zw8tlo8F2HBMQAdM/vVYQllEM4Zm6uLQZb41jS139INm/oFdSnFE8isk+L56ohrInadX+G5p0
jhrIkiCDwsQ2z26POHOD6o1ANl1FxxtPPI+2roO85rubMzbSsaU3Ev3HR4EWSfE7AiJi+h1MxbWw
WsyDEd2cfubT4RDJ5gwQi8rN5/X2HaI4dHqQsWCJ4Aub336tmSAB5GFT+Gu5YAW5c1eBkiWQ8jsb
c+r4VoHMBm15uF6QCq25bFj3N8yCTodT/Hbn4EopbaAwqzG8umxSVhyl35wEJ8LblGyGZgRAfj8u
bf42pqrO4WWiVxg8LR0yD+IhI8Js/3MpeOXD3V6lJ1IGXqluZj2xVGnPQ2pWiclpfh9cSaJXxp1i
9iPEg2hWuOvTl2DkA1/hgVDTYtYnJ8lM1q6YB2teJeWRRHWRP6Qk0ii4/TN7vyNpa8phrn6jUrXT
fqIazQFbfxxlZqPLzlIaTEdbwDZJs3z+N+qOlLDtUixEt/S3G0owNu9sCvZdrcPDUmKyn2NHP/t9
dwcRYxkmhBF9ZC3LZNTUTAXipMBNEB+/f31fxyUXBOdj6uo0sn+2Xnosy/pAluan5o0jYcG1uivB
MPo9GRXdyigpyBRVROE4DTo3JEkPTbDUwuzX1TXOzUdWrLASXpG3yoZaF2xxsVAdi/I/BWtGAIV5
ANU0z9sJAv1SJMh4BbsrTCQZX13NrxXEG3A3Bawwn0fve/GeCjMeAWTE8ZpLKEF/eUBz4zRQVRnX
oU/mgrutZixK3/m4SFDVFNC3NY0/wXL+w7uE7sNz1qb+R+BUrhE6/2aABIrB7zJeNY+KxwMqE40c
5AENU4ml1eHfTbai9Q1nTJ5nbsMNvzTr5Z1FHdYYK9pGke5Bis11HLx6z20w5u20A7W+RAzSlmcM
H3flsVfytv085I2qJ2tMD16rBMFo1kXzOcCdMzGZsutLrENs4w6wxrtfWOhrU6egyIInXUlUtwGg
X0oDLvFagiZovHhCAsJtTuD47/czNPfMDiIMn8tR5B73EOwzbVYvkWxy0QHs8Cru32mR9Tw511dV
4IyW6wx7SaoekXwPB4UFiFyRwpHRkwUNTHWEOMabmiDpOPZqS5/vwi5bwmCuzNF84qiC/+0p0pYU
JDwO7sen9HMZs7Jq/+XFfXYn8YuRKqqPeousZo1dtju18+alKwArlRbrWY5AYjkGMyGto+pGf3Z5
07M3u+7my3kgBu97ktHlT4wHBtyWUNEqfC0nXzLGj4faWoAbHZe59U0EOqzXhPzkWQOh0smL6CmK
Vi2CPy5w1ZkWIaAS+SykFThcyYspW/pbLQscSZt6Ql0y5Tyln2cCEGIFQUZqk4smkEY1uODGEFYt
pHaBJOQYGHLAiRbn8+4ONwtK+2ePfHaZIb89gxWivAf9Q4MQVfDI7wo9Y6DQ07yvbRxo38pq+Y91
zH8uy3Y9BZDkI3OIggDss/VUJufj8VoGbYqamLWz99h2AVMyDNElQsXIXck25octT3Mx9Gch60Ld
cyDB4zDeJrxm7+AnMg7xgYvj/jMe68JdN0OKOI6oTAkkID3zEX/x6ErA/cjWooGuEv2RdASRyTV5
YXLuzlr90bmE4yaG7EcZwr0/U7MbtLIgsOfZSmV+RH5HcyCdahxcAQHrJS/6CE/5oSbPCZ+JhvuK
0L4axxctUhQxF6AXN9B7tiwXeyMTvsXJyHr5vbEyPLdkVMkJW4uGBIDn8dKs0RDuVyQAsbb34HPD
6G60+5XSlBvs7KgbpCBlM1965IjBGBN22C7/2i+sHZA2Y6Ap10/9qb7r20A1V3nJoXnLVz3NlIFp
cA3Y2NLRsgdOhE3LqOfcl7CDAc6t6abNYoEKSW8qG3tuiCeN3Nxp46hxD/WIahcXmqw8RHTHajTx
JfMVJsHJZqdktC6m1mJQFEx5Lq9LTEsn1a+JtMCC4aE+tjA3txctdFCTm7a8fALm3XQ7fdI5otiz
9GOGcaC25vIDGl2sNRoFNEKXzdyeXZ6LqN46loVTwkaMCqT7KmUuxPmPqLWXxc/5x9yO+jR2ubFL
e1vJmTBU5mXZW0HTdQXrjtZcyK9eikvHRdemHZr3CmYKEuSfQC420v6R7cPbvfpU6DisXswaE9KC
vVPr49jb9cQAP8dBH4gYKJDU43NkAdv6ivxoRzObINWcoI9FXPbT0LCXA/NB5YjBcw9BSy85X14Y
BEvrtqV0j1foxh5/SM241yulMkLdVJz04kTtBepbpXvDSO8O8ojl5jPIz4TqlyX0+lYvZ4AXXDvV
KLgkisc0gmnCUExgJQiuMfKtJ9rN5DTbJZQjUaPZr88wbROIab6GtcYTMagx7qK9n016UeMEfk54
Jr83GQQoSg11Wb+jbtO7l9Cnn4hK8skPvHPv0NIlua4IzxryiOC3FFqefICe2JGAMH7WFSluENww
2s5tW2fvxeFlwNjlbmvbricEsTtpRL41zBS+R3GlRIchtUTOcYijA/ImfpTzE4XJC7XaKRplxWUv
Vn110rBTfv/9yYVPcQTeuIMqIMxPzh2pkWeajKphFfICSgCoAKel164UdzPf8aIpeQRby2mPrZxt
0uaSx7bvgMTEWDXNDZpFBAPQ4FaPUAptRYkNxIAUl0HyZMP/PUFEsT9CwxwUsVFq7X3teO8Tw08U
Ltm+7gjMmWOpz5Ag65zBRQPEFDB2Rd2I5uoqXAKQwzZZPXv8zzrTC4Ppket8bi4q5LxSLwbrIc/h
pyT8CKE0UDWIIvfZAz+DPo4KeMW1g8PTFgw+AeHz05A1XKPQvEyFAYBivhI8Ba/sZ0AnNe7sN9sj
qkEAeBEazDzggkPOiEFgduiqxa4TqLL3TUVC/7pzRvo9s6WIzgJgkxv3aXDPEH2rndslrAkusj89
P+jL0Zj+i/c+0Hf1dMjamYgxDod5eMsmCWdAMD5Uo+9/WXGmEiFEpqJ5wIiG5fJ9dW+iJ5EEeWnM
eEkYcnZ+ChaSz9S6bqwiQ4VWFKToNG1jluCC5NGjhpEuOEBjOPWsKe7/NH7l+F53jZC4mWkuxdn8
vmKScNAM9rP/EUMapywezMETuyLMgRybdTJzGOGr0DHrGYHvLifDBZD8827kCCAVZVlVDyvYGss6
BGCDddmbqfdQ9wmt1BPEnBTRhhhp8D1OuR6QGgr4hC1ujpQZ38YE+2jyhNY/X3dizlvskqF2wOuF
feRBdFBrLFcGSCOWMx3ev2KYUQtPW9KGW75lz4ggCMbN8C6vu3hNjP1Rl59V2tTsBnZkttpN3rPQ
SwT10G1+zWmVzxsVSEjcHXmb+CNDDksBVk0yUqu3NUKYBk85+ngAF4SyA2ZtcHkZGnB7Fq+iRddR
wc2q9wgFE7pFhZf6qaj8V0f8l9YgO6pj3exPLHWALXFBHZyi5kFjh9u/ANNEs2NFFu6kplfHFX34
7OHSHM7Hi+nOfOM+CG9K+7pvaXk0SNI2HpfktER0amppvy1WlCbZQiZwbtVLKl47xJLpskJ4uJBY
Rqc5L+VmWirrIkoNZoAzVauHi15tT6SXSMspjq1auJm+xiBMqqCFceDuvfTO0hf28n72TfUPMP2n
wmp3+lVwlPVmpF0q4DoncWlqMBMGCwK3It4T7HimKvGpyJcYf5dytC0dDewl8hc3dXKXmQo2BnQZ
sHdoLgyIYlhFqT0bojAj/3zM12tOFa+H4qN5EOWGxC7x/pYVfVE3VcKhEMmvMEs0H49256fkAPWj
hv9pWYE19vBQ6RFXtkdgFr2AqJiVOKIglWNMExgJLosc8TCQABfB3Pc3eQ5ReZPWXiHzj+Bb3wF6
Sh+mSJ1MVBShDIZ5c9mvSkhpk+0n6WOexzc1fQEXNgibXUwS3/CaSLxYZ7k/3p+biN1s35dzS9Iv
byGsV2kXGqTAfT0MnaieAtou9Chf0TySSNLgUHvIpDgUZLJQwM+AUg4tM0C2ZDq79hMkFiJ9+YqK
BYsDm1MmZ16MTFBsDw5LlmEQSVCVfBrcdgoB6mkDIh/FuUtZvkR159xJ1jVBuc/WHuxsr/TTvHuc
rlPGo+zy1Z/4OfPs8gAjn/EV3XqyCwfXq/stbk1c6hAPVv85+6ZXXVKMj9gAIVM4MZ/SnF17neaP
KL5cJEZKkakCZXf6DKyrlKOU80sFSpbEtiSqNfx6ItIXBso8cL6BT2lB2T5YPiIhNrXCn6VzSAqm
zwjlXPWaX+3Mp4blNZ/0XCg3slpD97/m9rQxyEzG3NnnHV4kejkuKsT0axCJHstvKNp9Chaelsue
ngwhnk+FJZbVXvluAdl3dblf+IrV6uRhYstqnOzUi/6wkJ00Nr1pHzQ0SvqVyVAywbTtWDa+CLp0
f8wXHJg9qeJgV1/q3n10TVWFJzmvJ6bo5clpWEHJkOpvx2uEVPOZdokz2hYedwumUOArJWhgkInd
KFu5THq5GOtDNo4NilaMu/KYEL1RDvdoXXrugDvPAoFGhwXRhPlGjgjXViEW5KiZhWIcDfkMLB3o
MZSKQGIJ9E3rGabjx2mEzvZGJ5VQenIFWSJIQtL3vLslmfbCgc1+7Mi0tsUj36B1eBBopgXZd3zz
KW++29WcutCFMfTWAmM1ebVH4FpeMTRNMMKmfsMzKEEewOmO5oZX1OyRtqpmAOx7+I0/4VBxDYRa
MVH66ZqLcGlJRIVwO8JMlU6k1XNMPSDjbxh/vffML+R9BbpA8Cw4IBV8yQGPJM54D0NlvCNSm05z
vcDNjw7ZOD/RC6998aHFyHnWwUrjnGR4YiyWqOsGFEvf0BrFvJo+F8Ci2QJDFMj+BAf5Ji72z6ao
M2P7Sibb0ziYME+FW61t1q+zljdB2mQocFkJ2YC28tFG51C28XWxT4J3MckzW3ZRkcxubaxGXQ8O
BRNzcihDnoO8ltiKV6ntMKW1cTxbAXXEHw96ITeNVs/W/aNIRJ4TeMgFL9IrCKbqDhi7FntEnpMj
jHKEsAmJ9YB/3yZvkQNr15ZYtzdI9wW+QygQkzK5i6+bzt6zBePD5c2BJXEZ4ImLTrcUZXKap8AB
5gtkfwx2ZfAtl+7Al25T43zv2R2WTcYTadPLSlScPno6lnNKAo9/0IvuBKrs+0JdVTlCJcUkXI9/
ah3KGaEe4ZyZ4B140M/8j2pdQyPbk5ppJ61OSY5erWrgFAeWoP8bxx0HGbC1dvtOQnEJRORcExcY
FO1z2Xm1hwnfGBiu5I7nE1u58vmixbWeKjSgLUg1U4+tC+OaQbHSPNoC6uTb7imuhocybgMJtDYW
hI814Orp5wtbM0xpIb3IAHymDlXZFTmUCk27Sgg5/K4RcXbVmOy4UYuj1angZL/RZrsnN8KcBD62
satkr9QQb/u12rOHiT+/R86KXB/z/02CikXlMvJvD/nT1YEA3Gv43fOOdj5jpDndKHeJy6hGSxCX
DTphpprUN/hmZ4lKu2wkX4BxSfRpTxN831/QbR1Zv6JPx5uaWsBgOovcBkqjPQbZ/UR6wK8zxIU6
GiHNzbeBcydNiEcHuUm86IWGnzWC4qWPwi6JLlCfmE/Uyfu9iYFml9qMtlp2x57DtieJqOk4VzUl
tUr52HCx0GwPoWOa8wNxNOpU+zmtfW2hvLRHbB2HnegTqk/rQMABqAEafiroDNH8UV1lfJIIDnts
EbexxG+VeE4aD+M68ZzRjVB3My6UMpFJ2jZhp+tVUmJyjuPNNkhgI+kKdrCgXxV0p3eASRMiO3RA
ADO75yZFcrNNlLeL8Nwh+1Db9ZL+P9QtMfCH3CT2/eRCMWznQx/6sMewXG48xNhbEsPpnj7aY86I
nbgov6i2e/FdB7i8Oojd5ogI3RwHE6LMWXFcsb0NC8MfTDa3iL39WB+a4jmoAZhFV6zKZhVDFR4r
rHiAhZE+KM81gk6U7xxS96f9G9nPITe7LBeF3KNd4u4aRYkvgex9sGHJJk728izjldIReZyXQdov
B1e4d+CuCxzFdiSRx7hMSG2kHStBHtmv/JYZAUDy2r0+ba8tpV08Bf0Y3cYb68gQ2Zet0+S9g9AE
e69BKk0zJCi5belZW1eiTPQFKpJgtJuBFX3Vv65JSgRVefHfmiCnzTvh4+jOuOGdtztPNETJLI4n
a/Q4lzbeHzaLR0YTN9m3x/L6KNsVE/ZJ5HtXyCXj27xghChHSFEv6VnHPzONTyB+GCz0fqxUF4vB
5sYfPp+MQNyzBVs2pCoRcVP3SB6WuGO7p96ygH3OLbQnDC24sKZHtWqOjACDZB0lseeMamD1bvhp
ebKHwYfEnyihT5l7+wqqExMdG/SE2jm0KIzJdXEj4wY4p6BKmKCXmX9F4mirdu49YGf03mzVTL4V
9VdaRqdo5A6Ip3LP2zM2h90TS8Nm3UpMQf9vE3EzAu2VtwWuOYJfGt3QAFctO9Ndvx0yEpuhMEWw
bMqiAfbagc2LGU9XwpT32HIewd64ihcuqf8wm+x0874hOp3K8ekP2RxbLVf1yJd3hF4eGx08+9DF
Z5Sr6J+RUy1zhU2qFqDxPDytFhajuPejbGAwUikK/SOoiO0koSndSkYd3egSASdCqPP3e3H4zLkl
u5irY30zXbAZ/8HnguegR/PIKiJim2/6gtAsIGLfyQmuUMa8DnxNvpIaGCdPXnZ6FdvthOZ0o5eL
BBO7Y1iMPhF9fWi6Xjj0X6Ed+i7hrGhDbOa1DvvsWrPRL0n5JROzLpi0CMN1jx0nnYehdxEG3UAb
Jy3kFv+aIzs+6q8QrhD+bAAaMhcXUKSBdDjYdMpJ8y379TPJX2ObXem5naTVrI9L4SqhlWFoJOGC
6m09JVkJxEKpkpwM69Gw0agmzuQI1JBo6AltVgKsFKclPw/knWYVZdDL7Ug4YxiqR/Hi+FYe533B
JFiYZ5YmaEOTJ+KACpTx2aaHxGU+e+wXG/PiqY/GPxMoyUtwdXigdVj5QYMUss6gR1hr4oBQt/yh
QponIvKA/V1MRNyERtOM0+QRlYJ9pft5WdrBlylHgPqSAZia6WDCWFRiLQl+w6h9qfsqcHE/EgGd
hmTsl2fgM9KCAqzFwyhQFGmuhmZQzff182tZxD8P+aFio8yqcgUUV0Ph4R6uMUF9q//4JW3Fq2Ec
R7reUVYCkL3W0SXpvxWCOgqodqR1X/HO6KWJu9BhC2EOyfig2cBQfMRzrzufnRb2e1XqpUKWs1Sw
juXYr3n/gsbJ8asRTwZ1onBy6BjKBW/oeFW8Tkv1qgcJiV5l279gcLjLVDGID4aJxdt+TuwMRsPH
nJLAJg8QNVRsuVmzWLJjJ8v6Fm+cJJaJHuOK6DVrza4bZQFluPIREDo36gtI0CZF8REc/gEA7Box
fnTl6xU5uyhMeMV7NvLn33tvo8ny3Gt+PplessS9vSMadxI4BHXV1pbGYBhWwdnXznpu6eUDJVTy
Eobo3tTUL2SQIDd41EYvCFFi49Nw3/r+uPH3u+7CxzSv9XVdjSGNbhGGNKyzRBpyhXBj6IKjKr74
dVdRA4/zNkGrqhLeIrl64CvRjl6lRbvOUw9d9eH4f69YW/BdYH6KATzWcdUW5lCcxTFJ5E1JOlQ3
t0CR6tdTsmxEG8+reYZPIJc4m+LMAS1Tsga7mB+vbhW7xkRf9/I0TiL/mt7LWL0J/alX6T2hnpKC
3Hvz3Ao6U1UVkn7BxGA9TgqAhiojKvallnVFxQ8HbQERj552nsYz9fibvN+uvI91dIpblbCshIPu
VAUxhH0J50YSR5JiNYb2kb2ABK5PC4IOLR/Fg6XQNMYGahmwwjHb4ATaJAxXaSLxyTdnWg0HIquL
mbf5aVFlK1rKXhMQjmBkvViFeue8wOElt0Q/1riqveauU9YFoqlxIceL+C8tPFgY6EtuUqZLLlNT
K79N3DunW9oL7ons9hPoaH/f+apGpfF4lcOJnmu/9DEVWFfOlaCDgDW5QtxYNAkdoWn6q4QK6RpR
r8BiW20J+ToeIOmIjS82MmAGoncWoFJuHRXO/r6VgxApbjVsMeEaHZVsACvXQ7f0fYOB1EtYjqPR
mOJkvrKOqKvG0Nm3m39wRH2d+e5LnvJRDYBlkRuGtUBRaigmqkRjHkdGLTwRYxl//RvAZDfExAkT
Nyh7e/Z0/HBs2ujQ+6ph751LXm4K+fziIJhShK0vTB/TCNDMtaGH3J+VNA6pLzhFpGzdjM//NPeK
TK0BqxNUAuQ4A2pIcsisQdybMPJUn/WuGREC2mRWZbOBXJEFIHShK4bWWngErQu8Vxpm8/VR5jUS
YfqNkT8JSY2olhxw6w6ZTFOPxXPGVVqG6m9/IgvHDiV6+57tDwr8Vlgscktdyk8ZSCEiSiWujK4g
w3v0yXvvRAM8SFUui5Bb1xoXd2ntvI6BG4BejWG6oeI3Cq2/E9e09PJQefUEYtHom4nmmqwlnORd
Ko+aT+5PXdzMJ5rg8OVI8M0PyCFooy98p4rL9ahXEO+3E7ErBaU/6WmLMdaMBPo1oTS9z+UVkU2y
Z/qIOOK91vRpI0gWll8iH/2yLzz/JQQsbtGi+skh2kDzO3ng63/xo6rS17F/rf80ite11vtzH8/K
sY++xCjP6F5vwCxTt7fPebtcg37wwm5Fek68Sl7UzAIG7H7OiZniEWEehFkWqNttFHhVTGQV2f8Q
+6bbwz36EtzXIJdCiinu/D9wAuxKv9sPNV7/7+9HhqZ+KI+PJkoTXNZgJLpROmqcDP7BA286SIfc
/gW/SJShiiPjhNidXuQ/XXVeMtTOGIknMrFzsXmHBIoSfJiR/wgx5wygs6z+70aQxCkw8CDTYrcD
jkQQqIgAaRF2LLyIkJBsfswVk/BK5I8hJMrIqG6GVCRvolg0yuZ9k/BxjP4AllrI0gqyKG9mcJwI
FbmWs50fThL1O2GDlF1xarpXqg2h2cIQUP2WqPGKhoyulNA18o4q2Es4F54xcEWMAqCmEAxjkZON
mRbN/ML991neVCnKzAbllAwqIdTYd7rM90y4B0bQkl0Dog/3RcPSn8BlTWMPk07aUuy1vuEhNwQ0
jqzZf2wEWzUd4n4wfZqxTRN8cWXo8Am9/uqp9uzVkMmKzgFmCI8aOAbpLfQ3duantJmBea3v71gV
J+dpghFvp7GkOirY+Z0V52jHNaXcongvRmJ7KMGZFDoRNP0Gi3r3ELuj/OSIrnE8BF/mNmuwXlmo
+dA7Ix07mwqZSMLFIWca2sFWqURveCAsz+bi3EmBDAQQniE6aL8H38IoIO9wllCdYZicWr7IYZku
ojPhOtNE5Aq6d3L7c4mJA7IylcYa5mXOTRiHYhjdWTcGnCZIjFLCe5SOtP8SEqvOPNJ7q4IcNTC1
K9mYj5Noods9qqc314ykdjTf7181WL5duCOBkjtMvI4PcE7/2FoVChJ0Z+jS9bAn7IFmMfZPxq1P
ptl4lfy89mPhFowQ8D8iQ6QqMoD3LlRRZvVxxaS9WqBtCI+VVdzip1Q2xqgwVubDKznzhKC9pav2
OFPsJGRsDBQlMKMOhPkT6IkiZePrJw4M7zX8EY1b8TAI/viphJtSWj+DX544FR0oH7g0q23syBst
LxLRcN1gZCVeB1U1Ep147fvRySoARag8P/eYsnJCllTwyoA1NzoPQtV2s95ARRtdQiSVbWOj8zKm
ell8AtlG+OrBW4tR67nLwetEp90XcuW9TN29H3BlOPKeNWmx+4XpWlRhgJAk9d//fCz+65dvIgKi
D0vmCiCRfPydlNz7JXEuuiGimYG2sdEVdgNeWQXDZQAiu1Yiuj+mckhLuOdTcYYGctJlKyaA+FkP
/JO6x2zlqGOZMECOE1j/V9DYI7HqeToyMekcxDeBUA8Ay0yzpErvONrLBDXb6t+zhRzKsCcMEi/b
fXgGAzEWJ5457u+ZviRVI7bmSD52vTLPVNHLR6cr5CyryzcrWDh+40D4gYFfSOW4H24X5BblYsSL
Z72zd9mg0VcqZooJlQHrdZ/zNelVw1fcZTfxutW0k0lnuR2Z3K8O+yvN8pch/jx83AvmgBCVlJly
Ey0PaKYk0cSawxp8cGuRtuInQpHd6B/D50UqEnEgjbvitFZDQWR8I+Qr0wyglmwgL6M/8CVNgymK
Q08GMRmF/NTskN1PB/Ksyf9EEkHTNO0FWAyxpn68Ahj0FNMmmKZRg8RSAn8F9+K0v2XcEy8ndypP
KjKHtbPRQBeApgt3Vz9eBLmyqfVFYwBBYK/lTwdUfGNCAVp6LbtwN8GdwOd7aluVcmygRh7shI9Z
dCmqdrbi+8HkrOWcQQDGXig3uaI4datWhUIXJMIZYVZpMQOkQKAg2Rpkw16jWyfOGbHvnDfmFcAF
+Mh03zOPFho/V1WzkXKavsi+/I+X/hE+t8+vPiaxqTCkEEY/koG9NZpO+Ch3z7hxcWa4ClXa49Nx
pR4iggrzcFPZTJ5uEdzJB/kkER+wYjh7kCU4fug//EtI3Hu+YEFlrCcp03zouroMUzTp0WtQJcmp
pFprLAeC6njTkyBGpMCdSHWrJr/e+3GBgRieeG/56Mt8BA3a4BMmB1R6s2i3OVgdMsIisrpKk1aN
DNnuLPrYjTU3TtAMK/LCrHqmBj/wvLJydViCrsLYGhnzo6moCrf1f8bFkmu6IvO+8HmJ8p7Hf4Gz
Hc81xbwr9hjs+aXYtfv8z/4iMv7oLQaEN69cfIZlNvvdpjN/b2VY+l0KGk+6KGiCTsKfLxFfRw48
Ox7zZtJMLM/r+gd2VMKhylq4tBLvtLDijczKb9jWQeMbAJUTMdSV8W+yfiwfRl0PXrRP/jkEPoaP
j9i/UcJ9y+7X8lQwByPGdf6p7M4tzLtPt5p3Tcj64o2zo3NGJk881TChtkjZIAZt0Sav5qLdDVnA
tgFi1sV1JmTBB/cHG7vwkiZ/jtYxDHv9yOx8+/VBSyrd1yCo5nI9671/tEZ+3qjeDON6zAZ6kNP+
WldFG5YDE/ZL7Ev9jtb6OcMSEVScK0LVxqE1shAB5ueCXMY0dSP63b3Xj3JLJguU6UubbVqYgOro
H6YzeD/BQyEic+Atk+lZKDufRhjNo40X+kCOpbv6C0bTd+wCKz4rqcRV6Jra3WqP1FyUhLvEVKXu
svItLYUe9g+j4VYfrhv3yb3giKYEjTHTiAVlGWnUexKT47fC10ZP5Mz0w6wtNbCqQauL/tcsod8W
HblfoWdrUAEeUwAiymvGQwhZ2/T5MD9KrIoxN/bPeLGFRG+Q1QtP0/aAJ74VljDsDIS7vuDQCs1t
s9pGGIjQUv//UK5LLhSVL8rUEkk01buYLH2Fa6B0XkYq1qoOBbZMONRS5oueLYrSDrlRIc0oPj5p
/7N7PqqUKDdaWPMPm5MTeOksMmRsMqk8x22098GtsiSPLeoU7qEVNOmKCDIjCvVJi9k42ZB3J/Dx
OFf08zW6pEDjUxPbHZSty+byOCGA0n8W0tH6PvooFGww8/RqTm4p7vyjkBuaOA5vpWdJQbyoUMfV
KVa2I+xMCW2l7BXK9Ku2TmXaGF/r2WJCvdZyMg8VphGqCTqiAOqysiajaLVzpjpuFNLxPQNF2Z2k
CvBdbZYNPf+xYDzOMpAA0J81bjeB9YcWhNa1eWc2kv2qL7m8T6MJqOM96eKzAtiI0GFnAj9blz6N
l+TfWzctDBwI9FfdRX11u1iOG6U6zXcmod36qzEAmNXDbQZcYvHcBWCgdBZavsVgIMegUeCuF8qM
W/RePYaGw+Qbkrs9Xy4jUogX0El+AtbVUk5VDZKlX9oSbRHwRnJaTaAyaYUYqfCx7c89RdePFfvB
B+2tF1rqrp8GRljA2CWeNbrF3+aNpk5yszqU4XY7dkg1B+jn25s7936H64P+FHImK8nuGweGPC0E
P8vtU5GB6xEQpdNgbu8UQjpbKbs3x56/beZpdG+7yVO6TNikjclHg2QVQOLbqat/JFsO1ljmBKjh
+Jf6NlAT5tfd8eEr8Rwv8/1YF6ZefEAgF2+mAN4zgoWVWc0tt7VFFkDfB5mAe0OOzSGFf2k2JcKc
EnjY6aFeggh30IvcbnVZ/1HZNGtwz+BAJljAnHYNYlbALC9f7LN3v7YKmFl5n4XVT5Oyq/zHNj05
q3ELPgDhBbtnooYSDbh68mlaAMKxuSIzDfOtdEZws2qvTspuiJHDWUeKyFEtFGd6C7Bcn46z6e/7
Si7SwSfhueUGcH17PZLvmviXb/OHudrPE9PxnBFyJu3rc/3uEEDf6BFw7N7sYOyx79eSis3Q7m2j
k9bNL0r2kZCjkTG9RFS7LJh/+vnSnwygN5Zb4sqn9+oS1cMTdKTBovy9l0zO2xy9duivDLOkOaui
NIVE9AXRrdrK8iSPxBgnlXiMm6I9BEBQVtJrz+LKfgmKyWrCZR5Enn2rOYoVNjMUyTqwH+hWonyU
4xWClJDaYoq+ywbwS0E3PjHaOGNN6goUqnkac42ZQSl4nspifT3jd48IgaJ96jfrU/b9CzceRST7
2hIvUfIYi5j68cmXWwWZGGAv24UeTEqRs/HWTM/7naE8Y358i7i+krPxeHMXnBc7iJAa9BQGxEzL
yzrTOX7HLrvS+VyO9aeRny7dpDIEvUme/1qEP8iyNiu76wk0TyXB5LporciZzMuPQ2WCUuTftD9z
DND/QIjMHxc47jAgMVs80Co7p1SEC3IRuqyGXZ1Sjgq8W5ilVu8pVlCD3kO9vARoy7goyTcOgoxM
OuVYxd/rIAnVRV1WmDe7jukxSfMLSHzzdj6j4Z7LqhIeqiKaz9+bCIcOUAXSqi7cLUCVaioUtMmq
MmCxvOtuhp+T7Qibot0jJpplr3kHBhjRsP8sGjIqLrE/+beu3zyhcame6hiZlmmFeta7lGR8W1JT
Lw1RPw9A1thAi0S9oKPdgPL36w1W6MQexigzlauCEEPrwQrs+TC8AYNn5VRg41u8QKFcCf/pTqT+
BEpAnHP8xmaRHdaze+oQDBYvpDwLkhzcfNOnAih4d7yj8R9iqU7xUcqRM0UUS04KAMCKRXX9nmqu
+j8xjXG6uZsCFZH4/WGWA+byCOtS9PQLdglxfyrjV9GG3CcugY+2OecGLvxuf0aDd8ctetJ/TcRY
HQExmW/R/dGMS9Bqg1rpNMoODUIi8rgWjy27ozYe/HNlignyEMPdFa6ETH2cM+DDwaaDFSQijI9m
diNLtGjJ/CIiDrfx6rjU8uC64B7bzol3TnerFuwewaAQPY5CgkOUMC1zr88sOatACdqELwHQMe39
6foVRR2A2hTSVQXyfR86RdrMW0x6oF8gbjnqbnL5xO2pS1g2WYJob5LdsDkCs3e9M61tZ6rNg+3q
LFtSKyCHIyYz0DHjc5JQPhzA6amy53toBM9KjHvf2NQiuccTkUB2jkOJSI4vD9yDFNLld73gNsPP
bV+27sKTVFSpsVXDc7NQyhvxI3a4as7WcKjWlvO/oDJoM2GAmA0aKdSXhVV0XSA8UtBv3jTt0UTC
Wy8BDY+i8W6p4IwEAyzn6FIr2/We2Tlu9MdNWKWud4En9TkbVaqasLc+JbVWFX5Ncrhy0jFXCQcm
9DzmGt32RB4pvN4ue4hyJsvb1jV2BkQ7/IYNnZJm1HwebtbtQGXn2MdlNGsTqMFgpYdPEzQtLB8l
rBP3XQqjmwMom5/y9vUrb4Q5yb2bplmAPvcPttoYkAltht/jNYZRTP8p7MjGBSsAvhAha5gww+tf
8alx4PJjFFB1OI96F7rUH/p/zkcCPYIfJvUzQUlQCtMymzdVxnPrClVNLhsMuwUgsWsa72fNp5Ff
oWXPkGySwD8bvDPC2RtEGA64VUVWRRgcW3feyGqEZx8WO2wKrAoZPnC2jzW+migDPUt51Sy7y0KT
5yjdmY33r3zjEULLixHvdl76rbcfBRxoy1O10YzFGbFq/W6ICcAUmKIL9RL7wB2q37hFGpI9nH0y
EcbMQw5NQR/xVpZqlEPDxHH6UsFEDiIEfe/vm2xQszrQZcEF4bekXLVXlXooZF4f9Fv1swpbwYCO
o6axJvVzI28djTe3hTCzSRTnVp74p0ACB44ykPRrDeMnPaLAWV1uA4iEIYpq8vwE32lOmZruoDK8
evT5dIFBCs2cgYX5RR4ywFYyvH70GG9c/nBYBOIFHXArOFNqxcjqvKu9ztQoY9q4AR20UlQb+tpw
6e/Sc8aPe7qutv+jjHhzwYdwq32WSDzBLZXRiJa5wI0A1IoE1DALLz8h7tlRdWKorgPmaTbWzp43
DZYEQ3pYiGi58Q4ADwORhFXcIKy7Xld33mHlr5kQMF/eTIvLm4NeYaSs0PDvLX2xy4zkvvoxO3DC
9Q5/4rP3toZ54lPYosQ6S9rfaDx3olle5A0DNpyRMkawhfB/kG1028ett1DflHUKzSkdUB30xOqQ
+9N0ldgf32COp1lFcFtj3SoNb6LrigDbJn/2+eFxB9diMaGn907zceNpO6D7/MWlfifPYAQxn1SG
Cb6dqwyqTEFbNnqHe1bziWDVZicUmyvXWeItY1yc6VdTsDSWEHCwU4dMcY2lg74eURVJIAQWeF0C
fnlJs4GO1kZlGekzAQWU/1uW7sJPagQf81C845ley+xgq8Ia1yHx0pr0Z6TGAXzAOL28vsiYrp6H
3jPhFrGSeLizp4hspDTcdWF9rsIzbdjGD2wHZLQuo3YpN5O/twOynEwrSXqcileDPYucgxCNGVvk
0YBFxgAwPUiUrDd8+ZcgxTkv58J+IvDtaBA0UTE53qu8/JOt+8e55EpxkUZRgqK7BkPNNgc/zKS/
B1x5NMaZVlt+CoM/z1PtalumhpRzvrWB1mxCzAFMrj82k9P9Tv+2opLLuzF1Dr1lFZU1xP7JwJX4
Y4X+opsZQ0sGwF3KgcGaXgYN2faO5m5FGDNiPw1q1Sl7gEiW6pGeE178ZhamQ+q2ifZ32TKKh1aP
EQ9Aw7PEM6ZLO1A9Ac09Fcnq72l0dToEcWyx2x8QsW5RO+ptr5lRBtTRaFcGCC6hTrAlpZknpDwN
d7iYpHZ80vPoBoo5bI6VfLTmrcZ6P48QY5Tgd8BkPQY/7EfXbU1ujADMBWafhx4c8xN9wj9YZr+a
HJuggGpwYt0ynwp437FkK2jUOLW2OHheHXNyGn4yi8xeZwRsSk1ZAsMU91TF/Spf7UbObvNZa3kK
fpQXpD880BIZ5DfAe2+IrtqvVmqE58KV5eoM1GRQdDp7FQyzADs/OgloCaSObuQAZfi8QwWz+KB8
ixEmYbgxbz0oMQ+5O9HI9UKXvDoJT7fVZdyad/gtJAGU0dmiwwJ6ZQ//u5yUY0OMVo6Qe1x7x4Pt
PMvhVPOCl2tYWDCSkVB48660QYbxKwm2nFUZsfH4h7auWyWs917vFnvsoctVHbuLKIMBnXmtMCqu
7x06RfkFVAznFYNnLh3HXFeF0TxRqXMiDpKUBbahNc1w8HpYiGjeI8d8OQc53E/2pLOJy5W+1vmy
TXCAU7TMus1/L7VPduly99AHO+D0rcQgGPQBLhFQr8bUIomc2bsu+b7sW2WD6SEYt51K88Lj/azl
5p98xydBHSeUFNnI7jl5Upk//RMnylwduPb/fFjhxD+BgEdGVoYNZsG5NmOkuK7aBYJaoyU0byGa
P7ytZGkmhaAsJfRS7yuy4fHaWoQJMeEBF+vVC2TY5IO7/eGkRy8wC+rQraJTB0PndAuSx+UuUEfz
bpeq3LAUokWBBQdK3IiaQK/j1gd/Hz3whVfN81CcY6iBSYY+nlnECgskL9wWiVDV/IyTHopziSvg
wWV0SooX8iJTyMlnJtaO/7ZrSskY2mE1TUuOGBOW96/84ik2FcJiZI2pbvHElwLK4rwC+f5agqT5
nkBzNp+mjy/TCVzMnLv/4qmlMHXKWSc5IqC88irZGuF5Jeb2Ez/LTEFYPtd5J3765zvdUzUCbGUZ
KchB5/d90Kb3FKvMPVJ3ZAoexfhSzm3NfKHgdlrdd4jSMgEVQMTxzVeLkJeCucqzpHtnMBFUr4NE
QhldBT39HXBoeeF5OWzI+NKWf+BcJn4i+OOyj3knWmZWrXAxO0jxZMjc0uzxmRrmg7Wfe26YoYl8
VhjeAhFq0sM9NS+qMeDRz3vm0AcrvtXsVX8OgsNjqAuECE26HF5YQb5aVdM1hHThk4fu22IV3Jm/
xEshtsOvOX7YlO44koPs+5e7l2A4MKIx936pFL4j0ol+cv+dQEudW761ep1TvazMRl7dObreh/Yp
dobENRtaMx+11JoTU3G1YHUELS0Phqwyu7UDFEmZBSqYrt2cnz2CPTO1/hCXKMVRmk3OWbGBqBGN
iGIdUSqwEJXZifJKQag+PlwECzDT0RP0YsGp0sKB47nZEcxRz5kFXfQaVG7P/Upga8nocC9JoWEK
+XpdZrsbF/8ke39slMCNG96RCO3teC4Dij1Dugg/ps4TDq51X893R5c6Q2EI4YGI959mz+JZugUP
U869dFUQrc+T3K92WXLruwf2ShenErSbRFovJE+/+/2TcUJMk8cuproSzVPSj85o+2IZgUEGDVJ5
so3kGOdKrGqtAxP6SBuHShqw5qQ99tOdR5O14ziHJ3HpjycFQ9Pw9C/HSird9aLLBLjbJpgC4FYf
BzGc4C5O10Eolf9V9TAmHtbC4a1MB7nNdLaYF31CsGnLWep/ajg9+XDPskJo2QnvlJYYYU0/EQAG
vUEIvqNwnOOOH8GFo9woLIoK/AMPZjRyzlbYdpt9bx5IbbThVkRosLjA91lx7p2h60bxVVAKpXdV
HkvEVJgiOzVMgXgoA8pEHmqsVY//++v7FvrOH8+TTVCfpWojtTvhT6KCrKssm+oqczGBnW+MEL81
GdQTNQEeeMBDEGeUe+bWM8GEDAMq7STKDbH772WJLVthlR1IGAvx2GAx71mDjnXFlLuxTkl51DFV
NBpVZGxglOyHH1eusbOzUKe3j+ztJZPDXEOaBgmp8OsCJY/lPeh6h3oeYvngNqaAY3PX1/lGFsOD
hmAil4TPd185x617Rigv1zDaozqthyW8wrJge/id5ExnZpmOsESjqPniM6d7eYINxZI7r/tasUVz
LvX2INXux2lSGNwG34N0T5KsKuI8MOzy7nlDv39T6KnhQgu5RI4ABX2F4r3nz9SG/SV3gv4TBnBC
ryw82YP+j1CsHYI12z1f5WZkmfKHqmeVKOADzdowa4IDxb++6iqaK3GJJpOq1lc1PSqc7EYszd4W
OXkL0z+ASTTNti5nQmfPnyE9EXZxo8cD+sCXfl1C9rVxtIxkyBkFly8mnLuz3/PXsJ4J0NfX4ABh
DcVHP2yZK7vzBWSRD5zk78fvS1mtch98IytLFDMl7esjIEuVHUkeqfEzQq1vODdMyoCFAjJZy/zS
FwEJ15ak9fKZZzyXz1/LXdnrBxB5+B+IjiavlDrtKY4WwrcoQ6PmRPgbCHtq75YNXpvjKvEFqhKm
eeK48gyktfmJ4X10AOqTZfcQpWJUyetor3xpvnbsOcyN30n0qlew2+tx6RyW5XjdQ/aN/NOKGm8J
GafMQlvfnPzcfw1Fp10N7UVpYR7YQN97Fw6WHBeWP0oxgjqAtJP8kfTuSXtFS+pT0KGC9kRG3Qgj
jqw0M6Udp68geoeR06nW+RdxxL3oJEAhKeATMeS3T/aZYYIHbkpSRVoxnUQq9zEI9BBfOsLiG72T
O789LZc3Tj2k60EPPgEvjFe6jAIi1mOfQO6HDtZAD5ZZ6UljuTg8Q2jRPgbgIg1FYcycmu8bAKzV
IqMHS9c4h+crqfjNU1FTRgfCApUhTk/Fxy6jWnt4rtEXhhwPp0ZcJ4KYLjeRv0dM49YQ3gYlhPil
ScYM9ZCFbM0QjZXa1/9gERW425SQYLYXWgKEWDst0EzQMogdvw6XP1RV7EOrA6X2niWf2AfsLVy6
FcOebig2JcIhQ6f380Gmm62eCiO7JVJw/m1Leg9AmrXC8hjqfo5T32Ick7tEnxGsAMQ+1bTrOoMu
PUfI3xuMPUd9NiWtjxBON76fMkwU0vY6JBQQx1cu1tlfW20qIXtK/hO5R2P3wUYlVPpBzj/A2bzn
su6qs9NrZU38f4tA6oMsClblYVN42yrDFshMiMh8jih2ex5pxF1TA+N6Z/QUl1XwmqHCjpA36bkW
PFyXrBdD8rG7cSph96M8isBffQox6tH2dsio3lExAoxAS3lyL2+OUr+EKeE6/4CPznXtiNQrEV33
EgVX4R0JWyZ5qexXxHYjYVOAkwVmtGchF1gyNanPAz0aVD8xetJU6cjfK6UsAT6ptSauP0c2/O5X
69+WHD5Eeq2w31H+/o5vbArLGZYTKiysMJ0gv9yezxb21r/g9S/ksk97M5YUXTudtPUKLCOqaRLi
sv0h/x0G2yjFhoV61RoebLG9lCcF2Nan9qRlNVfWOTcaKkZSFEDMU0HvTtgXsUbUSLCpvkgHUy+T
w4jEtOCzRHBZlu12SCx2pVrjSGS4UnSW6kLjUeBWeOa3v731WDorw1+Qtq6y9LJkGUT1X1YFpZ/A
LWMg+mlfs143WSybxpxbiuyJcTpxrBQSz4xJF+C7vV6XzmZpFipaddUtOeg3bqUM0m3NUTrYd71o
5YrTDEEnnk0iCWRaPvFJsVjY0f9eUBc6LrGLm/fAx0r32XTDL6xjA4/qSjUktwysqKIGCQhDvo5a
wIlsiRsBH0yGra3x/6XSWFApBn9LBYesIVJ+0Oyvsm+9ebIzV6WMmgHAeRWKaAd2MepFEKtf1y0p
1mW3NCaFaMj4qDaVUWMXNjoRTMxTqrfNNvsR8Bh89PebjJqA47kh4+RF59+doFl356jQOxhF7mGB
39h+SaewQrUmR8Y4BdV+yJp+E7BvBqYBlg6lUuK+nmQzy+OKCrW6U95z9OHQvx1yA3QJriv8/YkP
xeQUpP6KRMbAbIdVn6fd+MPtq5D8ObYOCn3gMNapF+6BfI6LQ5RQRevpH21CXQbo45Ev3DE1AFLU
hf7/x7fXL8mojV7e8nYXbdieKKTF1PyBTQQ1JQzDXU5P4ODR87lqEJhoPlZU25luLa0n1m8RYGZV
RqOVIN4+R1wlASLwqG5ZqGioJVMfLJLHSwJ/bMZaHCTDG7pGOm9Ul1+k/NlkJDkLOCVdhvFHFvBo
d8AYoPWGw+8eC3xDg3QyaHur6Mz0MYZkrg1zLWHZaQeOvWGFF4maeDQ9fXZNf+hKSEP9+6NQgvbr
fj+d+bKPDiZHxzBhn8XD5RpJr1RMQuwXfnNXLUUET5Tg/uWBDL+3mxfJ2zq/58wpZ6etCK77r/PU
m5ueK3VYrqlnLXrhmaMkxrYhM006DAv+JhQOcQSIlED9YOTlWv460hAmFwlP0ymyJIyd0MGCTuNK
Hv+W5wb9v7bKErGs61Ux+QXQ+n3U3MYAvPIKWYJgngbrtLY49vROJdwT/hpFQC4RapQ8Frd4StmA
2yKoVp7VSCOM9znT711P2ojBiOcS2azK9Sg/dNGW7U+JOXPy4NmfUEu3xfJWcmxosB1LUI1H5UI+
/WbEmTaxRm+53D1SjcaaSoTnqioY24V/hgePba5tYUNfAfgjvpEGkn17GfbtBzF4mdWVhz/7k80H
DVSuIbnM7iYZZ3rk7ED2XuxyLrQle+pEqkkRFIQsGvKdYAw41Ej0kNWvsFi/JfrqZ6FtDgMBsZSI
YggPyuLIFHi13atwAe/LW7Q4JeYb1dT1Vltwl1JpMcL5LjkK7oQRvvMgBxe8oEnjuvES7O5kKzhQ
E8CiSxsfCPn+8FsVTc6tFhzLDx5bLBG3uKESnHqxa0YdZge3G9ahhNZGnjKpnV7Wg0XXWin8BF8N
GzTqKmJGY3lXtCxCjNK94/BTpVBqXz8AQ6SSMEDA0S56jgwIi2bm/Rvq6hhUvJ5lqj8NTc4yJ91J
4VShPk6yLmbP55hGJyPLrG4V7Ws71jdBqDoxBx1WfGbBDh1c3PrkLUXASIXSDlTISsIWzsdb+ciK
mDNY+BixbwX2y2r4GdW6Aj68uU2D161T+SFpi8NwCjUx7US6eO2/hW+bunLeHikdq3mBcTaVRwuC
6Z6YRmy1hcXBK/l/8mV0vBeNfhY54KuBdXfalB4Cje32Rj0gwXkZnvOP4Zu2siKDSxaryuQ3Lr75
ZqaCzReM0gZrrHjHqgaJEmGYNuOyV63k1KwT1APJZXhy+C2ZcjIDrTs4OsWlnr3Zj6Lrfm5/3FQj
89kabjPB3fwWHVFlCXkWMKpGe9L24s3ITi0NkDOK3UaSCC4rMrFDGSPfsRfuKqM2LpSxAuN26Z7v
9gpV4GnX5JqmF3WLoN064pjs3LPE2PmKCOCpDWRrqTUyRTr+6G6o8F5Y2YB5W2NPedYVZugHuh4Q
IeczDp5q6nmM2Sige8MtopGhD3zclHF1mZ6FVUb+noxA0Tn38auX6hiaaasLjcgC8KRDLci2Dv3j
AYO6fA9he8cBYHESRTPg1pUR1xeUjhAb/M14AGj8qo6O5erpYDJNMsgkEBzmdx/3aB0GRWQkbNx1
A0IdVA40WEoMZXf08t+uqgYdak25U+7RbR160QlCzYA0Q0gkZErC53PTv8wZx3mloeSBH3Sngaic
T4l/g9izcycDrSJtqE/060KQtoJxgqvHqb85zwmMVxBMFWtAzb80vVTKdDxS/LtbOAScJ64VR2ko
rwCn9TnhlibwiSEjVCli3cDIjN6KYcFHdTamWncp+RBBPJfhCDvqIoRkmdZkuAM+N0HT7o52B1aB
0YT4tNv/JxgxPhO2JWDAmaEKVQTKob/fdE+ZsJl2+SGT8a4MdiaK8UokiNEwMbKkbwCGAbNCUygu
XCJzUxEIgu3QR04CxmjR7KyIPyZN9yquf7o1DNQqoRVYyEImj55HHtudycrVeuE2JhfcnoGyRtTZ
XSsPmgVAwDIZXc3KDWB90n9WWWHb7olc3kRv3mPDMqlGtrr3UJiQwaU9pJ+r3H8iE+DO2grjkUbo
AQQLxZ9g6Oo7OEhIp1zisCZ8T0hbIo4mF4+SQWyok5uO3ZZxhqik4/s7+mHXnpmJ7Shk/OmnEb5q
gd33vfsksrbaiQ6xK0ZuD6c35gq7WTtyP8ViGvWf1bkL6Ur4Ya7d9Pvz520agMY8FY33qCbzROKf
WDEOacQYSGrX9Ge8PsoRPOsMzfqgfmbMexuHKxm+G1fxAgBOoXlcICaQ0K4nqDY4hTzshYSAgFf7
4zGWuDHTI5jpzaLW06oCYoBYVClztllAusWT7ICKoLGVT+DA565NW3fY+sgh0FEu1v+OOj3aMUjV
IpEDYccKakSQ9kpGF1dXeKxNHfcbnX5sBIpxqN5pbkiR9EKVK9tlXcm6ZTflSzajH1CSm8mw/EvN
AH9le+UBFMYHLEaUdXeCusB9mu3nwwrimJcPmgu/ta31oQHuDQnyKETyfSgUIAZwyHb+ez5Vuk5R
bnYmgtcYnW2Rr6YgUJpaXaGwcmoLL8ayEAkLB2i7qS6tp7g9M0GQTCgXxMgPiKTM62yPS+qKJuck
lZFyNFCssFXKwBxBktldCPEQMmkSUBrKvyytAGrBFmB8kGroZiaTfrZlhDdh2txo2HcjfhUsdaDl
s3ALnDvFKBGqUJt3fSgXaRxJ9UAevsmnjCRMw9MWQAxSw8a3kVfQOpkw11BjzY6tme0sQudt+USn
UkDIesRwoN1Up0IbGzoZ3uy0m5K3LcYbgxyt3FMYbpitkHVmbMPBJ9ru+OnG+CxV2B9QSvBZSrwT
mYeLz/5JzmGmBQmMblQZz1nW8hc6f79B3uQB3DSgaBteoMpp2E+66PPN+oAXVXhijVnC6O1FY7bl
xlldTLU84td68x7hp4tG7PFqKdSz7KAqeELU+mhNKJl9zfulLOukS2k2fl+++v5Q8dn2geHoMCEA
ZZ1JX1KeS3w2eNOybt+a8JwMYWzceLlenZ3Wk/4RvJgc8DrpkkuxKGGqnW3kI39rCLZQU4XcgKAA
fi2mKOBJIpfxInJ4YlZUf112B/40rvUajRyphsXt/z7CeDyKOiVNYditmcDWAy20evlxm53wt129
q96l5aswfCxBs3E1uvTXVUr7qIgrJ5U9OR7uCJrId4hqwvrTgKy4qfO/iRBbQ9OlgIp7Htx4Goix
ywG4vNOLiFtbX7/jvCcHfJnxy5YatApJmBQyCYAfAwG0PzpFy1txNdf/ZC3LsotAHNNZ+jbhUS5o
nc4hiY/EVAxdJqk5BzhPtHoVSYJ7j2w5msGd9zIRuC6JABRqvjFQYTh+szNokhFfliqIqlTYcVK/
ffaYDlm1YjtYm+pfPe/K3LcVuH28c02N7qtHp/QfnZ1tcRPBB+BUvuGvSl5AATawDAq4vcwNZWlG
Y7CGF+uLaQX0WYKiRgA5WrkFEns0Ih8QYKipffNO/9HgAhlKE/nIrFgnsyd2JP4/5TGPPWvCbqgY
G3pd7BcCAG2OuT8vw+PJocrFVfqJnNnl3EvhYvE1iEoSZ1RbE/6CoT/Yvdu7QfFiNuOp6FiiUujR
yyw0c1AJm1l7d3yCRhxixj+ZepSDzFfxrO06EbuziyuRdVEE8oyiMM96b/FG3sLyJYaUs0873fZZ
5Zs3DFgvRQjtD6SChl8Qrn/tI6DGnKYKXDGz4P6p+xNA0LsbN0DDBtJTnH9d34G3nMIN1t1vroWK
0Y/WtctiP2GN+ygEPIyxHns2Od+Ih1DjMu9iKKn2kGXmTIGB0qBrL/JKOj/pW0aV9ltxI4/WCY/v
Jt5z5Vb5WvO/zhGGorNrSJMG1w6+PmPl8Y0i1MB3HVxb1mb6cQIGaLVyJ6o2uI/trgHw8qJB89HJ
eVd56ZMUTkNab/D/VtFLUHcNflhYnyZaEiwZ329kt4TtNSy57SbieVMJxjq3caxiZv3D5TWhSWJ5
EuIRaktF2/4L5o58GFVpp3C+ZArlIvYOqXk+6DLg1ltiEYeETndqw9Gc/Uofm9XfMzdNYQK4hhP5
OaN0QQEXrCi/jnJGq5TMatTgyBLFcHoW6SWosSaXyF7FF/i7fWfAHTglq3Y8gqQNDC/6ACs+qpVj
s0FqHenTW7FIEv7LdX0Sof0jv9uUvp4LnRN9+gIgN2K7FwegF97SNiglHJWECtMqV7ZbMhBVn/cN
QXxk6EC5zQWmdFCyU4V5rEiyki9WHGAmDd6nQTkw8Eppa6VxeIm0qYp1mzqLkwxXo1paAU0az5Di
zZhT9mtkcHxeWyXIOXzbCM6vBVbeEczs8+7V3bJdDPWIXxLpFmK5B0wHTjx0BfWZsMs8KIl4TsVe
gjSfftdKEcQ2tHY7mlQ97n4PyR/M0k65+J2Cc940xDNWmkaScWNNsSJRE0p3LGPDd0BLe9wXfBI/
7Z3w85iafo7lcnOqo3no4i7iTEUYbEVUhmZI/vcFwsKNaICAVRgtHQCeMQsCZkutpAZ2QRg9jT6a
w6pn8/UJM8ErLt4/rPzNswXY488UbR58QkjsxV51sIk8TCtwB4iIaLyww/b8tC0vjsKWy3vQTMcZ
wgTWsyyp54izktfHeXMAN1IlYv3jd2MJlNNNF6VykXOmKzfHjiy3mQSamAD0FYA9FpZJ4OmJhwSO
XFWkVdnsewP25MHS5MtYja8x6FtPtdB3JHpczj/6pupO7XOaBoATFthFKucgRt6/+mNAISm8023E
ok3Bs2NFGq3OdpwSBLfY2XeTYnlwUPSyAkZemQEqrSmbRs2m5bHB7xIYVaooSeHJdCuK2pVDsA/h
dMowMLVoLk3QkUHIKutrTND4NJA02vMXTZRcDoU4hH2t2vlJmiZBaVHtOHvL7omWD9vpVW2KyV0P
pH2SpymtDx+1W4ks+8lUdZRvZYRP+U0PfI/2mBKhx5Yu6FaBzvh1E+T2JqLNsv4L+SDUAOb90fOA
TdmjtoDpTuhvbG7IlWek2nFeZmWFiwkOI68P8lmcXNmwzDqyzVlQPqPouwXN/k2C1k+vR5RJ51n8
oTN6cG4d5RzgL3bJ/ZF+rzbza2SUUUzeOLAnEF1LWGjZcKEEr4cV0nf7QOsecTdIHWA//nrxlXLD
O7LpM7ebMDwdx87OeuDYNc3SnpAFqNazw3amChpbA6BzEtEdRMfAcUUhJ97CjMtRYUoOw/43wLlh
vCIi8xyS20M8gu8yIYCuv9ffz1N/7XM+QfEQ3FOUI6WkjmIl4gXciDXcVXfQgNl3LGPjuRpOBDoZ
wHM/eIntrpneZd8YcSuvMDb3dQspgdnQ8tExWnWqyfxW3Vixt7yNEqrhcHuZR5tyMh/OA3nk7KOq
VKpBpRv9O8Iye6JAWcU/HIx//YwD14BselOF8cy7S5LzOtKMwJBARhgoJyC/Vr9NYw/KeiiS0Kll
NQhcyzXHW6bYeWE23jQKW5s9uznlyZxkO++LjpXE4sODeQix3MNIv+S5MO7RSs/YVyrCMmHspCeg
aPiAPjfGy1qDpQU9WYS7wP/dEoOEjuo0c0zeO8meBGLHimIL+GDnnILlC9VTk2q61sWPwyPHRAnb
vsEOmBI3AFcn8xskR9bDiqeowp+XMGbXWmhp7ofGKRUNMXjxTAds/Ix9GEn5yRSbY2+N51nr1txV
WyXcctb30MHi9uVWCGF3batXm0FDD532VWk5I3aYK4sq5MIDLUSzAw2deT/7H6r2k5HkBqUHnHcG
uDF2ZCQswZC827wk6hlFkl+AZA+ZbEzF/hJTloDKN3mQ06L5bEqN5FRcC93H3t8N8nX4xQf4TIWj
G7W6EQRNJ1UrT2SR9HdhBpK6pXKn9nMfds6Epc6GZTpKL/X2TEK8zYIeuDd/0tl7altfbC6fsedK
NsvhSyL9/rGGi2xoXeM/1KGKre9kc7knG4wd/rshFGc3l/DOFTVU+D569BL3G/C8NYsQFA1iztoQ
Jgxm54MGAERDLEXGg5aHjrVHqqwVZufilk3Yfy7QRIgP4JyWpahZkgM3fKogtq8v0kUWIZEe5GUV
1QCWKhiUSB/qLHsRFOIqWrIpTopUNvpQXirWNKvewgQj0FgzQ/6BQ8RGSoPItCuOR7IsOrWgztqf
3tLDD8xQuki1OAK8uXmr3DmxE++3exGP9CTmCkMfJ0Ce3j08eoj/7MbDS4gJm1q9UY7bz1Rmm8ge
vD4JTBv64DP4C+fiRJ7iyyLTOWYDUZ5BtnPnh4nOerLfQS7g8h6eqnuu4K14EqtV+euXb+MIMSU+
QloujWPvjjCf7zsXaNUpSGBW/tDm2nGAXiiRT/kScMZHwoKZJWdIY7T5FjIsgldZRdhOr5B1syHX
e+bvgYZQ5fmVo7scF5GwDPfJ9z2g5ZK9K86VfoN4JnqtxCTEL89yPPkqtuYYPVNn9Rs+vuLJQD7T
7qdkgN8xUr/6jwkp9mtIr3dOFkvjDZSi9FRlIOpcAtS68FChT+nM6LLOzZDV5Eb49LcRVcDQrknK
k6Lu00lsIO/xRmETtc7uwiU9gVioPliMNzQbu3+zGmSYgJTzVUzZ5k6yXViK5W9LycHPY9VMaIom
hVjAzEiaoUHI7wI3nbe61FyzmKr7ex2jJBI7gKfB7u09E9stmcECppxiQJaAxrarJh8O3yEiAdOJ
JkZgSQ5st9+BJWqOsdhGSq2X8KdaIPfGFR21NqGapi9b4nKWrvW+80GBIkhktdFgWy4cpGtovOa8
x88FlbGZGd3kqPlPDnrL6eOQCowQRcmlh1rGffgeyF58JJ5gSKQR7kq2/aHJqoe7114PGkOElE5h
XjUTpUV3lo2SWU8fFpx5vv4/F4Aw6Mk63BuJK+g5n7yCptP9U9SD+MedvhcnPUgbgcurdWlNmCeG
kH1661/kpv26NEPv1sBDpiBn/BQvt+NjLq3oMOPkr3qcYqEED3zuV8hCoSH/t91BzLNy3S3CK1w6
qHwfMthaLctLCM/m6B9mRJfR57kKT6d72y8rVhLGZbCGMG6SbEoTUS5E13jYUhf6wgWWjxhMYdth
NzcKi44aWzs2QLoA/W9F4h22QdNdvSIA1FAm4UWH31uA9mU4mc21f8JM8nz6yDJQiVRZmWLmksUG
YRZVlE6a/cwAHiCaya42ettNMAnY/uGaw8SPIFBOEE800zecnHjfEsdY7moF1nkat7sEJ2X85pm6
bg1PllG3dNhe58QH2qxHLNq5a6wFHOEzX5x28EhRaeO5aJHoIpFMu6yxLRRrETi7A0NtOfdUMdkF
MusoXglHxpQ8fJ7wwSIt+tOfLlZL2qwQd/PqI99XBxBYl7yEP2uzkZWp9baLvgDGVIUGxi15K62X
VB6ZkgcaP6QBg97NsHk1C0aeoeA46RwKUV0N9VNbp+X3oFm7N8kOrBolrvn3cDHiGVAxykQa7i1Y
UXZKcfE4PbOfLKXp7R0GSJqNj3z52B4aJkJVCvSXPSWyfhN2cH9/+FzcDrrC0IbPCPgl+eDK2cLB
POovgqU8K8/fDfDJ3uBQwlJbDrkPz6iJ4BllnFe0EoX8apZj45Q/SlX2Rb0+wqvwfmqrbUgQNPbg
ZxJSb0PVV25PO16LHUJ6kJ3Br09lvoOUCb6RnnH89Tsk7V1tk6yncjUgV/uGpg9sP0WlgPpOWJY2
q5acnGV6wzTjxZG9FdCsjUyX/L+UU8xlNf57rY8CSBa9bTQJfKIGxL8Kznh2dhK57m723IP5J46o
S8bH3b1QMuvJTVWL3wYb8A/Fi6AQmF2YbOk+pfs/lORAy5I5GbcG7W3E81RiKIgBukXvxsM83bix
UaJ/AQEBOsK4s6D4ZNpEpuCgf1RTVAU7lGq73vr6sAcLMtfx/r69DBK1Lzb3k9pEuq8QfFoJ1CJp
6Z601/YxBjGZ6ZtgJpkpcq2Q8Ad0W6up+r8LxGqThJL0fiQ5vHSWIgJbQthVLhD8KfizYPSt20Jd
LMFCgMU1GwUzUFBXC1+KFU9W36oz1YLZiddUaTrBCKh7ixCCHPQeon438jISMpsFNCJsRFGvKsAI
IkAiSCJxkD8MHnWZagY+uPn2R97JvIsZbNi/5JFpxz307wcvVZkEBK5G0qNhjOoG+62ovo4hqxdZ
7hs3oRI3Tx7qFWjKFPlGODVIwTDVDNBqNGNNSzzkBBDCXnXJ17x4lo0bPEfyWg6Jb1MjcF9lKebX
gqnPmXwHpOuuy3dxt/n7FUa1q+hwmkoPAciMBRbXOfuA8uOZRn8TfPEC/b4KeNYaBv/94UF1WV7p
NR93mnuWuPT4jhPm73RlZ0hQfRCYM4yFZtaBUOdJM3TBNJl6Pl+8uxJEpUYvoxrZ/e/XVGqeguyM
lpUrxQNj9VESoyV4Y/woNV0xkTvdqPrpClTityLvevFnKg/feeSBT1Dh8CF/a8lMYzLBrE9i9Alq
GvY/XW134lg3rz0gU0f2hH4kLAmF4dqzJjDTfd68tpvPZo+Sk29/VS4U3ugxxzVp904qVczMoulq
uWHCb3uMftGuwjNF6TFDU9fNh1V5xdDSI0iNCYp4NcRnLTinIFHKOr3gG9JzorLMq2D6z7Pv6+w2
m5DKU4UNiQyH7GmPCccGnSDHrfh02Y0X5Bh6CrDOAcB5B9/7o8oyTs8Rklm50oNHPTgq5hRGmAW8
7RficdT7vcSYp9eK4tZDMeFfGXybmV7qHn1npfQrilCKNB9e1tWdIAS0qraM6P2HpqcKfvV42ING
HRvJlTKFi2FxLfd9SuJrtebsNcCMOk8mFmQ0JzcRWxTvUxHyAk2ZXU86s4Q56YpWtn3vR3JAlopq
+hSWcIkUrj/R4nSsHL4rpAKad9xobr84BY40V1GIKrZBcqxBv+rxz+6lpwNnZ1j30tgG0WaVQbuC
+LNTpweV0uc8x3Ql/flJHvDe6gQeRUiDlA+xh29XWOLlJiJ6CQsJxVUkB4l0yUycG/v/K0VQl76p
capiycrhTDKS+sYaoE+1ff1gct2MyzavFrHci3Gyf5C1KCc+wyogesz8pMEt7PAYvww7+ePjD87k
nFNNvkl1CfRGrjgS7VfpsWGbF4xBg6PH3BTxP5I37qM3O+Dms03HVIV3Ud7xqSy5Z702UMpJQqKB
hmwXTKn1wk7imQmIHb+L8W1sA+lWUn5ngDeqOYzMcsB7ysKl2faULqChnVcuUYVYyORZbGyzO3iQ
cFQtfWxZip68W77tQm1OmGeBmJPQKil2DIibcL3a5wHFjtDCZ3T9tcqGzsrZacBA5Edr6PFsMqqm
fvIallHwYWPmJVaUcxLAO1oPuDwwU+sJ6B/ppqTl5Wz1HEVgYpqion3bjNW6MZEqsDaLqIS+wayh
gI+6bO/n1w2l05wx72REH4P6C9QvrSIXxozzKgv8dQNagc3zqakGcZfzoR0YpLv83lzpOzEqkY5K
0JW9ozyc3gYw9wYKIPeV1pZSNPp/hRIPAGKJ2TGHfyvXxj2yCVjby1Ze0xrf3gXmbAK/89oCHTVq
aPoZz6V39kqzjszmmgpXFcIgjm0ThTU956h4MHvyQi3Oz8zbgJK0Lrjdzfp2V337x0/+wHcRPWrW
FDNMkTrEJQSspQsfdhBjv8WMo6wcqBsL1IzMF12fCQuAeiCDs6ew5OsjcuTT3Skhqm/Hs54274uw
SU1DYfZqdLHeKrwKp6iNaAWcjQKmX2Ba2LgPsN0NVFdXnym3U0KMxCGI5k/bkwhzpGyyah+uLILS
S2perRht1oumuthqJl3nLDsJyUAvRdiRjjd294LjbCww6KCMykD6dp1wnwZf4ZWwAn9jLmqhfuq8
bI4qqL5tC98NCMRICNP96eG1BW4170KjEw5sm91OjfpcsrjjBrXwHOeh17vRNXWrwBIDmDx8VWxr
oS5gZFnfEQK0Neg+Rr3igrZmhmhF+WKuVWihe9tr3cGJwt69tyuWJFEDp+BufFL4bD8mWf2CcoX3
GAChR1dXFN6GmkICEYvxDXu7qySU93tD4IJfjjtllgntgMWqAkkA7+yWxizZIGUIa0c4yihZV0tj
z4xMu0AENS7p28hKq3QgARyGLm4i1xiihblc0JsefQbeoDAG/YuHN0dJXeUY2cfSafF/hFpf6Ddx
HWKlvIQxluoqQd/vNv+WTe9mrKEN6+zamhDjjUQGi0I9kgk3uJ3CXeSAaU3KyjmHN5o8o5ZUydNz
vOLsoX0hN3cP/h/sNk/JGL5zEXZzL0Ey80MgICiFT5s+29KFu9AUO2M5NhrNAr2Mt82QkMMov7ZX
5OTuhUouEpp0LCh2JwFxmXtRpMVy25RGcULjC/863SdYV/c2PSvwaDrUA5XsDHFswYLvBYidWdiS
B0oBh9j7hGS7C9/m4UX9QEAHcaB1kNgHYNoypGIVdapsg5ttJgMooR+cvN9yqwekEG4sybjXEsSn
gde3vcO4PGTF5ht1UVlBzieATLFdDWL0/EM+DlkVZscivYTUl9oy66Wmam28jqyyMhDkJy8oP72q
8wRiUmXCo+VnxpFFal2cfWnZRiKLBTna5anmw3JZ6ZDUd7+CKvoIQevOEDke92VJe6l24W/ZvVan
NCOkIJ1eKvezP+73GJVsbRcK6SqaSIpYuPhgZ3ox1ATrklukbJKp68T0TZldPDUngM1xdgEgGQLz
9jyehyFu5Drq/n+ueOetg6HsoTMu42cTq7QOf8sZHdxzyokt3S3dl9fJAqvB81ztZUWUORFcU04l
Rj+NBqWPTjCb2YzwKBO6Dg36m0MF787PHfAAl1KL+jysuI2rAMN/0wGt57+kUmxqOn4nrnq2YgcA
+vWltEjMbWEWgi2iXgKQe9VODdkj2zloKj09t/zSEuEcDk0VXEG3z7+PkxxiFRqaIok44ZoPiKNj
Kj8CQlmyuBDShxFX5NDCGRGc1hu6mQx8V4KDL6UR9ZQ5RzzCfXnO/z4FdPwIjmwZATOEJM4JvjcC
2ISYXy2G9t3YvTM+DVBG5hfe+dF5v8VWwp7VvrpIF2rQ5nbfrOUxWJCLpiu9fcDVY6gnnSbM0nDO
KICCSAAYVqbOI/3fqfLU7YvxtcJ/CIS1cZiY9M2+qd2qCjdxjdCgCLCDhxqmdPgy+Pwqfd74M39D
LJ+y0Vvrs5pdHmPDc1N4pyt0Kdki0ZSaN1Z5BhB9D3K4WG3sFeQ1AXGlIf8RJsCyfPbpg+f1G55d
Tvb7YnlVlITNWnH5sES8RSf5ixo1StvTeMs3qTYu0oBKkRwq6wt50eAFAe/fFi0xFziVBJKDRwFX
S4o5SR0ASHlLtTFMPEWIj8qDGeeQyApSrukQV7b8BERJ8rLsmhd4055uWRW1vwFY0JEzepzC3e1+
hUziOmJ7kYZ5Ip/eexjfEVxYAY1BXuaa5/JwDJw194L48OkwRu3j+MjzuQNyuFlwzh1mKvYWHRUv
A7Zxz7OMmmmJESPJT//5PuVVmn5OnB1R3Hd3T1n/Xh4O3Z2bz8/etmMkWpZ0G5RNBjwgn7Wzckia
iSh0kzHK+d2J8GWvLjvle96bNMOGc5VfSXRgGtyb5oZKqd+gawqbv3v10F5dqcQncxwcUjVvRKhD
HDUjzoeg6TmzSURbtNb09dF10DoSBm1Iv63gNAJfmkRyB6SwAK1YhRJogSQcax3XAyAr4YmnatWp
t0y5zrb4ocBSpchbcFZxzvu9Kh9rT3m4E40+BKizJzRCo2JDeYTqfxtExlggUmlXNkzrOvQ5khKV
TkRJuVN+oRquyBat3TDKfjZU2Zy7OyoebG7gpXkUCBRMSC/ZYkZ8tv3VnrXeu0QSRb44PI59GE8U
djmm4Hy2C7V8BcHIIQyoZn+8F7BQhX7huo/odco6WkfG/aXnYCSmSMpFef72mj26jleJroPtpixq
StWilu6k3ADQZsLYbHQXF11A2u8gAiabO5RM+aMfL2euVi9YDmShxSqT5aRNdT502oUnA561fBpq
QLuVWp0zrJLN3wz99077+zhfCuEdNR+JQ014pqWq8DF+OzTxSrxWpfvQ2r8ycUdcmhsi7zm2KKfQ
ml3B4WxknIYZOWM2mN5oe8180ON3J26FVSV6NbUpDeG3AC6qQX3o13OTNu87qLNjwG+/cy4DrDm5
dbe3fqBkA1ZnWjs0Xq09/V38FFHsOO9560+N6YYU0v/MHgihDvV982NakfNnMqgGgSB6gGCBC/+2
IAnuUMEsQM2TGqbV8jGZKfivSnhwTdfXxu6lQEXO2dsGPRYz3CyNwe1CdDYwHaGY7DBQqFy3+T3D
ZhVfVMKdfIwKbc17UoOAKVu7+Sey1I2qVXmiNzAcXBpMAvbiKrWssZuu87xaJOXFGSphvANsFBvB
/yDIGB2wwSO6gBWTevhkLJqqjjGdyIDSzJcPA4VLSY8JNBx6CLQG+WwoouLK/7Thxnbbl4/phEiI
XQrMUjzsKCpmmTyXwvTGPLG3xWFlsl6Rxo1u0kUPqvr0vZzG40HvZ/JoyZJoTgFkwRjuNuQ6F4zy
j3KlfdYIaNYT181eH27zl8S/vizPA18ptDDn3VMuNIaCePHh1WzXETTi+SJ4QXiMhSK9LEE3NRd7
498b3evVh+I0aemu9lXaveg9qcCoLHxpaIpbBz04hw9VjIXwMoeCoCDGMRQ84w4y7zA4KKRyjPA/
eY4/2UctsMwH2ExwHICOD9DvhF0K4sPq2/u2sPQfrb52f00wGwUXK8HdSoPa7Odr1VzOup16hK46
jqFZL5cfdDIiMM9MhBxYurtIKPI/92HkqNOvjrsyr8BRnnhPg2IMyy+LizYKxT/sJQSI3sN/87Aw
Hq+6k4XqpVZJay6viYtqqyVMBND0Ow7ltv1mnUPUDTByvPRYDphCSuDlATrYyevthAExSxE157BS
C8L69MCOIC53MaQT6Jm2cPeX5ISBKqlc9yWAEtoIQmLCzRwNs1tjVrG0EqM7Kc+w0+QVE7vhoNEG
lkKmDmDTjSx2/WUh+TxLQ82x9dDHceFkSk3dRkwo9tm3fFxTC7t4SiMl/PZBDB2RPdWGkGQWX1mT
UT4E4kbAI1mYsbzAHrLoNSPKyO/8rbqogXbJHdNI5rox1eb9KRRgdfz0xGd4apPBog4Nm/rqHxv7
1nSOYZ5ZpVBWa9lKuxYLzBze74LVciah69k9kbF67eqODcHIlBiqRNNCz1Kze3rEKpvVvwi/XoBU
ioExOuIi6ZDLdqaPu+AUIaU13WtBVuKSXT+kBQhSplNItPaU0kg+bGI9X8Mstsw8DGQXkxey976z
RsjuivbpEp+T2hxP7ct9zeVfWPU054TzD5rgxjKKUM9StSRXoJKUdoFzGftXaPril922c4i/Mjlt
Q4Gf00f4On4SGTaq5VxlXYuYIsXFW+yEDD4RxZfMk1tdTcbnk5KlDWZzQZ2poUACe6u41TQMTWiX
U8q03uBngiD2NrhOR0p8tfCZ74CyNK22CATWXWCtG7AJ22JxD+b51t4AG1LlSSi93KA0QOftZBJE
Ltz+kDNiTA0wf24mPuGWzT23N6dhDEzQ6aw70M+iw8HMbH1n+Dy1nSUnFSxrXFfJzEwSQFK9qc7D
GV1NqhzrAIoH0xLv60L75wkPjVXLnFAe9E2D9eE8GzVNJh4biMJ1Y5Te5iyjEOTJlnfGjgfhmxKv
d02TSuE41oWub3cBE6fAa8Ja0XGX5KS4IVKfLV/0IwIJAXL79yVJtVnyVLApsAh3+6SeNIePvPbf
fcdWO740E41El1bBrY2d9Y4VTSTi8WcAGMUGOUPBpWyeH5jwYAq9ypi0ZuRLzjDNEryBO1nBC2ho
IQv+hYYZUYDrHp1ZWKlw/6xRcstQkovzVGB2kN+cEa17SdE3LToSCWSGvEOpiNzavA73eO9ATddE
gxlmd/5kirnfhIgFkpR1tyepyPebJLQMxlrIB5THk0FnYNvfEU0caPKrtZ4OD3Dpsz2vRhIl1NTT
MaU+RX6ayl/mkjxaUs9RlrV/Ll+0tQqFivzIzjllnwZv8OI2UIqrM4Zdy9quO8TtaOHqhnP4XOif
WnNhks89fp8RO9Ur32VsXPuY/YEjDmDeCMk0w6N3gzy+6lUbp9aohhzgHajsjNBrQc24rc5X+aVQ
KU9zTHCB7yWlLZIq6GJJy5IVuGUGmriAajqjkgOgmUczQRMGmxeimMLNZTC5ulP44Cb7zJQ2zWa1
DiySP7RiUFGqCcEydTyxHFnQx3KYj7AnucFvzVs6BZP0Dp8d+3QXIeYLAq8Q6J5bdwhRxzZfhNIP
DjsqKT+SchciCrLwodwS7jNaeHXfyzcF3yZwoH9FKEmtf8CJnH1/348BHerHJ9rjz69D1i23j8Im
yqAaO8rNFL1fGhgzWLcfhX1ZPXUSyQBCbf1X9+k3nOFKFyxlTjBP9Yfq2hyaE+hlFCzRS7Vf6cWy
BkpVpcNUqUzd3Dh/tVrRKBU9vTR8udhYYiZNC1JynPEifW0X0K4ILBlhdovWi2K4nRA7qD92nNRd
sHcUXPHszAPoXwpfN4jTBc9tkic5xqC/tEZPBEURIrXJQXLQTkmSkcnLmGXjGxEbpza3p+2iYxnq
zQZg1M0jf+HO9j/cDfpg9uhKWl6L4rK7ISQGrMG0TD6IDYeoqp1moxZ1ZchFM8Fnmgz7o6lJIwZD
6v00Ztb0IHVl10OJHvROXvTZVsblFJMXp+Spt+hsqtiZhBI2nj1Gg8U1cQ7kvgW+/u4hD71bJDvh
IyxGBPB/EJBwAUTdMQW/ULqWhMYhQBjjKyl82J4G48YASZ7xzGzqD4l54D1CvK/OSvzYMuWkuX5e
H5KU0jrw++k7pod+cOm0XbnGngcjJ+OGDThh8PLh0GDWHS8QJyj3ivdHeQf4J9+qx9Vk8SUtSl6p
ZWJhm177JvnupJ3xWvkTkOrNabU6najlNNCu58IPTFsxrAA+TqOCqtQPyB99G8WxP8ZcxokkJclq
uAwW6k4APMtalXgxUoZ3SgLwGhxYJ74d0JPU/6JwpyO/eN2/PnX7twFRzYw7MIH4AZtNyXRRByiw
94Q/bTIRG3xWxJuvBiw2fB7PHUGyK3xO+EfiL+KzBADSmNfZKdkGCDIJA9xGLXauBA6SsC8SZrOr
qNoxSLBs57SQgstd8bUUPBmBHM0Qgu0hSjL7Bk1kDQ9DH+SqTz5mQmrSc6K4fwLC9/jZdeQ+7eOT
0J0L7H1Eu3CbWNnKzV2MOsay7kPat8XJmDMdG4a4c4PNwh2JeVe6+sHL/GzwoYwNKLAaAF9x36wX
IM7VzRQxlfuqXHfCM3virJP7DdHuqNY2wYGaJlvuklHWaZu1fYyLygXMPfUNW5YxKISA/I2XNfaS
wYOGwTgl0fWqB/YdWzDhGVFVAnOaNfZaid5zB3ZZzkC1ri0xbLF0PB+Y9zQkTkJlMHAWYTS6By9t
lHONDK8mVqkCFj9oaNzKWuw+96wIYy8p/k7UA4GxrWrBim2+jlWEfq0AtyRHdkzXparDP2NRi1Kd
b7uV+Zw3/epOILeGlcsgSLl6bgMBKq0QwVc3CH9b2mC3quURe/FYyTPuQKejRAq/4oEA4s5zoDD1
k6SOIV2DkbFeALuG3YXCI/oPdeeksI22ENhOkpAqRW0KbI+CzNKIPoKjnYY58TqOldwBfBGSc/V9
qiEvjK2x+cjwK3MYqoiRYGHS8sMxtgZ3zlUD2UMSOc9Esrm4lcO/KestwTVAQLEexvX8/ZLdUO/U
XfolzuMgVbVTrGl9HmS41p/cEHykHc7p25vpo7l2QQSPDwsyuU4AkuDM37xFx+MAkKuhNSgIXQcs
t1O82IwGYtvC1DzBBRX8Nf9aCJLYUaWehQgJCgYHdbphWpfC7tb8Ft5DChyZEtRVmjMLMgFnFS9l
MytxZ9BD4z20nd+eSVaFy4vX2LeZDqJ/gT/F5foqLTXT958uVITPxTfXgC3R/cHAwi/uIkq1nhj6
X/AlPSnKQXmSsA2RAErkEZRqOBfmr6/VkB85Jg8exnWSxT4PUO38KqgNcE36x1CK0GAtJ1THPGb0
OwNYUpLXpiIULuLy7LJ1tGIefZ8txieUEe+I5lNpVGhToCQAxl+Y23G16Q2yDQZRmyGQm+UzIl0a
N7zShxt0BsE004Ch/HJXMrqtgpfEixtaIVbhgsEGoVluzEPkIn6Lr7DPNZOhtyhx4kaeeUU473eV
momUFU9SChap6bp9Fjopds3d4uhkGDfkvbWp0x3ZxfKT9WpcnI1UlKnPoQ/Q8GAva31js3dvxu5P
/pLapuUUO5t9Y37SN/hTHjy7+jFHs+BUKCfofqaEkzuoVF2VXAXjirlCE2m15f0IMRXaUzIlepid
mIEMdTedwJAYACv+BP9qrgdKDD4bAyKWZWBcLEYjSavIjZSGG7g4u7WduTJXr+Frwqw414F1PNny
Ax52FBpnpEn9YK42njXFdE2YtzEAKKAJxyFr/gLyun1gUF9GgomfL0cHUglOtI2Q/lUKmxdTnXFj
iGwGylgDK13d0zLxzQzbmPEGvXL1S8zQDniWXWAiTuTrc7VZECngRfpWKRbJIemlquupPgpA+rf/
/2pgMEg44soMVRVq0WN7B7d2ngqJNHa3hdQrYFUqwtKL/xT3vzE/3VBxCJTv2vuJrnEkf8gGl2Lt
GlkfyRw/viBbCp/HrVnmygNrAytrAFqlD7CrBJtYlD2/mpiSTyS3WI24vmumZe3CXIeBU/14YfBI
TZk/F+Y76YjM2upebF3J/6jmRCWdiJNKwM7AL7jMtHQNCMx1RvzkIn83snqwLHFOvFZdVVFRsdKH
3WrmxkCuJAd3cOiR7X6xpOmqD5+/sHNfpgUJyn4kpg4fZTNojj+581BPJGvirT4eZ8B3LzJACGBj
Wyq+Qg+v+4XwAJXhQHIoew6pmfGHek7GL47irMwRE2ZM5cwzul5/dfEQ29XjAoX7ydAf9KFCBkun
AzdC3asxwrthRPMAwvpTWr4VbYtWgmhnEzHzSttRm01zrPUA2uG2WoCfQHNs5nrqGHoyYPlbYKVe
fiXTiqFRavoahxX5WKu0W2qjON4+xUKe1mDi6sVpGVsxjxfKLl3CUDFsYFzdWMRV9zW3HKcUBNI1
61gmiDiYCe4gAZd2mUPzhrjCOyQtbzKr+3umO+JKAphguFjuqmPGr+0h3kmRAKQU5ZjO3gdndtcM
KFqCopM3eMO1s7cjTz6p6F4LMF1oDzmDdxNbJkVTNGEdxB4H9pboNZwGKYIuoeAUuUnCuUQn2Svn
ZkRgpl3r9qO0Vhe3I7pafJMe/CsniCMreR6s0ylglVzShQtxqcOIUlHrHDTWkciEflIxUwr7D8dp
e3uz9uBuLn0kJASPfBD0OAeyxsgHXerZD4nePSMb0FMY/syybPj3kT12vKZ1FPxvL12SjDfbK9XX
lP6Y5gwmGNODuzjqTeZJcRrBQSOsg5A4d3yA/QG0aZKmE9SOMeEPW0dahKdIN/M2bNOmO04/huP6
1ym5JiwaGq7cDmfJWxTaxc96KqlP/+P2+2fToUtMGlUagYEl1Je097DUD9XxAcEqqSjjD48oaF5o
KM3FnFKHlUrzFwgR+O+39KVEK3kNCD8LDQD75JwKQaqs1bjxm0aIxwIyaAtLdhDAm28OBtI5V8+w
Hd6vmKzgbzxEQEnzJE8JPMg2PRQeYdrn5L8xlVS6paDlrWFEjbQsfU5+ir5+F7a63V652hGbPqa3
24hR2ij0UVf5FzDJ2sMyz6CXPLswIAPbrtby19BQpKKe0s5TvcOVbEg2lRZ+HuJesdPogfyrOL1y
yJY0YV0/UyXF/ddlNtApsJY/1ARMAPyxpMQwZ1z+czg0CPzo3rO2VX2eJZtpWwlSA+0EhIFwIYY9
GJ6+lRWBvel+d5FbWmj463YTKqf43sdYupAm8E1onHI2WFv8wCf8yuKf0BVkj/scOYJHyvsd9cNi
u21WWYkWh6enXAT0cKkWh9VmSNCftpcvUFHrrjuvXSnJhoCJXu9Kpv40kKFR3YQ4v2SDJkLyxNnn
IgdenRq7BNQc6VocHPrM25OuOlG82d+zLVHFGDKbjWP5ggI20KkswJ/yUqmuHmZOKLA7JScrJzBC
49BD7V7f++Ck3gtndXWi87SXMQCX8g5e0L9w2gR3g7+X73rOXjBZ304K1XuvpgLB/9TsPH97GJoQ
5KfvmhLkHSfStcklXJ7eNLEGhHpzzW656e6FvpYqQhOXhYt68TZRNtvLUB7bVXopU0zSmLCN6YkM
hkfA5mv19HNr/utrOHo0wdwg0UEb7lTyIKQWsAYts+En+klEShueKqwvuYZWelzXlDylMePAaVoX
5E2/+NcoRto4KNUQDTz31GFwnWXpwqO8BY5VqLqZwTEXNC26RAr3Vx5EEo7IOi3FIq7Je9RfiSXZ
f78TcLPuB/rNEgBfO3qfDQyYe7k9W80mv1uqxdjhSfZrcbWC6/syjxpZpZ6EYv7Fqb1kIAZeTdJa
foFXMYU34E3czutotekTloSCIa3n0OGWgp9YyXOlLIWRgTcNNF4bTmbgzsL0ylrVpn6+As10P3V+
Iw9J2EL5TjM7JsDjRAYbBIDiJ6fi2rIQJAsVVoUUJ/cipojSK8bBnnJcKugRDLrtTOP5YvLK20PB
p4bqE76e073D3SJnnLBh42ojznfHj+Ds70so1IokYGoBc9j3hVapshqNrACktBUIxGzL8buWkjuw
JmFsY6/SOTA06KlgIyCz0MdqS/A+v5LIkJ9YpPthVP2CN7Fdy55h26taWVxKiTpcDlMJRogt9AL2
BOdTgICn1h6R65GV5t/Tvm5fWX2qFAG0rKE9wztZtStbIC6Vr8uZsmhW3YKgHrtTiFdpPIgeDBlv
JtQ/s7RSsdW1CLyXBGRzPcB1sudFTwV87VkWgE8cmoRhuQ0m1ioaEeIleOnYsNZbMBDKS9WJI8vS
OrgtNngQduCCQACcB8BmiRoyZdep3jB3yS8xLrqp9fzLSjJsHfdJbY1VFBBoLyFHHczNvrhhjOeS
ZWCrPtC5wpBh+RZcjgLWc6w9aROBY2IuWTZuQGD0uj86TUqMPnrHzoAzqJyD01OLzHl/zGspHeWx
5T8RpdX9UmWOsQYdmu5YMbB5UbtkdIcfOmHxCNN8kdb5XjUvXUF033bjJcveEAh7/7GI9N71PPE6
MZzUBKFCWQ40blaegOpQTFwxZ464NsBWMRQYbt8AJ90rk7/tw4VPgIk5VPNjzALJ8AC8PRHUrtfx
V1JbX9VlbWFyp0DN28tkAeABRujkdL+E/F7EVSYPZ3AQDaLiB5a28nixTYVnfbD6d23QsDmNlqaS
oFYQ4vjOhdf+kNxZssVAghYIawM2/7ii5vDx9YBAk5JiEoewLnt55a5p0h5OLqlBK+G1+HyGntE3
hASBEd6SQkBOsAkHuaGuKLPg3SHb4E6PptMcDkVXXDVpkqHQDrpYBwEHuatf6STslBijwUQiNMK8
oyQvncOb8fqriv3R7iPjczqiOsWK+juMHTx8dtWonkOigwLOorLK7cgwT8z6INT5ebgMt/RzrK/6
i5yaRTpWlAHTL0tx3dHHl89Xr7cBmFIzk+bDjWr8yzRDfUKtS4Uj0ZtQWAlFVj7Hds2IqyCV5Jc+
i9lAnwlGANCKVm8yHjBoP9Isl6x70RazoxM2dz0ph3dEnym6OQCw598wKwIWAjWNUDDg3OG4AKcD
8TxGgjv8weW7awRIePzJEvSQ3Ui8kgdYhex2Jsc2ENYcjEAclzE2fGSwi5ZElptfnRgeH4ULupxI
hQnuhYO7uatyRZIm8VhOF1azwOH0ejNWcXm8pV//zBH+nBXC6u3vGcG5NjpDfStMj5eDct4cvkeG
24a9XoqCZsenABCQfMjon4eJt43vhuslY/KTn8TdSJpmGoQ0VBCF6zngJ9EPWAxI7kM3yROVEBbQ
RLsxhT+57DGRNurRWtTKH6rodB1MbqyX4SMC4hTXbcpLrSgx2AN816r3Ia9DjRA87wYdhdY3d8mv
vuOG1CdDHZeR4u0pxbRlqZas1H9AOY33GEr08C5y0sN2o+qyCc30vUf6zU9ZMzsFBv+1h6+6R5kb
yvuVyEezvcdHQdStOZGpXmGhmq3ySLrnEw8UCiWn+XFIqiAwA7cSvZ/CETQVPuMxkxH1X3/EAMg/
vku+/vLZYlInI/4fOFD/raJ6d4vI4xYkR15eBgPrlP+0KVWDHT5acLJZq/3Y000fI40wCR4+1Ngk
H6G6Fe6xJJrqSBO7WTAYtnp/qBW6nHv1JUct/kC6RaotyDatfJRSMuVkS+8wGCKFC/0by/JyFR+k
ej7xGHQQXmBaClRHpfBJ+GYjClPNMP8lrDeFA30We3Rp6p2A0f+JVpv3b4+UV/2hjngmNoy1i4im
x9N/K4UwaoKJLCxVIGNainauDjH209XW39K8av79OJiadgDqZEWbiaDTJCv4vrhYUPCGV+GdqAAa
kevmEbX0bwML1yynjGMglopJmb4/qDhfrwq/UBHVjRyGDEfi1Lixwe5/j4boX2pjEpg5FfBZokiJ
1XhrtT2WMfyklFh3OWjwtu+qj2rCK1FUEezXipSIjeMkA8tL5Vh0SwWF+Z9vZYbqtjriZK9zI5fM
b4U1p5zTyOxKX+3FQmC3o30FkuAkDtAYGpChsIoUpOjCwFY64Zlavyi/Av8lFw60MRr3D0yXACWC
OrgXB/3dklYF0dJ8ndxhIHqcdjeb9sjXShqTvHXu8CVepw00uduowJ9APPU2oQVh7kG0zq9mj7jm
DHpkgnkOwZbjBUq01lCsB7T41rUWDj06ak0lSNH8C/ENfupGSaURLDhbAokC7uTOmXYEPXn5HAQ9
RANzFaqqtAhlD/NjU4TE/mv1wUrStIGMuQtaHBNipXWzliApIOgNN4gQHTiOTLmPhbC+j2zB5dA6
s79RNyM22SSrHmQTU3J2NVKG9s0/Fnk5sAtYcodlSuCPoXMnXNe5qhe2jQPbQ7XCw9TNQug1uGWu
mcDYjsNB6Ctx/XEWlIvqrdNfr0g4R8gyQbsfQMdYLR0Og9Yd6Fbid700xZxBZv3EmGXuUi9VotJb
LFmD0tRawFYUh1+oiCIeQlLpOcXjAyTkV18eQQ5vdBKHiD2Xn566D7IfhNtvIhqlTtecUN0ZDsJD
rctbM9XboMKc1x/hgcNbV7YPKg4len2cskFe3zO7g0FaYCVoLtGoa7LICBN8g/fEMV1swwEOuciY
EQbWHmVhrabTGckxwxzze/1U/VsXZKhvCZ5JXvRfARe6AC69lcholToRWKSVj//IN8RZWp8o95nG
oqw8WQwIRmzPgHmeIQgt2CUDc6hRdvYOqa6LDlrRSB3xnP7v/nmOXLDF1KcpOEal1zDRBLMBiGgU
Fk6RCHLuqlVP8fdadMFQPCYxcEo+8CK6C6xHtQ29DY594/4SSazmYDaK3IWEMrRjzbhE4azPo3jO
DXhCfngwGof15taXQYcSqHQZAlu+xj9yI7tNCD699DJJPeQcGX6bd4TyQk8VwLd+rW7AvMuJsLOd
amtYYgr7dyNN6eBWHEI3eVmh6TWG345dGSz36xuBQUNWOZxSaTg3XmsdYvgzzrdpG8fjSO5NWNBX
ol+6DPN5wF3lNCxePbJxxyep9WYak7oKTs3tOhtDn/9bYs3pEao8n7dcfe5ioDb2DWrOsa2hi1NW
XzxrIVLltJFHDCJVrGp/s6Gb0SttsJRKgnuz6ds6e1nuYUVzioiovDDmMmIKKSiuE1QkSD3wcq5V
+dXzmwx5i32p3d+43CGiBZYnhspjK+W7QXlrLp7x+CQ+UBf94yj5TyuwS5FJd2Y88ArtUa+0LiBP
/sleevlkjPQv64uw1JGGRF3VpjgVlwm1EGZKIkktQyH/a3TyrWPmMO5TDsbO06JxggARQ2cbcy7N
Meb8EVDUYkVU7sBMx7k/uNHAvW1U1EmFrc3pItTXyoe5W531ZDlWeXyeyxoo9gZbZrSE9ZA8xkRz
XXl0KAdC+GsP0sdTzf4G7Pg0v2JtqpLKxzuFxRx3G9eKPV3zjPRlSXljydU4bees2G9lYS45m1TC
YoRCseupdOcCWgoagNNC2qU3DsHoRi+vPB3eyCYYXZszT9yR/fp0VYTLbyN9x13M8q5zW75eVxB9
DJ+IcQBjQ+spbFcljsYOLkQqJvGE8Bbs4EE0+v6pOGGZnLbKxAh4YPuZQnDxzx5uDXCd6tG3ECB7
f3WwV6Kwlsr/Z3V02y59pmRgGMdm0+02+L2IKfvXvtjuMjLfLyx51TYjfeC07GXySifAQ33/TenN
wq3fMKdOf9UXkg6vq0Dh+dXffr1Dp8g3Pieyk6hOUASmXAkuTv+znzSh0FsF2lmUTH1VTrnpTaL1
olugYdpZwN6C4Rn1h2K6EYf9qtM922XOk9ps9/Ih5WFZf+KwrSXYTcJIOnR8vnEm8gLJEj2u55J5
9tSu5rtF7WyhSju9mmsYyVpywjh76H4ISOV9i+CcF2ILfOL1XbJ7geM96zbFCdKJRcxPzu8reO+l
j6MphgiPCD9zPwjS6/uOlKJjCbooKWlriGAc79+YK3xY2d7qDPKMlZPs+gupkktKOYfoYVaYYAWU
DBuznh6v9ta4gSLhyWeAmlU0hxHnyyG+rUp9CRZFxDo/eeiO1ehsLrN7plXRXHjNMfjFs9o7xRWC
tH3nejTqU8dCZNo8mSAQYnydIAZzWj4ZgucVWJOo+QMv3+AEZhVcCbRzdsBe8ZTrx04x4riTNafr
meaXfuOrnL+lrVvwKdPh2kmlUR4UdLBt0Ff7k/N+NOILXByF7JX99wXniblCvM6pQrx4m+13XCPW
1MZSej2MH4XQivFH7uHXcLIzZizJfldA59XaoQqPKUii58vF+LWu12nlS2wRaaSvEpIWB9gdKTw1
8XROJ63SwCoBDBO3S/RaePCUll7fWdQzFZxE8XpcWum46ZAuOhHKQnwYH2jK6PPB+YNJSvZAMqWQ
RtkNu77+Ra0Pk5zdI01HK1BBa3Sfz8KSEE0tucDIg6CMP5MLoBSUtvlTD8lbYAy0GJp+TnI1NusH
7efi082LIkeVYRJVZEba+0Jj7X50IOkUW2UTTRDyugSx4xSe0DoCjtG6+iozCTAfsyZM4vdhXl+Y
6h5ME/Foryrjj0nZJIdZOEf3hW5filC1XnUFcp3xazKAdrDwJvL6XSnD/YtrLhgkQ+eLQz8gdnjF
CaAMOU1BoQUpjNALAX7NUEEkQg83aY8LaOLXsD9fSuP4jtFPGCThgAp0SOTciVAYbHEhDxg74stf
dF+TTTlsTwP00bsCEqv2fiDmyCTpqq0X1UGTomnoBtXgKJ4dXeAR7Nn1FXjNnz2JpeKcemKC/9cw
hQ5PcmhJl/LJ7pz49GYDj/0li4llPvar78q1Kbv1pluKnquXnsUYccZ/nnY1eh4XES+G5JKJthwx
JygR9ECHvuWudiNLOSDldGa1GoazM2/SDRjuWCzJCkMpTy92HYey7rTwVj77GkOqxyCIHHdP0Y4E
Q03RwsKugfXzZKvf+5mNTTCY9fN3Oi7e2zoV2buny4Xjy3RpO+99PrmhAGPyPUo4xFo8cEQiTQBV
kmwtSWuWstqeTsans24im1jqTrV4k4DHH2bDITCbE/s7KVv1zJbqGjOKyVH+yNOq+2YVtaJ4U0tK
iovvGc5bDF8Yo02Cr6zqtUkBLPXPw1FDudq8oW6vK2mNslmvH+PGgTjpa6JtD6RRg6WcYJSHW+qw
xtK3pT8u1RtrjDWk5gvMyiGEDWot42r2ln2NWXfQHmrOyV7hIBJ2nlwJPfW8wC9m9h7bzjbpfe5z
/g/aLUWmecLdEXn4cLdZ3+D2Jvh6zNIOat/MvKB+q/VoKTcosj6GC5nOjum9s+7tN6U54yjAou3l
zi91JTZKWoKjGGJQeQ4PqxucovwV72tXZnDllMNuODk4C9l78MPoP9LUUv42hQa/cZXwEyL0gpeC
nWrgm+lrPWYxI3mviuIbjbLOEJdivZrsYRVud/X8IW4kzPBnrrE9W5qITx3+U99VzUIHTlU6iDeF
R1fIu2JRGVPGoBSE+WVZutXTrH/cJkA6Hb9/YKMM2KbUpyMPQkZVh+M8Z7qp4yWLLE94pYWHYlxG
UKinjQQPNfMiZkuql42LeKas3lnp5FjuIUM0p85IPON3KdgzlM/Q59j2gDB6J+QiqbUOtgCGcAId
vB58VzIjJdr2UCwbLXCTOUFHBSlgJqDkhCzElfHBebNqkdMaSMD1qLtNOa+91lOC2kkZobcydmlz
Wm9E2uJOABqyE5XC8Obtwk+6VO/q+57pjDsZ36jY9Nz8r/Kgy5afeUxFbME9sVMY4CaZEKm4DgIP
dExDJQorQoJs3uKC/5RUcwKPnOoL7Kpq+Wwahvh8w7pr9FeV0YOsuseZN5Jn5Tw8wEadJGZJldLc
6kyvRFteSZ/0W4u3dcBxB/3Mnc302aF5BLwQYHHBtQgO2BgzjkHiX2clKpDecb6tHbj4VqgGYCfa
5NpdOweLDYzb1uHTHFiKn/BF1+dp3oZIJUk0CMFHha06o/jsZmyqGlmrbHIHrxpEyCYE7LJB0Sho
V+Kcne9bKndXnYxWglacAV6UTEV4GpHWXC3CCAJSI5Az9vkRDUZGcz8OQlpbY5lZ2ah07oh36giV
RjUAdKh2cDq8hKX2y23RCKOrepayq5n2DLZjcaS+TwwFkPcpPXMWO73C16ZLvkdek3i4QhlRjx7h
q9uteJXQSgcRX0+MnuYMHRh1EPZVebNCjfb1NhLZg68bE3BTfEpIVAWuBRlWY6zjI9BDehBPOi1x
tjhoAi94NVVdU9qSjGvVN7mzMi++2QfLmR4OtnOo4oAgmL05qfAnHKc/r8OHdXCx3dl7jBHLl6cr
Rs3rbnNpUw0f9sUnUTNGNdRaN+ergM+HP3vccyfIOYewvQXYos3HlPPkfG27fJeVcV6HxZ2GVh0x
AuVNEI+AsXb+ZlyNbpJKXyRjKzYqK6JzAkbCmfSFYDmxGFFWFMC2gKV0tkRHTwtVMMVV0iLawNGg
7/hi8RrCbNELrq45oHMWtgvZ7wpAWoK5wV2+zeBRcr+nzkB/kbRzV3TIh2oHgE7JgnIVk4YVzB1U
/C4rrFK+6A2z0Lck0Yf5/Vm8QPnnUJ5pNCDw9Xiz5uXEMzyEE4a731OrtZJjjHBteXgmlhfzcYWs
nPRCacJB/WcSi8m6DO57x0eaife3grjAsPtgpT5FOM4UqUX2PZ7CVmwz+YTmT558UBp1cUWU2B/a
7IoBoesddvEt6aeiVsejw878E6jNpL/gdfjtifVx6+xiQJE2TPv96UPSjtAivhXLgkZs/vhQ15+z
WBoRgBQ3V94w9u+wGgc57TZWrMr6ELDk0n7Moxu/k2wRgDtHNhdsQb8NB4TZug40S/71wg5FWK1Q
q9tNGzN+kPk1tdxOoLca6wirDVXU0aF9KuGnVAjlJb+DWPEOzVFIMd0WP3Yo2wpfl+7uyTgrKeUT
z8gn0hAeH+iIgTkqKfRD8lgTQDqWklao3MyURcMQ9yBmUcFjRn4DKxQ8tVgNnHLk4G0FdG5SrVO6
aTxJf0hrZziyAZx5PriIAWcPA1TgYPyiXIs5jSsqQonOvRAtYxdL5yaOZ/sgCrfCAfnhQaWvGszX
c+UzSV160gLwrtQC2UxmnVjTEQ3qhcPpD6Rn9OKjDoP9tS0MPWijmaer/NvpDidSUOnqyfwwmg0/
SW79d0hUceRRM2oGli6TwpIu4vRfcGcA6AidfTrhoVrCweVKBW8KSwDzwNJyK34aSPmpUPdsiyRc
Q8znEilPGZWduY0fUNOA8CV94WaxZz2on/0h6TpaCZjVFAabn9p8jgLF0wgFHWav6S2JGYEHheWh
Ez+ryLmzJzmFwiZlUAuF9REoshGX+ixlfo+RdTV8MmyA3pY9xjtlNEsMzo9uK0Gw4FjNiK4mpmeW
iVoV45YjuS8uhzIzJawGNBg0FDKOp4XhCzNgUphJ3f34F0s9Ah4cDZs8J2L99V9YqajzIr6BuzCz
7Byi60G4ecLV+7ArqJ9cId4ZmTb90Ikl0hD3O1R5CT+K/qOv+2tVPZ+Jwch0Wnv2Scv/WldFUbTb
4QE3LC4yzRMHXYoLX3t6T1beBiTEkI/bV2lxUKY1LZvIkGhQ7kykm1QRzbfvdMSiii/UD4xk+jCN
Mdq8fgDr3xvmB5ncGgPkeAMzzFpuPtff0ftlcLWbl+ZodnFD/7J7ArjukNTZvxxJZ0gJugrm0ljy
PMoLbosQBRIYL0AaUMAKY/SFhGuYf3CsrS+cpiIxhZcHjyefDekuyA0t8xXplDIicEkWVRE5sAnG
Y6F/4asIh/Pl/9hzS/nmuFrQ37pENviALTM7MwOd2GqrnlJwgFM+jFfJ/NSIKjCp0s4COZ2MlIzH
m6Ge4N55pmfB6Tb7OpVZd3yIrXw5ghOtf3jmistVOrcEQaGd2KclUQFOFWa87KaZEaPiSyM3yqNZ
B4ifZPTMRJ2B3k7z869CU75NAyrsIanzH+cDtFjZEJSKKErSoSudZuhfbf9ZMovt1lQlNxsbDUZh
l7Xh35ZRlyuyNYK+PgBrWeyZY8LZbyaW/lHSCVEnF13s4Uh1GGYUpv/fkaXWZdUGWo2VlV+7hP/X
n/X/aFoNyjrdkfrHs1yHDG3Pwp+KyltjOTWjk5btZinJ5zffQzY5NI4cV9bldJo4LhiXJqBpC66a
5n+sggxjd8MfZIe9O+A23cC+tJOXUS/qS2lJwmSFM4DuPGgw2Darjc3stMhbKEivKaJQZt+GerrT
yL8Vmh1cpFYhAR+IJiKvbhyPKPn7WRIf6Nt/jCYSWdRriRtdeZMvVkGw9yi+fRKnIsQX16lHS8P/
c2IP/HH0lzyG/Ferh2Do8+HeCL5F1SGQTS2u4Nwq+HUjHrZcnxUH3cDAM25QpsszZaq0I3M2xzGb
85O7NUEsghF0uIUHeZgKH8KysQGs9DwU68W1kZE7Ww8zd/KcF/d+zwl+KImw7ov0f+aTSxDUS2mP
92v7eKmYvlp80gJp+cm4gTgnkKBzOAmNteIj/sUJ60gJ5A/3KXMamI5nZSwSQtSIKr7f9/z5dux7
3N6CB5tdG3ypvbgdO15Wr6j1opHG/KVK3MlsyN9O6QMSqTotQU3QJxBPhr5r9ErRIJ3wmGr7fOa7
r3J9msLe7tdRbkARPc5jiYZwF9h03VN6e7dTYiY1mihDDn/qIpN1amF2SM24pD0HnNyhzbsOHRN6
pDEq6VpozYSkWnfh6r/EIZ2Ryaz3EW3uMb3eoTnscNlygYrkZArNQKu8Xy18fEhjLUeTLGJk+y/c
+gNwWEtR4MW6ZJ+AHdhvLEOoHhacvdFuJFEWhbxsD7u58hBKUOC8j+KTY5i1osY5mCA6TEfcC5SZ
TvjkznqNKRbAqHoYQsVWUD2fyFN0xJSSu4ynWM0pCA6qp6hIY7vUKs/Q1KBR/ROLRhRWRgZQfynY
HzW5koh6I2lk+FpfAAONKlQdK8z/J+xPxK9U/7EAsuDVW+poGk3OgMOEfBwmxWfCc5RoRnh9MQRh
4cbLzWaKMzPDXuv28f2S2lImYrGYPobcb92kru9Vyw9z4RHlFJuhtAirimFGuJH5IbtVgg8dYfqH
r2KV/zfd711Rzuv8hsdPPncFzHtbzvufIMikLcGIAN3Q4gT+cX+ciRwm5p9GYIEnutDqwo2HhYOj
MA5Csu5P37mhQARUX3+glw6qdutqk0losiDgmoKVedKgW+ryw7A5ekn7CyMrUKYDm/Npj4B4i0hH
EnlJJwdXslWcQUyqAexnFt8ziFAqemMDi85v++BjHxOeb4I/P9KoHS4ZfcWadVcV4b4ZFzJ/0MBz
ZeBY8e4mXXNZ+NZiP8Ff2bJKoJzJ2p3DUBBBFQdz//XxlJyCr1hxuHLkgg7uhjN0DuUSr+OnLJD0
IrPex8jOAAl0qLT79UJQXVHOlWDyOtaeMsLww4k99d7w5SAAe5lReQZgHf2OUsTTzxu3SLp11UuJ
Q4J7xT6WLT3uaVJlSaUDwR9+UuijIguHAHLZo8uqrEQl15TszAjZg/IlrqQMfqMU76bU/fPWmzJS
ntfmxBJzvrrnvvSh2NsmgkEITdi0+udJDC2G3hOPnRo97PViTFdDftdUvzmrlLF8CmKEff8c4pB+
xvtuRPe1uexrnWlKVs/YaRyjfo4wnGLL4+8MgVobPeX/r5UzXx686ojTjYK6/R9V6KyEnej6ERBL
mSy2a9kMCMEq14k8MuZB4yuX50zgMM7Stea2rm8qil1zf7fq+Bbo/rCm0IWW2MCnZpUUqym9Zv/3
KN8XoqGPLUSn4aLZ0KdCt8uLhIlCqwYT05ZhsEN9NRyjLecA2RhTKE/mjNOuQ1wuP9d+klIWQHJA
+190yptaQZIiJKJmjsygQNoijashXDAUCfv206ITARhIOETvSTR5oUjh9sV65HDqMB9XW2rNjMZD
zDq7oNRZPTJOkLRAPLtwwpcMD/al1pvrdKLBAsChtVqDKY5ANmXueymaNrS3GIbPuOIMiAYI6U5i
37/H5WSn81ogNFESKsLvgJ0colSVMJs/NA6nD3ZYnxsw4W6ZBT2p+pNFnsNmVdwAAyJEI81VorI6
qqVd0nXMIp90wrCcx1q70byKn8XTbnD7O4s7aYjjAEMPlst/Y7TSTmy1kUEJHNCYzbM0sxFmsy9g
bfb6mlxTHaFozHjOxvCuMCy500EWs2niXo0lEUPoxxKelb3xVUF4W84b5Jc9JBuUfr4QmtRch1pf
tStcnkJkMuNwYx4j2x/KVP5Zm2QEAgbXpWOMIc4OKigqXmJpzAc/qhiVzgG0c/fsdvcnuSY0yW2K
WEzCBUH3+PJr7+svjhGEUU82H2ZPcX2dJPQlv8ZPU+qL3upJVWnCJbmy3Hj96T5/hskVJ6ClCr/l
d3J6exBDIQade8i0wegvbIbWAaPLuTjal69x7ctdPYmW+6JJxOkgDtvkPxctmm8SQEILTIsbg/g3
3El9Y7aKWs6ty5j3smdpFtP+E/BxVYVliKcNlTsrtz+4GcL5Gpz48nWLtIVBWFGO6HdV0BGant7r
KxCLcE/POiuVbPLmtYev+BQ84GiRLr1Ld7J3WNzki/+DPbHa9xpNZXhow3EoViwaDgQJUNpS3t6D
RI9J52J33t4jNN1mbXX/gHlFng7P7qYGdPkw5OxJqBUCiPSGSfaxnA+78ins9aiQznKQqludNUCg
B4IU7ORYlyllxZxVF+3/e4ywk5L2I+ULWU+oq6jvIGPsx8wVE8NTZ9A+Yj5bZjUQe79yDcRxWnzF
IgTdSuf2KK0WxInacemqbwiU8kNYzh+nKBaYNp3/4CEwKSiDrN2+63RyhFhMeWBvIgSXyvXW5QHd
eTZS/SIshlwL4o9YoY9xZkbUeDumAhVLZsbwHx5k8VtcgUY+2ws0ui6WMM1d9X5uqxD17r9r3zHr
SbLtzhFti/xJhD/fjfShwtJenK76kJyfrOBfrj5HaDOusPhBcScbl9d2J8ACSH8cJzqlRvrMeSwM
yyK/OQSY6+KsuNCiiwIIVteVPVlCbQVvy0uk1V7ADnT+R0v+hktL53ogi4QaP2gfnTpj77oNhliI
5xt6aSoZO/RCKPuyrk8qpDH4n9k3OYWLlQwjjB9l+yTzpSsWJpAsHtMEZGNPdhknZhJlbSha+asU
OgQ+UAmXWTRqMvfnr5Hvi/6gdS8M/cgMFzXe3gnw//QBMMveT+edXFCgpXi4P85q6ul+jhq1F+n1
rEpQTkQx36M6/VcRdj2nfhJZCUrwYX4oCQUs8kmCYVeAw25gbTznB6p3GJlnRc7dfBsLHg5PlGr5
emCH+vy4h+mJenHbPZ9E6B342QWJwQDIzBcstoSQ0wc0OvJO3ICsm3JxtSjCLh8yxtqa2+xQMMRe
yAqi7zGvS9tvC2MAexNWWNFWMWBtnkAlGRyfUux8maZ6Yl1OJtTFCbq24EpxbSKMLszt2uuVSFMh
X/bMIg7X9olckyALbsYrP8ztVWVzXVeczi+QFHeq5BwK80YowVRrwLmRVqeHgoF7TqwGrzVkLAPC
Y/YXydYtDQQI2XYjKY6hA1GsOx6dAqCGRlIPcofgDj3/4qDt4BolYEiDOHsrBQ8qUi+ticd/Zh6n
oslO8RoZ2rPzCC0EjVK2Tn+EhYObiPtxbPvEDdpDAF0te1vlgGCbhvR5vWE3y5AWOTKWJ1EnZK6F
/4uyDVa/CixN6vXX6mFIA4IK0jd0ZtcFUJvNS5oPzfvIIiyP1V72fQQDyJf5WvCPFEn7GeVN6nhI
OUWApsyNv8vEfZ9LROzGSD0njyfFM0usDUFOwSn+3OciBSwSVfkFjFk8sXQbIX2GhlLiA/YWsy8C
u5Sf7N8LF0W4roreU4i/iSkZwSsCPSi9WjgJoS0PcoMYsvdMdFvbn8sMIzvYtdLWjPdHiUPMiVC8
rgRddXEFIJWWrNaGCBCfJVVzxRcx+n4m3PPkGvA+ll536ti0tV9ApKhKYLRmOD/AtMgIxuHGIVAX
+KRlMx6Ot0VjfMiegDgJiWf5b2lpfF9p4MkI7DnIoFoR1AMdgs8myBo0yV3HDOsUgJ76JIWy/WDc
Cswx2OxX6tFSqVjy2OMTFpNZfeSUawneV/BT2V86JUQphG+BXB8Z9KqNYOcBFL5wb8l5wmXWmOox
esXpiHjWkpEYpg4t6x/SECLKiMgikxnirWCdxwSCXBV8QcAqhgJjGP8ANm5aO0ZrxHIDZe3hJKfs
AMriITqBcPLnbXoIs6HGZlCZPZmhtDpqcFA5oLzWYZwKpycg983iGOTOi37gXaRJmWmEorPKbULn
HJZ/1cPMQS9zGrXvXjdNGxRfRhMx38nCM87jFxAYSpHCQZ3LjVUizoAPWdnDuOjcm75fRjPtFNu2
S0I9YIdgLWOho2NfTb05YC7SjH/D9wH2ZZ9h8WMV080GXCDRgO75LPeGzz0sscWJj7jE7E+j3Eoj
nlo3L5ub11fsjMDlZ4DXlJOD3kCzxDsqc7Y72tgu5FC/pFxPPNNg/XIJ9rLKNHQDmyti8Uyq+tNd
q6zzr35a2J86nYKMPhxiD+b7RvA8fpU/WR1N8g6cI+E9r4Ei8t/qxTP5rSCM9N4dK7ETikWC2ZJV
PQtwPOEk4M43Gh/DSD6ZD8FOO2g8BlauBGfDFAeA/IQzDRjxMmgRmiUwFGuslQEN9rCzI41+oZoz
vN54UIaGBJWdZZwSBt/fus14bb5BFWW4yEFblkSbMRxH1DuIgwf9QoNsAN6Ojv1yTXYpfn2PzElZ
4tb3oeafHT0m/2oUS1LzWHw3GUNLwWa9GvyUkOgzV+lC+LoAhP44QFhg+sQDYokAc8ieRqggxdIy
rdXJLtS81fnLDHqagNC+fANJXH2XIMDKxCif/DLzrHUPLJAEVSWOzn5VCXiv8XfGqYMxdhhnAkBc
K3S07ek11UlyVDkzKR+eRz8cIGzpcpKo9zbA1YvOXD38lISvA6Go2j8taIEkaAf/6zzooaH0ciYR
jxJhWs12sy0pMHQvXrobrA843e98JbcQ8PEUKERsqbroyHFGtzge1Q5gNuI8x80Ybhe6SCMBYelz
r6Mq+goATku193apmH6EfuITTT/qHzo2GXDyReY6zXYGrm3X42jIemANbm7yGXgip8yqo4q+nQAQ
cg1b3DGDu3w8qiIgG2hcihJCq8bxOF40Z4d2JhOxWMZaGt+nrMAC8nGmgVoqpoFdJ951fJ2f1beU
eZ1L7OwTFNKiQ8mHQ8obO4zTz/eWwItT+UqU4ULSCLSMCw11OY/ak/e202lKW8gh1hTEswbsR6Z4
bN/m7142r4h5CafcfxK5GIs/PtT1jsJ2KJIeAngc+6Jktt7FRuOSBE+EQNrdggUduS1QbuDUcKEz
sHMpYSanO8QCjy0H4AjYWNIexZOsn+u4kuwBfNPK/Fex5DxsBX287B0pJK2WZxTF8y1e42ZvCMiB
nar4sfGQZcQEecheYv0h1Fhcmqjkt5tCNLJf2IWNDxwGz4WwCuDPVNs0kuBsjVKuXdy4RJl4xyY6
gTH2wDqaNfmXZ6cP2+FPu/5SikWFapspcaNvv0r+6SJeHJb8apjt6SWJ1lC1oty0g7/cNzIyTiyq
VQTcvkVZnIWpMS8lGSsVIl/37qzezVh665OIPoz6z6CwQUyytiVgI916FcbJCMlxuWqx4PTiPYVW
50M5smr9W8ozMXPciVflsrMCDh4utIPewl2VPxiJ0+QEkhGnOs2jq/i1Rrd2Ec8No9vurevWWELu
bSy72sA4Oyhe1i7iEf8PEMTUXyM5xwU5f1SdvHqtg8Z69lNgdyoPLL+ewrrv7nY77sJ8wsm2m5po
8rmKkwtbuF6e64LNxY9hEgvZCJHiobquSv6snjLHGTyzBXPCqtuaCUhOOCHgfDTTXXtNhdBwKDDa
YOjPercTysd03tLHLlKmLUHq+xgkDVFlzHMoPP9sojkOc7jr1yvrXG9f9DsrNdsre7uRd3pDWNt7
xdCz8igPg8523OwbXHW2YTVKEacLdFfd9ECTJDZ+NCuKMBXwFacCTpxvfJfaGxGUqIy00QUvmXfT
9QjnhgwzmS4o8SQx8taO0lsvp6SOwvDJr0oxHiW2dFL47CRgKW9n9pJsfRycJwl170ci0CJoZHK+
F7V9//wwU695nW7PzovA+F7bck2e8zJuy5sJTa7RH80n+JjHxKZvra9iqXRpgOL5t0130DuOy+sE
rZPfL/XgJhlopYnu73pYFO+DmVl+pWH78v6UU8oDr2jDKBc4gU0FlkTrdMkvTZeN29j3r09sfxLO
/Ix58ejlXVJiUntgGgpto13OpqIXL3tiYUHWJrqQpBrIFOU48JUPVGAjoENS2y3hS+4Tyibz7xUk
TtVxDzo8BqOlA3XBP7OIlcHehUK1HTl/kI7cT/RUeJqE4ixvw+qRyNUJbxS8XIVJcdr5I1CzkGCN
cbTPO+Tu4HyC1mmXslsDJliW/dxfMaPpbzGgyetkxdPr+P9f5NmFFl4rn9/ON/ihGCrvdXpFJ/kV
dbpmbEf9os8SGwhkYmM/XuZ4UwXwWj8AFgGEz2skdVMOeNJ0l76HRyul9TOZyZUZCNo8gykEiape
SxhnEGcqUYbInos9OW/KLnbkpmM+69JjA9/H9bMwfoc89bLQuJ4Lt38LBtoBy/5bXjEVQ+aMLVOD
Pg8A7ImcspHXgKYGGCN7ftWjLQrgXdSkSnMPft4K5s5GsSPitjqXqnOTo6nKG0nuwCj79pvhddO1
KTAdryHfjz/8oYBJR2vTdHVnHCqulAcbrQgBQR2+tXv9SL0h0/MnOkRbW4YJTHb0uioVbqNmvXh/
zIgc81ZiYMYXBU3juBzat4JluurgpwH4HNDNXkhA5ry/T7xfSwEFurTI06WWeGcVJ/zxYA13w9aK
LbIkTLoGXl48C5zqZ63Ee6WGvTS8sKR8aj39EmtcjdV7VSAordqmG+Yg3yDmL0SpkLgsGGFLF1Q6
SpHFrwGuxGhul5leswHJoiIDkCYt+oo/k1jODlkjig5YUrleW4/Wo2ylncOy72+mzKzAjwaVFy6j
6WGGLW+6RIP9dMlhUbdhhnoWeAxinp6/HYLn4Pptz0vxBqkEsEUl2UdWRcIU3xJoL2Ek38hNZiOK
60Ov5YS00xkbKIOn5Gy7atS9UWqTO4t2nKNJdVprhg02FYkDU1VP6gEJkEtCrIPq9xMFh0Mdpvcu
cccnvwEB+uG4O0sjYJoMVnJ9FcNtUxTn9+AnTvfhuRVO4b2i2eiLnPOzINqZ98DUv8KfK1qRvvMv
yX2DS0bxnPbmvEgjAcFWCCdnwr9gPAcoyr9M5b/meb4NnUWSnJB3Nio7KpKBnBFRCnrj1sqNoXjC
pJxEQ49mHe4q3ndCqyPB9NnXp7gX8jkd+kbg8NdL8esG5do9LQJWCwU/n2JZVFuPXDb4Pnhr+325
mH2BsR1q0guvDivapCseZZJ/6hVhZXolf5gVrU91wDjTWAREeRt2o6AHGR/is7KvijqOXq338d9W
0aBl2khunTVSm9/VmmvytaGr5oNp9/VBoFGJabCbYcDY2QAnG4S9j2Ufz7ZIfydY81mC9ZdD91yh
7sTkynHulpWqeC3Iq0k5g9/msNef9320Fq8e5d7JA5X1doELFoOFLqw8M6+wDdAgz6vKa225PBc3
D/GH//yBDhY8KmL+X0OBUZJ75eLzuFwNSJMDBfwUa0SS4pdmb4p1Se2Ec7g4xX0YOX9yGyxtQMhG
MPfDR3omXuK9WY07xqlY38v0PoS9WEP8YrG8LCAbcAj+L4T1j8glmq1s1mRurFHDlmmrWQPUsY8s
e2A+a26bljyisQtMVG2I7wMH8k9HSxAkQ8F5A1FhmIKgZDGXCbGbPMtfbEQ6OvcAMNlN/BGGVkCL
/pc04NIpLshXSVbBvcQ2cTr34LSRq7OR+IHZ26+4fc79YpiZcBPVaR9L1BO+9jyfD3m9BW+8Zowv
ksMiDqASsruUBymaMH7KQM9xauKqOflzZiexSP6DFEHEUo4WVM35i4s7KoeNgjFznAG/Br5u2vKK
t1J3TPGGnUabrmUlJhwVjMMOkyx/4t6rhi2x52Rr/mKX0mt9uwntW9yXmidopG+kTzHzqEeaSqHA
AcOBGRRXAikMtZjz3bE11J0zRF8WazHO9hPoDlBikTTGmCvINw2ecn3q2L39aJpmXoxsmObmoh8N
FXNGxOUkyEAYeNxc7jQMJHwFSlCRJ7g+BMU321Jhn9cxCk1y/HlP6S/OwcBEqG5zb2P1e5/KmQrm
uUauvQRcDue6Pc+C+xW9SS+zQVWnBsDRDf+XnBPJkYCxO81iNOQW3VsI20j9WXykGrPS6O5mNeXb
aO6g+Rro7OOGOmLYrf5goATW0Vlnr7jNP7YS+Jz7MfaymDLvnIT+H3eh3sHbO884SEEYbL/rJUQw
boER/o29mzYbqLWFWx1mII0ARIap+iJCo2Y1W5ZCite9WRToFemdXJvJk+L036YlWrz2yJOnKIaZ
K9ONe0j7+SPuc5J1j7BM35GiJGQG6Pae7H+3ygM7xEoazdr0U4PINSbR++IhGSJIG2eStQ7TT1Ib
Z5bAIoTEOCLQtwkMid6XRXavlAc81uE8Soaj+tA164Q6F5IoyfCpH8qKsb+vxdfeQ9wnKXdRVT+d
N9IxhNXiDYejMITeHpd2mU3NhoEZr4alK9g92pFFlnL12G25nuMrkAWZ1ZdnN6lmyngeuU8rkNF3
TEswrIQ8j7+Uv+K2BJ2r78M3ugw6WOJyD0xb23XyFNqsk/3f6NcupLrBHowE/pGNDMW86tHU2Oy3
Ha3HLQNnPNpZAjmJiyYC+AyAffaePD2beV66vXCUY3xgVB2eg6pYGXR+ImjNHszYt/IKBzdZT2mj
H4xTl9FLw5LPYOTpG5Fx05RiqTMEc7w/RNLuRnAuUWsIDE1Ro+r/QgT8uAq/EJ5/2LFF/hqg7Kt+
MOfZXup8Ol/e9cOerCSY9V7k2XYuOTIPPvVKK0v4HZE0+zuHSoUxS9ITa+jI6zPpbY/hyvO27FO3
KuH7veq/aIPL4PhtzAKXslW5h8Y8oacZXFhrOWhiR+aA0a8eHxbLxLIcfzf8jsfnbfja5Y7nBmbp
d39Zgry3aPSeacc646UWJinhpe1PXoljT49nyVEz6fOvaVn9cm2nFCj1mhInkLgACr1LrPe6kScg
ATi1KpjPUfgNx5lrEZ2aE9ZVgu1HOgo6tIbAiQ8jYrQYG/jNGiZATvlfXMyrW9uJY1yP29UKxgAg
T8u5nW+RAPWSkHRZSxRoHjteUD5ttt1AJy7y/AC+D+C/m8jRQ/bjXaVZcnrlPEtRu6ZVjTvo2eKM
bzBpiaJyGHnoncBZf1y9LHaoPlmKB8SJVPOogra02uK+HltH8M2glCEfrYwjhu0/05uWTmP3uBbq
tZN+9NvwlFQ/vsCG32xHW+4PFEg/yvcWr+uhDw3vgttOFnA0qWjYOVbFzNXsmnKLDh95PgZPJbqf
SjXGbY4YYxtnS0MyjX0xUg1nawvnrUTTtUm+DpiwpfEAkKtewV0A1CfHNEu7ds3WufSztiGDlpJS
+yyrs5Sc+53CtWtxCBFrbVgV9sIZ0w0sZGtiHlqL5GxrX0PzE3uzfJM/YXzjBFyjrH1sGLurS1Yc
NeJkR0rT2Ik9YsqaOOPrdAziWJaGohf5wLFtdqa+A4EeQS725ZhsI/oc845/np02uVCHFOg1r2dH
SKybIfh6lPsCjuh7Ss+QA0ODXobrM/Ol2w+qdxv5t2BBT+becch9oPII160/LSozR3Zff1CrTmo0
dmq2I4Oi0bBWYHJi8FodqW0Oe0wuREWxz10XYFXb/Odgus7J+476dsX6cyycsFPHgd9oocOnYSZ3
Er2c9ux8nXyAcaPmnF9mtLIFhsDMfpLSPxBMD7GPwUFFvjr0Ne9rF/EJqADfXfqI/SmEI6ocht6q
4icXN2whJ0/76+BgtoOq0nN5kIawg3MFS7YI5Hqqe0ILV65WpBCAv+I8Mu5M5P9IX4CVAF8QhezR
AlEAy16MuELm96gES753QSAYazfepMxJLRcPzI7VLMFlF6A78lC8boMwmRbbVkCTkyrBVvELHyv6
780Z/FVTiWpjwlOBcS4Qb0vzUeIv/rkWEHKA1z+X4afOibSwRBdxJZZHTsjqpIxTGVz6JoH0Jk6B
dhMDsYE4tqVn9UuCkruESTDcjNMUnCwMaVKpiID9ptSzC+RCZ89KarGmyrTF2/7mSbqCHnQw9MU1
XyEMw8xGKGSwGeJOKHkUG83Jmv/JFZg11SosZ6Am6QDHHzOumb++WPzly93dSkEi3Q5HuGHJigvM
y+wSyUg4U/QQIcQlgsuwyh47aZphd7335JEVGO4admbsWCa0gtrrSK0bwFisy3Z8qWwzuZ25YPnC
vttkZ4pIGWCqtiT4bcBGB1MdzK7Kc4IBLF9qzXW5VcZgnRL/FYn5m73BIt6ghRNInkYNnLBzNN4D
qi+hNR1f6/84zCWgvK93tH3Wtt5i1r6kD/j6FJzi5wTR6rAXG3m+JRDJF1b8bcua9uhIb/6h57sW
i9f+NtHLxI5t4MUeXmTOJ0HwZ6KdUVUa2SWhRmgQInbT9qHG86cN5FUhQD0XG82tXmOTlAk3IbrQ
tRELENSn34dT90PZ++rsIzQcu4rtiOc8Ox77VYQvpmw3sqCSq6mCX7ijcn9bsKFtV8mMbcL6G6wD
IjSmMOLZfBOsPJsk+SIsI1ydKo40QSFi3e55+UFEP2umla+IqJcSH1Yy9VoOgh9EiAIP12Wqt0kI
2v3IwLCX7CI3GJ64b+K6QSU7Tom7XbAnIkuTGmUflTl4hECzLTLR55sYqyqr293NcI9TWiA6DyVu
avoIrwXKGOYbnvB/Yfc3hk4HoUjSFhcB+so1ylwwmMDDAnnxhzRvjhMWT1IZplqPi3qPAHurkUN3
mTIHkQVtvf5rwbJWj6Qs8ZNxzmhBWudkVyri7KMwGA+wQeZtQcB/kjDDjMOM51Est4yndiZhxvCV
prQ3n2dadOYDNwost+d5AJMvQg/XP35h95TAJVAp4BmOTzNRx3V7UQSitbbFwM+1iyT/8juWzMrn
iQJvtjq/0ewypr3V6FASxiIMsR2quFkCejmO5O4foPk1Yn6vfyJUOZlMmfQFntHgKrs8rPzkAj9f
BEwAeQOA0BdsozYcBHw5292CnUtVymUmmGMmBjxWhrE02GgFFgSuk13S83NG45jWq9BHWFDONNWE
DUc/3KfMU2HeE2hFtUgahLx+zR5p2r4hYXh5On4PHAQgmpalUUwgBX7ELZCADJKSjIMYgsMSrZW4
7eKkZ8d5j+zSFvcls57ar3/O0LhsG9ly8hkNjXnf+wX7nrdXn/06VYcwb1ud9om7aKJM+2YL3i1F
AoCS3K7I+36OiFV/of1K4wZ04+VG6lcSuPxxryOZ6cG8Z6aFI2kVS/G8KilAnx3pPnvLs/7avzuW
/ecDbNI5IdJXKxHv4KDKW5s34/aRJeZ2jg/H1oA0M8zvWYQ0nMWeeCK0yM+i9or4g/e399o/kyzl
Zf7tkWjU+QoKPbUSxK3fK7Kwx+mFfCCFv+S/hRjS9C8kPtbilpvdY2lqGLzxfSZibvaRz4dBb6sI
K/o1rO2MgdtsnlpROkxdhKg7s5Ka9tavV6g6JNQ9NQ5pqP5vAHtG5VT9a7CUSHokIIiWleAF/C7T
gGigUb4b+sdBj1LOkeuhuzDvPhUVjjdHxM0hprFpU6mzAu/KplBShsqiBr8iNAxxcaqXTuli6YMA
z/AJ3oXt1W2hKcJ+Dg8KU52ZZott8nTDoO0Gv19XhA1RM3OJkMWLAqugUExF0rGw/EV6ONib4+Lz
tSwruMx/Ad9dvKZOiPxHN6o3r/YiFfcbDcPsFQFZJ1+9TXZao9Up6tEsPtCeHo7jOIKblgk0f5/m
zxo2rgOoNHei1lD2qQ9TrWi55ZKpMsMgaNy0DTFN0myPac6hoLUh785DB+fhi3E+eTl3lhfuTZdo
7ZaYialiU5rgoJiO8QejymIjMNw9G46m4v+OTlY/2RnxPCZntl74ubNRAcjHmxNlmKZH95BwLRKs
O04zmE4/J24X2O/Yz9Y+5VHhBf9+OW+Ngeuw96ASwwE8hFwRYx/g8Vyvd7YPAH2m9kHkE6zbZ/Bv
4/1ZwWZnnj26kXBmCxqN2+4VfKs05bfiSLeviO2NKE6HF2d5Oxa+QgLu+JomjMEt39q8NY5J+evF
hzY4ZfqXRiXzGxdaL+RtjWY67V1mIxl1+U0Zs0RPySXEKHTEsTWTY57SkUdEFUPJwCQ46vIhmjRQ
Opu3OLbFMc41Oe8gBodfrz9AYYT8Q2lHY1+xgL001O+1EK41kzlOl13jPj144imt8P3TRv4POOpN
5slLmcF/hYLn8locx420SwcGwhGgQtTSjrBvuk8RFPkEic3ZVFPJCoDgG2omjXuD6zgmK7tsmpHS
Lt/JoWvuc6fzHj2NHxdYHNsEqF7vg5zx7kHJowaeuJRHn2ETr90ISLz4ihKfOL/Ve8UBm9RU8vh4
ypLcmTnfpAIyiNWFQu5rI9ApFLJiBBs4pH7e7NDly1XXrCyqYwrgAV2QQZmvo8LBwtTN0XzDeGLx
ZzZIfvxikrXUH9OZDZaEUKMP5AfPfNyJk8bzsOhk2yECgsx5Vy/bNfizPeSMz+eLgj3h4V1H/dyx
8mmIujmD1+wf0+mAoniQfL1NgDvC8ASPis0AEvBgT/oCLrtCTgTnjKlsBZPt1qbz6pjThciHuKou
Y9hqjz9dz6Ny1unFgLEv2isutTR2jPs2bJeB/Fw0iwsDqbAhDIG35gvt9hc5MSOujqMpAMnev5dp
4Od3WwWXJwqxGBDLMYEVJE+N1RgsiA1RNGi40H2sYIu6XcHrZycKIv4v6KwuG/nf9NMPAtsSa1+0
iE+QhCI4rxTi2EpRyDWkGJxPJMKWIzhdwL8ugYC2+tEv8VsoJJiHBPoGEcwVPVIltFWKkcHP/XDL
mOarogqX98MMda2xDll7a4KO5i+Q/w8vLfi/c3akiZhG2SKjimzeiY7uBw2ffXOhYFLEpJFvQVcA
5o1WITDFnM0Txj/uo/yXQbwMDFw79XWVPkfxxED5G+B3HIN6obenOFlNTKlSc9Im080R5PXzfFvi
TKssBKdUhjRZMaR+FNJc1hXFvk4qwYHPMlbzADbvhJp5w0EztkFv0ra/602lzNYIZitlX9zdFxqF
tNekz4A1aH7tsPHuCyDB4XavIugAuRPMb7XoukVHN5BHmRuZzvWKEPNvs4t2NRIOvt4CYcS3PR7D
S3oomPe1AEAq7YltRwg8yrOu+3yDIw1Ra75tNp+hunDej1KjaIgN2gtKHFQ3LIMklXPuL3ui0KDM
+7/AbhhFxgcs7dBS3XnX15m5P5MINS0JUS9sC/+iwnyGqWVkZcxgYpaiMAullaooVbbOXUN8FTuA
/mfau8bkGPej9sjrTFTQveNOS8Mc+jglH43DYoIuP/h+DurXqMZ7H4MkahMYbFyOQ8tdYfztCZ8N
jXyeM7LDISMFnwZnYGEAfe7hdLenpuY+tWe/HkBKq4XkmmqbOhjMXW9gLpi544Gwds2vrLSJQMTx
agpfSAovkRWs+6Uh5hkchjMnWKRhNfZwLmfH6dIDdRf+3goZhhT07titIgamJ+4qDQGIGeW5aqxU
HorAhu8+YfETdqhBLM/Rgx6hzaaftR3QWso3DrvzbTcbAz+mMgCGGQEjkAiSFSnO+hqdqt9kvOWA
8kM9NJ8oJ0lh/3/2aOmLq5GafFZCJMIWVuAGbloC9KgzZ0oToA5/XFYLCLymwaSZbyF/BNh0sRbv
THcafCP9fxrJq5zt47n+sDy4ghm7OQmlTvikxfAOvYYfLKr/qm9eYDCbqGUzD7VQG8m5ttB2ejEF
6VtIne3mcIk/begxYdlm5Mv+2FiqFaDars4i13ogpiVLf9XiGVHz7VqU+ZSphz/jBiy4Eg952K0x
DLCnUC182avOtm4MxncKLEOTBZiSpA9jD3T+WlX6dRaovog+gN20UNkKakpvOw0qyZH/05WC6ISg
7UfwDg8vKxkyEWnn5fZE7GvTatLC1XtU62Lv71n65L97dCdrTM1i47pes7KjGw3Tk7S1/uFPzvTY
UZ5Gt4pRtOJoB9mEecEclpTmFojp+hJbrf1ZDQS2z3DwqQnsg8Ioqvx/GhpvWEzgFC1D/07TK3e6
6TSgoZkb7EF1zUftaUkmlwliK3qNnYSQVNxJiVWK1HTZoBpHe9XIVbLuCF7IQIn+d/j86BhJIyPz
8sDWqTwCpvEhocw/t2SJv9k/lJSFdXu13hMSqq2r/GLTfdojJmopWPDesXmRr+fiI31MbURfALAi
vI+QNAX34ZBJSm6QYkD0wfqO/X9MK2xuf6FVBuGwSC6HqkZSHJubWNpLA1LXvYVCONMhRdlR9F/u
bP4OnqIx9YYB3IQag3z+TvzlDkKxt36KmwFJnZSB3ndG/TlK4/6vj84jrzSCDqKj1CS+0w3e8uHX
yKGnbxwCNj/5gpQZtdCD3kvDaOcO5eHzj3lauDgoucex9EWK7XQEmOWV/+h6FqMZTIBv4RofWOLb
Cn0Rj0+OzQsdShFco0v1ltEdBqI6sTwyzWIUI3aRtYrTUcdEbgE1iea6ZCyCzYn8z2BXZUHUMGqN
UICTjXfuU4dcJwBKHRsbUm5WUNzW31wvj6Jiq47LBh/AJ4xh9fPRXARZYoieHzlYfHkDzMgtl77n
SknAZ9mDKQUmMKglFfwaGc5LI+L8VmmOwMzTHQXsqkiq9PhUNg/ehuk7XCklkUXMlhgDLY6171Fp
nXI71gIVQMp3eMwHaZWfD4AMKZkIHBppdp++mCS3DZMZma6u2In4ho5fVIql7HSHqj79ULwedF17
+bznRJT4kI7LFxJgiHvlJGcOLaaz4oEf3GlHma+aS3QiucFAraNLy0snH/U5sbezYrs+onFceXmY
bQuZUARSNmn5CrRNp4exW60oLF9cMT14uHqh8eyh2/++mBnPoVsHjSrBpv3jyfmvsZGIB0IVqW2T
sPFfhSrYNUA5rBrgBQUKxDBfUXcL8y4+H9uzwnbvmBCIZTU4NImPEs+2JRfOy2Xuy7I6Arls1fsf
yyNSuwjZm2PbLu1rclbKrcJs/Yy5M2xQHmyFVL9jejSDHrLtYJ8HZk6gRru1ieQZgkY3K0HzzrkC
9k0Etwh5tZ2CDATNDsgu1bgbI4NyE/12tYaLsSLOx7HFhC76PV5G0X/NAs54sLMF4mC5XKX09in3
+rO0iebDbeN5MMlprDR8KUAfR4ch73WgXCsZrIu0pbxPpjkE7SKrpq2wYWzjgBkjHktMbCd1zF2Z
pzE/YwT9wxJmOe/U67mmMPsYRTSC06X+5nuEP/Qk4cYi5XMCAc2MOCDfrgXP/eWG8yUGarRGYxBc
BbjntH+BvjGf99hjVRUOtIX6ofs6ahbcI6WG6H0ZrMQt6aZcoPdxiLPzmCOcSW2qFkDlmLIAsf8m
KqwKIZK/N96ZfiVfQweCZJz2+RHq2SVblRY7w9V2cFM0PVVCoQdoUxz6nGUjJR1OIWES2+w75vZI
VwfEWJy93YcsnvQuXQhL+c+/sJfXQufst5Rqe292dwvlRLAbrf2hIw0oNAtZv2eXxB2iXA/wMb2g
5jwvdbUpW2tLfJC2ZZegievc2I8rlKiRf5WYUVkjJMwtnk16SmkHhI0z7rsUAwqNdBLsKwYULW9E
I1Xz/UssIvXir8cWpDwrplExMjeS9uos72lcIgg9ZOlqkQN9fKpcEZD1DFNJkOGUS2O7psv5bMLM
Yzy9cV1Yr/v9RCf785JIQMi35oOPb3+p/ch0cEN604a0YsLRsx8D5uizzXFMZas9F/SWJ6eVpAVG
CgY+1hIi7MEqHluMlzlr3NOnEe2osXuBPEMArLICp9PMiFYSNnJGIBEXp/srOItWFiWd8VKRKDB3
pdjkoZWhY4mxCUeyYdjVAgnwNr0gm8Xk64XFnhjZnVFxTgi2Xwwk2jvDGV3r8VKt/x5eVO671DS3
c41M9vlRfHSqyGmul4vz1tnpn0JOq6IEzpFn+psRCXdq6zBWeqwo1wUs8ss+Wkr4iXI2uGDT4yF7
vYcWY8tGNiRY1jLfjVDIUiOn9VsbYABttsCOAVTHfFMvoBDWt1WpfI8N5UsPJxT7cEMoQaX9HLvk
az9Z9GJ6wsb0UDwvT6THUT2nsu+W2kt/KyaUruztuVF9I4k56z3LweXZKrqFLrrmCaxILZuFgPy4
xzYb1EhDs6BzbzyOs067vFRh+bdvO66ZdqpLGjpQ0XY4M4HcZkuDqjNlfBM8XCzqqaFd0IHygGoC
3lh81RJZ1idHFVaQ8ZcIaLVqXDAb9JhpyOTnYRUlk1lWaNN7/6jl5itVqtcKqj0bQMbHwy9aN0nf
vJxIC3MqFGVzdTrwYZfdPxsXQjm2WWlthXtAEZwdsTpcHdJIKcHD2cISOqFWzXUChhhdwMHXnBU4
noinLDxp9Iah++jW9O80BUHLUn3iSCS4VlTgjhbPZdOG0z+1IiOOiAKNCqsv1deKkPdQQ2Lawc8X
WdGAKag3yiXZOsKkFtWwhg+ENveUzBXmUHLPnAqDTlE683cA+7paVrl+D/+SjiP1Qm/RXLBCcv7/
D1mmOx5EmXtyeDpKTHk9fyiKpLhRalB910znBn5PARXO2PPPHfSL34LEFdsgCJ9j4+4RsmME0Hgu
F1uK1NNwTAn72pXOvDrcujrZcCsTahREoFgPV1H9giOecRDSebNsLpivbKUk3lWmBXDQOYdzeVDs
S2HvlIqktJNJBaHSWnIfdpWIvalcTQXakiwFm0I7ARHNPMHonH+8t7eUUn4dN0k/4IjHnzVFpvfh
ODskWXLQ01VsP6BW5Sb3eUSNdvZmIJxrrbKAprjI7rTThYQ6ro9B2YJElxuLKYjeyQKomYkpEcL8
VH9vKYSd9Pp2el3r2v3FTNqmljVIMLVxD7CHTcCcy3r0HV2UQuZRrdDe8Mi66s0uW0RV4IJAM2dc
7gwbEKO4FGGeU3Uklg5uK2A1FJUa8RFQs4/c+tWVoqWtAdZzgw6nOBlrhpbLfUGDwZvwTlFOqodF
rPynVYq51zEfJoDTc1tFSEr3bSJhnKxuZx0WcIoIWY+UvORq+1QPPEd4epag6xq4G39QJMdTKmOg
M+vY9GpIGjVvKz8Wuttjk3ehls/tQkLzKcKtEbKv4hDOOxdLDkLk7CoWlzrt7sCpja0pYXmE6XW7
G6+3S5mwZ5FWByUapG57e5bvcSwPlEevpLDh2b2o0Scd9zT/eR9+Oq4QCAlOGVF2BeS2mhGAH2zh
n3Yy7ir5JWh2SNVSXCvTJ+X8lGK0SshCStlanu36jqPn5S1BPC4CMLpry1VRurP4uZtqgIbKBrmF
UpJq4zs5/GN6Pw5kqh5d4wZpvgYPqpQt32zgqCgzbLciRYk2psyH4xXMdVUAIb1zaQJE5kT6lg0V
1M72yrfFBqirZB/ZCF8Zi2XQbegCVAM33ATrdk6ECo+jhU3JGGg6uV7yp3ovBtRgGIN/lFuR12GG
BRgzdqFC9WGjwl/Ns15cOxC8J7MlW/1//NlXTXs6jafRLVvirUM8h8GYnpwtlJWIDZtgejUXnWPM
OmEfBqZKqlEQCMcz+vJE++w8pcGZp9Af5X2xmyS0HkZArHtbvmNYgLhm6YvLNiLIpmW5kSY3CHN2
tdWYAe4PwApFNQ+fAUMvwOF6/jLZT8Q4QazIzRaF4+m1V1QIWDv4vGgSj0EwK/O+DIKP3yBgssX7
HaNCZ+/SBEZAQ/LYK17RYMi777CM+gd46rsYUjEASBzjuAg6WdWexh5nE5k/abLSWZZw8Bm8Lvsq
sQccSB18wbJcEtrrJbw55n9qu5TLsJ1zqWb8EpLx0T5V49NHJXZ7dlhYLi356qsfb0lkqTT6lH/5
7sVqjLpg9/OMUhrxMDOlVMEDZxz9n/B/yTjfQj252pbFuT1uAJSQFCzaZHhuttkqg5/vZz3LuAVN
UVyVXADhXJ8lhjqAbMiA9kWv1dYHlvtO7jPuhue4hpzlygko1Yok4PuzoGAT5BCVgMrKf67LZdKh
lKQTxL/BgqWFCkcgDJB8rhUSK0/Ud6j30i/LucEHYCvSmTX+aCbMEdpwJrVs2/AiwO3iRYSKEZ5i
p3Ht6ME9M9lWqnLL5UF4u4D1S+V9COYDG38MckdMgpi3GBcgrslNeK1hUlIu+Vls3NAYX01RxIlS
i1hwYKAQhbM2SaifT8zvE8xzpmgCuwdZf/725cl8k1qmBSOJoKLRvoYbF/0++8lCce6bdym70Phh
4B8CDsgffZqVnb6lVYos0QKq4pd/cDTiQPxQEakJ+XAhXoSyDxoo3pIt+i5Ztv9KHJmYY9Fl69ji
y6pLKx/VJ2eHZUw/q2/dmI1jkSydJvWAuM/+uFFiBYhHEIdLl7TrI9cgn2h0YPntNQTiu+IdQ4Hn
xFnzemcYdaVykYD5a5OVlhQ9rrIUkg+YDW2zHolQwwiBK6uSRPF8W4OMwVjx1t+iKjI0GMmu/03E
Rjn1KVp9a2piu+491M9NyPUI0ATpgLlFeuS3TikxVm8/2tLptFqfGvnZPbVmWxHx8jhYKYg3oT6U
7VPfNAAX84bbpgREUChFzOpe5EcbG+YupwI21N38mvkyxjQt4Z4Nnw/CDvVsSaWRWjnDIBv56elv
nFJk2h39IKASE3augYAuOx68slrXOWIg1siOSXqOiW+SVdIJG3ROvW08dPgfKv92SLjr2rF+pPBQ
Tix9aLxxGE66wI9220XHlZw0tEtad8MLrMG30H5nV9PyRwLq/y9p2B7WvepnOaFDsTlbmjZWovB+
dkBQVIClRrqQC7Yd1I1sg1i+sDe2O2bBOVh7lRACFV4Yg7nxv7MXMeWQeRB6AqE/LOJQQdXpHT0O
FSKMx3fTjOs446OaS0Yu+hb1WBkMQsB4oVwaTPJo1KWukmLbwsiniNdwoVIfqBOalGnpWF4JWUpj
Fst6yalW9F7MpsYz4ig14bQhNH+5KVsSaqTZBzE/ml/4gfvucghHnI8RZ5b0m/hvUVeU9WYearcS
25KnybYmlFjTxUOHiVa7Wd63lF3islhVrRM5oqyYUZeq/RdYZL9pNpAH2pgmXch6inzKgDWar6NJ
u82uYyYIUnkcyhNKD0aP06+Ff0JhGGbjSWiCulWI0vh4S+7rXdiK5BmjLX5uoYP349MkVy7fy0NX
Bj74H2SbiY4eWQdHxQrfFzms592ZNHISNnJ69dFQj/ddgfd28b48836N7A3J6DMxazdUUz/XwP/N
XXAkgtJHsbqlZNgIiYt9U9bO8CSj/igl+lS8kCAq4Sm5GKaFPOxfW3aLFVB7ZEMeFiM7lo2205w/
24OnkeM9sgPW3M1pF/Y9uSQNgYRHMU0OlhAR1NkD3xqVGQdixhfFXA1wSDtE1cWn/C0hKohcDvyN
XH1ro+X3AHCuLmFJyO1j5x4vz3X8uyQS8pSS05jtV7WraSFHqW0GvSVQeuPI4TvoFKUStEib0PCS
b7OQmsNZp1Pjf6ekfe8wJvr3Pb2SY94xziIX1LVgSLdaURm+5xN75dg0S8HFdO/XiMu7SDHUhJKL
lJKVpb0wsGslBP2GVmi8DTcb64zpmIsaboI8mqssY+jp45gSr2wnuDOep9riSb3PD/J9ssDwI+BS
Ah7TdDr+nuAr/Cqox8ZwKQUAQ3exBRTxqShtahLZ0waf96h8ho4prFyFejSdS+gAwL5VLmijRVBe
4SIJuDen19e2t6C4mkVr+p/Li2BspAkBPFB6V7JdTa5+qea8nahpMnpsRf3wjw8mQrgI8zIKaU/w
keZmJEWfKKTmuryb216QQmn2ESzTmrOPENEw0mdV3Y/uvXdGtXMxG41AYJTnb39015sC7uaJx59f
q4/hY+oJEQBXPqaBhWJKt2KZg4t/oyNFcdeVLwwWEEFvcuZE7ma6/q55f6T+3xnnQnExdKA9ffY7
w8X86lSqOqKk2QUw9r+JW9HmdyofWOtzWvkWYaxXXQKwtm6lZ0lN2F3FAtheqBE4rD0A4tUEDsc1
MiSjXPljC4IP1MA7D1Q7iDEhON2n54tnpQTTr7hiDONfvF5tgHSJNQW4O3uyMi4y9eCthn/qxFVP
WZN8JLPTH5fI4iOvDcMJ384foPx3d1KNntDCKwyj9pIrEyV+6Ez2YcJ6iDzYd5MGlch4zTBjDBOc
9GaLIZVH8mOFBjI1TUjU08lF89cVfTR6DR1F3VJiD/sjpIp8IXCgwqXj6EIIBGlpddF/y/afuwJl
w/oJCQD1RiXgoc+0UJG2smEA4UyM25au/i9V7giM7t1BeDaJjPb55z6JeNj4Od82WSpM00Fjv5ul
1HaJFdP0Kop8gbJtUFWtX8zMxWGr7ILgeO8BTnrUIuPxxiYc415nodyFawDV6fAQ6T3SVXaXcv2p
fz5bNCU2pKVX+w/XM/xot1OJzeSqqytIhvrNrcRH0KaZIcwAVSassHKNvFG03nSaPAM63ifJUXUH
GNsmeUguTS+0yn2e2DhM9+XaNUzyBfD5HDLZ9+mHjk1IXldGRX0VU82ADuE6M9mQJzthgKV5cZO2
/H3cqzk7AVJyNw0CLstiKDB9ZFRTByRDwdH7RhnUCW46dEmsEw6S+jztu7DP59KoDxo5qN46wJGN
QmlE652Xi2G11Keb6MeorydlDnQtWhabU/YL6xX1k5ucK7x+f+SFVuh+gf3LluTFTZ5mOQlonE+O
/3PEATgx2ZdXWtUNaU3OhYC9pAUn5ugvtdcHnUAyW4r9TGosRT9NdJla5AKnNd8NZJ8sfKonzEGm
TA6T3/Xube4wiTZH/rPI2cC8FWtjamLQgUhbanspxTrPQhzRzHU21pbFnFVfkXzykC/gB8FS2iKM
zAbpPxp4sjaFRGoyJsQvGkMVLQVC9asI0Zg4/hBxywK6JblldfKaOiMJyCs3gkxnG4e3VvVcRlu8
E72ns22rvaF9RkJGaJEm5xGLYbLoYHvVALouOm4QbHDeprcio/nAqV4Ubfe9WhaBPe+QGtG2/JhU
3hBO++1YKPnGd1nWJocjrGaRSevg9P+8f13alnQoAN0CSD3QGXr3j2xy5xvMajnVNS+n7VfmBnqe
Qlz0VLiEwfypgFFoYTCSDVmywDx8wqK3NDkruHhxUHzHSORvbTQRFAmLdyyYgSuB22F3KopY7nyI
griaAdmhvyxQW9jz5bOYkRDhhcI6VGsd3ZVZMT+epZc5iCiwBOlQxu89Df4zLAP1YoSFDX8yMIim
yKLlp7Q0/QwU9aDiep2VKuhfES7huQ7n0NfEfwf16UUuR1QhYtjPuvir0AdlC57OVbZ6DDk7guY0
8lrPmciG4WV4VYmCgLBW0RAyPkhmlIXnSiT/Ubf4CeqJ285PEIDmUYwj6L7dKBmXMY0qXzXeUSf7
gE/AjZwkpe7l/aYgsivh7xkEijT3gypDIogB9YHCmYUnKQaF8KTDw8xP10LhRYwYtPxxIvOoiAih
rgyAp5jAgHjHwNG9QStzbqqUHS7vvB3Cd2jPCL3N5N5ht28dojg75+88Tjv5MwqXA/JvExk1C1Wn
SjYw7JE0AzDs1+JwAnTveXA2QNwaDSi/v7Y58NWCMm81UEXPYfosKL/lPTkKBb/RAMYJanHNtHqn
xRv6sangeUjtY+MbVM70a5SOwFLg4sIaWPn9i0cF+TfU0N1Ie553+5iGm0gGSxn0H2O00sYdlzor
vHVBJukv4wn/NgDMEuN1INug8GZs7VqzO5QBiC7MawknSr/Yh/RRRMa01ntXSwMWL5xn4Gju+qPZ
KchIcPZvAP9O0r8xKVBrjOvO02SJr2t5Pi19/S6TxIgiQgMjAhiu5UvozDfjbG7rBXRhERJa0M4l
9mPnDodAYKC8kgk8Pjlk2Tdi0Gn3+9juf2axtviZ0ltM8U/WtTh6mvBYDBEaarjlQf/XVsxEAJ+/
JA2/UrnDNJlx7BihCxqkcJ6dX/0lwBtks0DpBENdsG1wF/2jN7K0k1/TQQTKFFjZ7v7J7OVYaYwK
sKFZOw9/L6a4Bv2rk8CeVY3Gbvq4qDDNBuyOhgetwAdg3IPjuzNuWojCq8O7NVyAkZCFUWjWAJMH
vfFOt4x64ug64fW38ceVIUWUZTUGd3DeAPOFLmhLH4QJJAFyQFHx4NvsIy65i6Bn8SZXzwGUjT27
VLzwDn1Ysr2rNDowkeYUGaKkG8gSEjIvDH4zm5GQ34gdtZzVebEnhMh/IlhvSw+qs7J3c0y1BhfI
AXbSJWk6rES+EN+5r+UcN+CmXEDM7kBIPjL/gOQrpg4W0fVtoGgZfaSCUKfeiZWTDlzA7bADMKGq
oFUMybxhtifQoepDRAXLTEJJOEetcmv55hlW4rypdixA/UcDyX54jvBBbY2yDAQyN1rdOl5kQddP
dCejF3Tcg/289zsHdWsX1Xgs4hePbgRbuajqAqpiX0PKf1aRAtxnhHjgpxo+yRhOVmkosa1zZCHc
uVDS/kTbn/mfX5NUlE74JHx/14Oc9Z3jguNFGE2tdFVhIQv1hitGCAdbnMEnwHJFfMQiSWPkYf+G
NJ013ousSpeuWAnm75K8oOsdPZLsmsHa/VBWSOGmNDk0A0GGkJ3i60GOX4J+VGa6B+/yId2qJixG
w8ToWWcQdTr4Kw/4sJv0KRAlfy+0NV7wG8LxThZwNf0bFAtdqbAVdGRO6GNxa3XzhfOiGAPVlVAz
KYYKJWBCKdv/hnbwCMduFjq+5JdM726KhfyHGeP4daZsxnzNX4D3+vGdrC1pmgKYOwXRw0CFlSG2
20f2iDfozGjJjKAycZ9pDAbpcBZ7vs/Kg1V33wFJgo33WH9o/4Ovn5o9aYHtKNCttC6azxlzQy/a
LFBcH2Um0aUy8CCfprREYxSd5FWKNoYAPDUQgQFKBFJAtzui4RMi32J0yw2UCpi9bMiHdOGyvcnO
cVYAzfOdxMbcbeASfTejzMHhhzyGR4LQrnIMax/CtGrX/e8AcAbrnAEoLXeZJfdHkUILuZPghg92
hEu0GQ3kIhMg5QG1PtLEAzSnrw/5LlXSQzALRjDQ6AIMxycSb1Mhg04Xlwqv/kbW9MCBbqVAa5f5
eu3dp6adLKgDVtFg/GinSogohXnDSy4vZahRHm33ZVicC9JHTIi6BhFZyK2ASLS8+EUH2GJYv1gU
HlMTPDebycsBf44GdQCEYo0wp+c0mMiZbOPZvFZE4PY76TGXteIw+7ff7BXKQEjQCE5A67Ni9Kw9
AEM01bHbMgvxv2jhZJeNMNtexsohO5Mtfw54dmKwjl1nvB/HNYAtUUDEAg5HXLh/iwROLR2TkIut
llgI5+CicX10IGgQ9HafRibgsULMYF0GZPk889IjSrYXzpL5KxFb+PB6IcpltYqmCMHhUJxHMRMH
bN3+sZ88YRkNM2cWoOnw55KaG6uzx9LmAwYrJTjRjttPQyvrU/i+uW9+91OSU+kagK1fo5AtJVoj
H3rbKs6urIfCRbYFz6snJ4gBSZ7yEi3mEd4/tzT7R5pfgPJF6ZI2WIDzwXEZEejoJDG5hJUrJsQj
mggF29RLN9z5hGzkJDX0o1lsmjD2duP8OU2Xb6BTwS34OJOKd4p4x2m/DWA6XaVJfuPTxNjeBU6E
iMP3R4IC21skQViC+2oyUvKFRMTY/J5FL6AOUm2Wi24OCfV3UshAnBC2mNzfphMgWJzX4jkBb4g3
kWUXFP8jlLoXBmEEpJ23/kj5Y63tRYKwN370IBskSxhH4LK2IsRXlDow8LE/sieVnPXQo++L+csH
HFus/xo1gx/I3li+G1UUdSq6wf9FtjdObtTuxli4h5SJceZWN3Rqz7OwmejcQpFb4ltV5hHp7wg2
wt/8eaBocJ7NBupNW+uU2GCD/PcVPaHi31svxi5+6B9qoHUl/lQEsMN6nZq7o2msgJrAYYyoTpy6
02K1W+w8LqITT8zuMOqGyovypgytKvysCbqqLJcYlxN1YYOhp/mdZzh12RU4W0UykucxQfjgsCuU
Kl6M+2aybxBYcp4J2zqFj+AyRFn+Vk57ekOIZHgx+RUKqKgB/GOQsFxoEFcxRNM3AAHpISCKmW3l
G7YfOCr48FEZNNTC+66r63D4FFy7N3BTiuAgLiW7gjnRAFDtUJKK3NgzANdGb9COH0ycjfgZat7d
OboQp5Zi87AxQrq6raqZBxOh6/BjsQyK/t1urRBIjCh2KJyZ47Mx7kkoI9hkqn718JfU3MDJkjjO
M5H+JPnXE+5m0LqAnGX+7wKNAMGqrWX4o1BZtu/z3dKVucUlxI+Do7Sr1JjiGpj2tbwI1tOygafY
opfk5dtDF3aCB0uNf+J3nLNUUo4ELiYNl/nxcMoaaYakrFSwGpjx3IjH8S4gpYZyZuUsd5AR0S73
ixuXptRUj1qP+lpee8nYNRDuYeBbYD5vugKcHdc5LXNtLduGPqIuoBEfBy5KBSr5FweXkF4pjXWW
jWUxB7WDeoPWvSgcLgNRV9Nb9aiyRuTEqgX9e7rsU3PucqkQjT+ypjrKFhnuEk+7kiWZYTdk20K8
/MD1L/Akgl5XuehBnOb8mnw40eqxkClTzLStAPUe8wU+Y882PdFnDLoMersOwjkldjb8cSt8O3uZ
x5ZlqBjzPCcdoD62U7n7CWJhHgCdVeBHrWorZTIle49FaMrQJPPtKcCAxxQb8MJR4w5XBEq9CfMw
iKVD2tEU0JnZxVcTUyqYT5tQKoTuFP5rp4igKjMAMP+P+LNFuaDJ9mpi2FB4Rr5di5Xe4cvRwPNR
spN6yP7wXg5PX9NfzK3ghJ1dmN+ElOnI9UkLUAl/V3/fy1wVgX/VVakCVL8WEG8EaXHVYyyH3pF1
8hJdw7N+J6FYgGlwdRZvbcvrjUFXuQaJTTRocPEoLFn9xMIIuT7Zxcn0Jtc8rTuLyWlz7pi4UNJU
TDGIDEcZkgfkdbpfPlQjjl/x7xDWQG4WYQRfqIL1bfx6HwXq5/0BiSxmp4CqhZLUHfDzC0JXX3KG
RC1Nrmt5koC4XULKToXNDzcqQj9ZKYrJBqAZiKNyPpjsmThS3HrKy907TPw2ZPmpp6jbTa9paJLz
KjbCpWniqxxg3YE4e6T3nHLAJxSW+v9ZUw2bKNL9tfwr6lRyMaWN0VwRqlb17sI5TwWHpiu0KIux
WP5Zhh0hAhRnoNn/CjxlOQAiWLoh4SF1GlNXiBJYndzSlxDE2+V9CX0mtn+94q+1YU/7TrfESyb3
3w8Fyfh/04Q6DSkTlbQCm2jRYEm5swObIXkudcrtHex1mw3V/k38pMbxKpuBNp7Z8QPTDDaLnrYv
RFDFx/DMDcIB5qPd0Vsd/D+y7pcBqdvMLzPsBllcSqNGccAxI6u7pVRdnrHtXSVMswVyRI3St5A5
PMkOCt/sYGz9XcQplMRU86SgYicPneZOgqfgaXAZCj0Uxf235Qo9Ha49cSsNvhzgTPtsHzA/aLwu
OYmvypORJfQqfGDtpppxAeu5POGNXnKpXzCL/Y2qFyAI+GTP3NkuSh0RIpxGHht6FTB77mFITPnu
iFDzAweafoPsmNbuTHOYAxU41smCEBGPmUZBw+Y0sjg7ooe6OJAMzTQnIdNIXawhgAzEp0CB97Sq
C2sQISbP4yhDnt+AjON6bagAte5CzzcCRpGhR091pMsx13qkRRykqhWTd+41CWR3qB9F2Pn+EpBA
180ejGO5ZFMYucZD6l4lQAc9IxK73OOaAIvORQ+MNxx/3mtQNzxkfeo6ulTsb9BN544scQTfL4bP
qgBCTdET9fi+RpDvLzJ+xfsSvqXnptZLWi6+JTC45TjRPwjh22XZ7+XXnjOQoQlBfUERwKWW3LvD
Xww0TQFnrgjBFJIKxi9brjkPwBW38gwNeyrLUAgSc4r3CULYtmv5Vzxz4ZCRuOk/6uN2H0IQ/efp
pKKurUZtC4vRv8RxpMsxCVR8XAbuJoE1CmSU5esslTxOwucTb/MkzhjK58QB5Fu0UKb5zDK1V7Rb
5w95htuGdeqt08+2tOxpB805bFNFD5l3c5P6UPUaAhlVzj/pT5gQ3c9awagHu3S3Vy4DsOjbm6jJ
P8C773LFZQsEhqdlntm2rO6qjfsdw+uVl2svA32e34wGldMLjJvJudEsr6FXw8qKAh8oCJgd+l03
KzTdlHWBWUSyyz6JXPrajf0y/hBYGqJLfI16EAT7h9GPsQYYZmW75KoQVNU4bpw6+L2AfhdhxS9a
ljKhchaPyRnjvRyEkrHqT2mXMdqj9lxIeTt2wwI43P2cbaQHGd0CN8x+2ykpek6rOoDVGcLUDQmm
MdpYUBVpF6n0yzqBJT3ODEyvN9smPb/pnY7zDiTVrdP5qJeMmHcXHUwVAAE+Qz7nBgSjLyWRL7+B
WCM1fDtk6q4FTv73zIiSfPFaVfDeZw8wHqoPyKLj0WOcZuvMin46tx5PzCeQ3eVF3PumjHo2HhyM
6eyhzsQBeY/2LBahYkedtl0ZhIrQdaSz0J57myM6eLWFE/6gtT5zHIoF+sFbQD0dWCjzBH5uuVXm
3a0JSYbTls4DRJWRbn3Wp+1R0+nxPzH3moUUg+nZZTX5UB0yDZ4a3NFtGzn6UxyyrY5xGX7aHMle
XY44UWRJyqFs/+kc9sQyKem1kziR7eL+u++3Bhz5lTf+QJMJ4A3e/yqINtJ/B9BB7QUYmebKJhoD
LpNCe3VWAXCgaYJi8wql5RQV3BAFYN43eOV5iIiIubH3DfFDGqvmUCXc3dZC2Ke3NE1pJnVMjNAz
uqNp34/cODCXTDKSMDxZgyptnvKUYqlzIqKMECpFsCf489FPgKQKJ90XgBFHSaD9vWp0Z76KDo7D
+BMBdk3QwtihiUoj9s1lcB+x+zleMLElzfIaydOG4D4E2FsH11QbJgUMI6exM62Yxd+qHy4uwlvb
M3n0wAjPv9dzmFea7XdDuC1frC0XzmGbZFm1efLZu+77hgP/SwdYZc6JxDVYf37cMnd++Vr+yzCN
KtsOjf9evxH7O+ZOOLoKdp6cG9l6IG3X4CiW85Bnq1MApDz2AOW4Q46mphs9CoOoQ3qg7HVHQeBH
g7U4Y6lqYGclRTsTjlZrbIUgd0shW+nGb3LKraDumhFND63EzS/1EdagwI1VWAA2Mwp2NAqK6fmv
R9rJMyGVm0XoBZbS3fRwHHMvgf+VMHLEl83B924FhyPZmiSIA6L6MqekuMRnthFzidl1We6cV6u8
n3QSwfbnC7A6ePkQC/6TNRIZY+rj4yMFT62Dhoon28lOMUMHqNjEMfj7pa9LshkGQk/dApQTBeLg
+0mLvQRgoC0Qvam+a2E2+itBSXznKq6b7n65uOKIJuWeIlcdjLR11wLpqY/SnWWTZO527ioyI/nh
IHpKjFGOaXQ/PuBAizMN+B0vIwniR9pl7kVx/cfn2+Z+9qe3ZK0sxUc9ZOz8UY7vxnrmcLy4WnyT
dSWvP2Am0OZ8n4me13J/Iw90xshCYsPK/AfdGOlGQO0cQqH/b8GxA2IPoZshDPM8xRqz2BLeI6IY
l/vjFHC97xFVQUUWmJ4fwYbeEJ6kEoXn89HVHud7adaX5y+4ha36SdqfXFeSYy173YbPyIqHgnIE
z3OzqUDyQPccrNCYnQJPk3Hx9KjGkife/5/McPaa8jVcC1BbmoIvRxUSHLnhnUKBS8N+QKqfjQVP
VDen574l20k1QgJw5Vs/4Lf40mzW47qbO6h7bB5gHYYqiaHT4oN3ADCe5Cak01IhcyN4C3FHxhyn
DB/ThUH3WAwomSEyTuAvBCClYAWvsSjDIPE2WCs+ln4s4w2+9CQPt3FANb1DbSfbqb05jBdn7HOa
UWQfebWMcKPsAVBbrIgq1xMiEna9nkb1/+dRkcQ4ioenYojJhSjt/7kTDfLyvJGMihT+Jdo4VG/F
NYu38qVtiRCRQGX829zVe2KFeIT9b2TdnzVjYVPbGsIIN9Nwe5weAu1axghnDKPJvC7M0lnSqs+C
f0CUme13b8tYtNRceaAB45nt2Mk1t89IdTCgHgUWlQrStK+IzFbIHqGP8jUdYYgtkjRZ0nJhL4z3
i6HWV43X88ZROBu0fL4JNLWTvRFf9hyHb73KFjdfqRF33mcpA1ZGmA4CZpObGoBgMnW1L8y3xrvA
+LGO+HK6HYDL7DGIqvadmJnhnsKDkvBmGD0IlNgyT1JjyBgE4jRaWElmqF8RFIct38ozPaUkxqeC
2C5X2qnjFQozDl3xsLYygJzXzMjzr9YuwWOY2pBhSH75h4UaoL80K5nc17o3aAar6xq4cmrabpEK
b1eQKicnXZY964nYe0nWsTJG6yR2vT0TG/YW5f+Luw+T6mxp9gQ0A1x8h9LIMdjU73xNM4bhfzzq
021aELQB09PeYrHILgvsqM1z380MLtEx8VRo2671qun8PLh0rJ+A9TFPzRkIB3i1geMZr3A2O+FC
F1LhXSAKgmEqL7+0Py0eWxEdFI0UwaOjJwZg1uJBU9QerNTBld3uz8HiU+WWvnpyayfKAIL+cq+o
/C3x1wBqTFCRlB7Pb+BKaX002fJDDb2PloF4OBMveLRSBxjxp0n8zp3v9MpQo0IIsvNzpHymfYRo
jRaJQGt6zfDrRRJRNvdkBei5Rq3Ezsv9ECNT4bWWleu2PpIWElc5n9gW0vKln9BFZBDbbDS34irh
irOYXN9yU+RJoXaECaezjDhw5xOPYd8fMgvQi2A9uArN8Sda7JbSZardEGt5eOvooTTmByfLlCzB
x/kNUOkfwa2Fo8oCmKfdWgn4AGsGkzBLYZYWwTIy0E2dpRlwat1Y0HDvwBjGAyf3UOtxdJA2WaWL
aU3bQOjTCSubZovBrScDxhqQTLwV3Mzvv5u7VAOZXrdbfezeJuadEriT/v5DPKDrUyf+Itdf21Uj
qZ+MVpv5RxbAvJWmJ2fHLb5iZ5BKfZxNcSAoIBnfpnibVa9IHaW5DgdWCEuthgh7C5r40OYhgjb8
4wqtGzsIejcWrHiLmdIU5bSPuE3kYurrdwDwfhyRIP96kup9shlyFPZyvGASzyO5CEoUdYFBI5wa
V70x1INvOATkBaIA/4OSoxhN76GZH3E6szXLoql4OYN26wS8cAIzpfvF7r7ve4HxGdgX87ApXWkQ
2uEIPXaiXP3CrXahV/CqA/RySjQHprrYTHz249+xYy8CCql5JihGsOJwF4vV511FFfuxIlRgMK7U
MEtDUWk5A9HJQOK7zERBIaVejM7EouJJ8qh5iSk9R2Gm0GLhLgYSnSbh1DgWVycVJ02RKqHQlKlY
0qyoZqaBgR3xbNjiaTvevzzdyCpPvsKnkOCu5HQpdz500dIsFaIYJMPzvnc9hWB7R+NWkHxMKw2+
IO0Aj37sTBCnEW4graw78qiM0RRQ4WqsPiekNSlLuvcq8y9rYZVSlnqeNd6GnH5fDerRKvI3QS8J
ZE9FGxGv5r6Jln7oEPsTEWclWUcll5GSVGg+cNZK22gA4FHkzVR6HX7QefaKADgYsJjHo99EwM4t
tc8xycgtalNMifptblXzFWtRLd/y1vZqeYrLq7pu4qHgGsJ/df1ijEKUQ/Cm0Z9xV/Q7RbN3RDh3
Jz9iPj6JcWdF+tpQRD8uYqvuOitXob52Z6lXPLQBV84PcMWyvFccP6eZZcTVvwpxUwt+OgHiPFXo
kwO6CX5AJrGia4zMXyGE8v6YGOP1qAGhJDFBn5RRq6kZyQEBRewz/nnKTK989CwJCwNrTBUUYJtH
jKwACZ3Tycc0GwYmaymSP4hP08+Ze146yZKPDPuhNF8hoP+AMVCxa5pImR3oZy+y2LjjplibPCKR
TfUvWiLhY5SGJzTtIB0qhqJ1Q79W7kbhZk8XJNEJMGc3TfO8spQJ+CBCr3RA12ofXEJ4sbBdk74f
JK5T/8h7I82n7mQ++6YrB1cShl4LKGuvVA9gbXapS2cti/I8QofwC3hhKodCXEZzjbgMM1T2b2By
X1izrlWDIgw9gBYHp1xLrlmlE+ZjEhR+PSK5gdsvqHz6L6ElelJC1Ogkmc4+proZ8N+pFy5qbY1N
BS718YpXe96sw2zfvb5qIHxpv7r7S2f3sOePlUkIqTp9o/IycytGGUReQuMdFMwpteYhz8ODFmIW
LD1odA6nx7c8ll1tjR7dcvos5DdQxl5i8wEafYvQ5m+ND/1jRtat2znT/3If6C/BlNqKwCLX5iwx
ghkSw8dLGFPYSnx9HfyxH3jLSSa/LCElpNbojNCbeG9DrfalUDpionP+tEqLsUZ6esrK1MHjbUqd
6n0H5pXc/PxnUiZAdQY1MDFTPU45qsZ92UIFMQsdV444Y+sDp5LNdRCN/+bVPuRL+3+WzQKoP4NV
C3GJ17wFdFma2f3uRx9DJaan7lVbu0nbWfD9HK/aUAGBPqP4n6EIJCtQqetv1GiUvZm82WQ5NB3n
lqO3cta17HmmYNdSEnDwbkk2k9g9cJR8DHqHIEueJTActI1ofgGexb2fWNhOn0p48+63gcSDGXfS
3PgkcXc6xs+QR9QBkn4RFkxTm90N+G9YQ6dY1mje5e35QcfX9RGAkrf351XauFSVoBmt4eoDr4HB
UOUpSuleWJ9dcEtImU+LuIuY6mJ7sbhYpUuu2QR01pTbXjgH+qf+C02IOSOTSmfA2ryH0YvO7FTT
LZ6X4HoRxOEXCnBe99vzVWy2+noKT7vmDFGvDiVdWxYFOgeZOCdPiOCdFeOr2zDuNgft6hLUA4jU
eoqSFIp1Cbv8HjKJXylZLPIhz0JR86NSB4k39s99y+Du8C9C6S2Lhpt1KZedmTGUL3A5Sypbnjve
eMcaY+M4v+NXHGJDC5k/LVaSYO9KmbQw7D3NB4qJzI52YpKqMNyaYtQiLf1wIy9xmnmTI+waNew3
8J+fA+D1aClwaXkRdFX8S3lQPCabBoKLSEfW3iu1nxNa2jg4x/Wuy+me0YnTiWEK+5DL0+sOQGo9
/Y9eDfHYCpJOcJn5x+q3xRfHEFiI2uam4604Pq877qp9I7W33XSPrMj6ZzJwWrrKWKk2z9Bz6Ayu
1PAlp1+QKR60RJuZWHuEgxljUEATEFXPZHvbBa4z2jzHkgU7Zc3CRIKdZgQ7CKXYp3h90jz/BnWD
4sjX+zg9HbKC4jv/uBOIYT830F6s42HkdSYQ7PhN+m+UeGz5Zycd/Fh6rdu97mpXSt3rBCPmPbY0
Ykkm54YozQ4dA7z9mR5udT8WQUnCFxZ/ds3GVfgYUNK3XB650VcYhenfB2YzwPz0mHxRBh9CtidR
S+EN7luGQwZ8fYtWsSHXXiQiGLVNmdWpwQ+AjdhmPsSpyVewelCI+AIgNoDZmhBpj52Xoahvpubg
LlXTdHDtc+maoT8pbnrrrDnzcr1GhLEq1cSBQWMKny5HOlx2+napiY8Y1EgtoDtB3ePhb1bhl+IM
fBlN37bul9JAjAcEP3s+/tS6G0z469x+Mc3psmbr3oOSCuh1amMYViQkmwGN+R+SN+UWmSrkNWQc
AN79ESUoCHnxP6x2QFqVhTQ1rCsSa9hQkCLALcY/I9KbNVvRPj4CKRFQ3P+zByA/CAyL6Zp8s8c4
DtdSEXZTtHEQneeRruXw6ZIltscZrCmvxtqzJoJaC24tlmbVWBknyu3bv9sOx9tk5TX1VNDPJAhq
3RjkfbiJXSgT6vJE8cntVYw1YOv0Idg4bloikp7P00+6aRQT17K3wCm2FMED/D7/5cDBRSIsTCUI
1wFbSXY4yTvWewae08hSRuLaaGRwgybe9xbIhyQ9QVLnJLlGHUrKBV2cKuamU8grhmTw+i1uQMk6
qSzRWi8ZD1cdklmqMq/68tCOzxFc861uyun1WI4kgAYbrnOEglwwXubwRjMO1XP6wrXR6Ete4FiY
PQPeCS5VJW2RylZz7mpv2rAit4NuSda3AXgsUCPI91P9fTuCWHsxpdxiB1Hb9i4WTg3mJXr2sQic
kQt3G5SwSFLOPCr5xSlI9XIDMSZjuAH02VWzGY1uD4eJuhpe0wSs5MHwpTnw1u9e6Pow6y05FPW9
+J6HqzoJqR/PyVqG9bV6bL5ol3CizFxcjJkp/3Nqznw0jpAIdss0jgbf+3hCBfBYeoHzCcrWdOXV
Lnk/PUynQWBsEGvkx9tgaUdOkMSoDrcCyiE2uhM9aZdF7pi/jekk33Xw3fpn4ul1sWx0uxdA4LUa
Noa0r4+SYavHGeNbjugGCw0DKsOxfBY1NLwRvjjO/j6VuqPeyvi1FLz9bQjsaCOYbkGYEFw75tLK
Oyne3GqNpKhqqM68pXyi8LHKZkQo5hxXeFL2FEuodPVSjTUe6N8rCKDN5dFrGOKH5iyycE5I72Ke
dbpa7aM/DOh4T98/0G6Kfee0DH268b9ACcBEa9G1xB4kklFCe0Ij0vqJmBG/ekUSm1Hvib4kJhnW
E+RqmuvW0sh41/YbnpUuRtJO33XaIP+FwMTBBKDeBLN7/i+FH9/Xn/LcscqGp/Gxe1rs+yszvnxm
RyI6rPUchoyALQOwPHoHocL6ujAmEDXVpRnvpNawfpvRK2fYbojGg12eeuO8h17ZPZ4G2tg2zdjA
BNrOjgzcXqP9q5yJfVK4URhZjUo6xjhn+a1Hwd9TVrhq0jJ4LytqGVjCMIZ9EQJOIYaGH7H7DBvm
MBkLSVlZMQPK+J/OZh2MU7n2nSRtNyeOwD9BW4oFiN/KW613uwu4TuCUQRkJVbLwb0zV9YIbXU65
xjceRcuAi99hJem67uxcjokhkMLM7UHmpPtJN7gG+IuSenkk7kUTqHnJjylJttK6ivq5P4K4GA8U
6o1GWJYvE7K4dhmzoRXR36hDx96gtSgjttGq+yPMFcdJyNiep9Mk6G2HtCvwpFuPPWFDWTVZSCrG
eHovhy5GW/N2pEfXHyNqVyri5m+kAuC3qCHd4E29psIE7N7/ZBKlH/04CiuR8hSu8bDrP1AYjq92
cy5p8Trep9z3ELNDrJtbU4NO+H36kXQhQdYAer+aN4bYeZoRRwBZ5sQGOsGKEVQsd4bqlR8sKJoP
2fqCoAwsaZnlZl+O13QSpY9fbny2yJ9wITQcQTDcwMyJ0rG/4uV1RM9skiOT4YzKnY2N/pBQm5xi
DVNjr5Hg3tULrvRMnR1l5dp5+YvKO3yJrbc1KrshNVVvGyO/gCYT9uN6gaUU6LJ0r2nL65fgxvpg
vygxpvEAAJcX5pXsCeWYpexgm7HCDgaRC4insu+Nnj6CWGcfRf7Sg1PaZFY9LwmB5rXAOcvXKyuA
cbfPCjoL1ntTBXENCTCrn6ptiPGoey+utnWdoMnMkl9FbEm13LFz4qZzjmnCON2Xm4z+BR/OgmYO
VAU/hMkEqVq3V0vs3uPA+OeTM8zU202+Nqke7wAY0j/MmRWDFkhLNahSI6JDQON5LDZNB429xLRq
5MXUmJSyDMhiefHOrhZTL+5qml26IIGiQVNxrdWlmwx4fAEnpK8CeDg+SmYfNffLnatibtCEUsCN
YV0pD4Uo6gKzmB60Bccb9UhRUYZlFdlDufdNeubz2Ez2ycBrsqN9fuGpfuQXjmUAGav7l36dVrOP
9XBWRr3/jEh5c5sUCCAggzivpRBpBcHVsc8tl1Vn6TubXaAZfSS9SmGLdineciHkQIPgX2s7zL0T
EsAajcoIjsgppkfWgsaV+Bj61JkSqLvHr/0QOiAcvCnnzODEaEuO9J5vOOlVpqKOFBOhVKW9ADSk
JLbjoV2hhJWjTP8HylOZ/WBuzjl5fZDC4XgR2GoREp9dWbcnky8vOq1PaKYkHRmzpxOpt8Q7Zsyn
5XnCFTZ/Q6BcyKWaw3JExQoOQnbIDF5alGVMm9dnl1e9Bt4f6dgso9rc7sq2XUnVMBUK7jEjhvMR
OMkEp1GK0AdKhqVzxQcPh4/wUpO2458FDk94JZj2+V2rgLLuGiyh1T5kT88kaBUFTEwU7msTJ66X
QicZuOqDSKJH71BYYVtBFVzI5Sl5m6ZLBXY+dJQxMSZR3LyX0nH4eq5ypU8QtGUCnY5L5/wgXzGb
MelEGK2MgxwZokXPwoXPGX+m+vd9JyV9ah79PP5Ztd5OKyePuxnwCP1KjbutaUHBDxpifA1TaG4x
AkPeIPcYzmT3mZaM/iR59trdpTAEtYc6Ue61WfB7RLumqHBkSw53340i4VSH4DUtU+Pm0xoZ0YRI
SSNuZDGJRnWPbts6+e8OwT9TqSGtIM7qYHqfI4lDMPeajmiQZMjOhtfU6fCflrWqjrP5Ah7Eb5dn
opcM2IXUk7k1eet4DBsZkZErpyFtlQ2k5kXaSpek98tpAQLma4TmEBnylQE5U+dXlO4Dij2K4gtd
O6UGpurRJenvkf1NBlaDbv4quBD5Dhx29LZLDnSMxKuR4vZ+ZsRvVde0DwlmqviSeSPwI/w/qnvr
epcDlYMPhUJVchSBF7eEFvIKzafmgSHAST3aMC6TCi5qapAobbwi2Q0K1pXW4kB9OfJ+BY1OfAll
+Anh6+kCNm8PWnRKcQ2B8+Rosq+im5vLG6DGW0WezMbgsfQ3t1WpIoIGNZ642CBtVhc6cSd8YplA
3Y41TDbt6KMY7ct5nmYndHwCqi3jiCJqmrIEN2i8XXtqbbxbn9cZDGRqqgcl18kAn71GIw2t/jEZ
os6xFW1YTRS2c/ZXlI/WABkeTbt79ziBj730ho8Z836Idz7lMk0Q2hisb8Kw6FGcrjrA22A0VfJG
Wge2QXRNko2R11Zh/3vXjKf5HP7I+nSkVpkB0j7X9tojCF5+9OrcIdkYrsO2qKaaBiBa9Oebpwek
F6oWFeJ1JGRE9uQiqOfFIEvnRXnuPYo1JMSA8scIMhOohaySYZ4BnKu19m2DHH2M3zYQ/MBgkltL
ZWi/gp1qMPLtFa5pyXDktIEPP37vsoPH1IQiIbD2e3JbVESjp3oh3o6Sn6tHCIR12AMjWnBNer9k
Q2DHIro69Iqdf1dI8uSFzv5ya5kwi/hxLlvWmZ1GWRIzsIf5MI76/Lyc5+dwfWqLGQVsOz3BR7AD
00JIcIQZ020UlCcGNHREkTaQzoqvCe8lZONRiLL76BCJp9VWDVwi+Wf6d9J6ZIIrsJaW0FsyGFdl
+O84KD43nv0VAMCdW1bMdvAiVhz8vNVelBASDzPqdVeqyrEQJV1zKZ0txCmyBU1IbIuiNnuBTtMg
4SQCNUVgjl+uA986k9csG8btF3Q52qRSXmw79nPulm7Z6Fe0rbhvMrHfnBw8s+VhCpx/2GiWdMop
iZ1KaUzNsOdw8hfa7rJn3towGpATMtE4LcQY1ZQ+aTDIssElrxx/v2b2jNuw6dPSK9BnXNgaJPS3
9Ga2xxM5cP+eQvSIaSbY4/J6E3afNGTiNqvZ0hcvootNwKXtBmB+9n1w/6aOYO8s8xMch3x45SNS
EnFN9Lls7shTCYQoBuayb2RZiGwi9t910EEx7X7FKTI1F37ewM72Gj9v8Ld/+oBRTmrQkLW+42Ab
LkFfQmFqlYKwen6OoGTkfF01kmbkvLBkskSDTo46fLHUmyAcGhI/33sAR+LKkkLcB/49n4/oCmWx
/Oaiehyd+CaDD0ZzzwlmEfOxK1gdX2wIaBQkIcSQAxODvSKuoj4tecBNy7kZFhDphl+42oIjpc6/
fQqvT2UWzoclKiEjw81yMZO6+X+ljy4ekOMBDCCm13Cp6lPluSiyl3Tw1YyQf/sPoonLGuXsQvhm
3VgvybOWms3DUMu8s+CIuC50f3sVaMCeQVCgmzYU1OX64tAcaDaqJx+FNIm8cZn0Oj9tENWzWWz6
4CCq7KwMPxrHgeyD4NaZDHhs14rSSaz3HXMqGdaBpbAumBuitEjJhQdHxrt+djt7aKRkLpF4B/2O
pWdtGv81yUcpuMxCSA3CmxoTadE/9QsdacpYYBirDbfwNV7LQOs1FdfgjEbe+yTQ8ZN9Hp7vKiDi
A+BRdC5iU9uFL5M084ATN4Sy5Bq8mOPxWsKen0lKfHR/BVcaJNYD8mcBob5zlTlIDWlIGZTBe9rF
eDBMXfsjUu61f4z/P/K/bPgqli4nFlJ9O5Jv3xOrqSZbx+dYhBYTLjM/aMeaDxGt/yRoVM5t5Lvm
zzoAegTDaxcCnmfo0r/9IfkHabrDPnoxo3APzB3FY/RgaMDZikA4eYYcDxlN5V0yggsX49vsq73S
hNagD5pn0s26XHYn61ZNR9TEKcAgyIRv5oXXXkXiyl/HEpaNs3KWCKa3jNJYaNJvMf+kUodWmrIS
iyTh+Q3HT85qshn2ztwbIzxefxfqCcD4jKQLbgZT0GBPjctSqFpItYJBvhcTzSV/Cr1JSjxDGaNw
JoyVhwp9FkOXnl+hri/zIJcWgmtsKeycbneyT3++ySD3Do44cY7VRG7RVhWLyXX3z79mEmL3/STj
0Whazp1Hxvb5VMHLrDYU9XV4wMARuY8X1ds3M5TP/5GkBK1Anyap6KvZ/ht/g4M6oLMtVHf74138
rD6pyKGjJneBmdSe76MlgeXfnUPu+G+20FSJXcBdCgMQUuRWYTSdCWNSX6CQxh4adHSsFs3rxDL0
a5LQlq7gjFLYXVwgxrbudjDQG1aiAqm8u08591EMX/B89mX6hGTcjDeYeD1bImdyXfasn7nNxeSG
R/lPyhoXI9CZ9etZcpK0ObSoIii5FflUTkMwQhHlJ+Q+g7J8kShSl1WDqasiRvLUI0AUNZke9Huf
clJZbPR3TeSsuSZaXsGcHYYQe0x4Rb9s3WlLmuAfkRRV/YOvw5KNmbRvvBIUEpcukP27+Z+DpfDo
S4I33fON04+7xoEdLrPoAWuNf9LcfipPJtXuu2kvB1JI5w2zDgAB16LU3dG1RTh50MmRTN8Iq2tv
NzM7jSHGNV23Cg08SPmcx3/B/Fli4za55VdrC8UJrXItWTVBy7edl3D6smZ6vJLGKGy1B2aDtlr8
i9YXQkQQXV0M65NL1KlxPKATnVhOMvecZqze7jk9xMQTASUhtliLekgdoyub3WWPInRSVdDN+acf
sgi1FEz0Pw3tOEmvbtKH8zCD89UMlz35NHzau4QEMz+xljLm42qB2WN1Z/20pLJVsjqG+8UJceew
zMwhb16BC/NucCTG4nBt35kcCOJulKmgfymrmpM/5FPjLs/gNoEpV7HKry2Kx5DwGPaTlRlWvf1R
rVrlYhfeqmp8jGNXuZdlDN2NN/MO0P/aMAfagt7NX2ZNhwdIXHdRnLuTCEHtE/Qim8Dc885MuyMe
XR1IaYlKskMlJbvZN3k/6yEKWOVycludjBfVA04iMKbjdWrteDdzFTXYmtxJqdWpmWrsq3s3/67W
C8PIjLSnJwOq1QY4v4UxN8dQebJa/46vjDvwINMruy20nmoJBMaQCjwJT9PYlPBa463BBuaGvcCx
JrmBGPUcILUVFpKjDvciaD0tf7iTQuuskd+vZjXooRp2DAmFJscE3i038+7x0CjZruZK0hf72+nd
JelcKPQrvH/XWjl1Q5pWPPKdtlBGbTTl/LcL/OqETjwabPC87rY6mjvRe8PoEC0xHt137mZZoY1Y
tZWqYDlAedm8kiPi1Bio87gaf3aradLANTMUJWDQ2fl0k91O23sSqcqMZTgRT8Ovmiwu7H3yt4Tn
x3wo+DH6G6LbSWvTpETS916GJI+wqwEbC5aSlZy+W55StM6+EXREq4eFxWDgbHzzdQOE/ESai5FX
yci7H2yuWsCEiytdZW8FnNFs7ku4GxcTlDAWN+mrBTTJHL39zuxECOVTfgEIev93hsHVsk65gEMD
p9RqCo2DDpK7sIPsHTtj9KjNCYylZQT3ned1YfFQT6eFZu5FuuCRIMqEcuPfNiexpa40TnVhrOjs
xiuUbH3lbQNO2GO8Sm3L029kKquVrMiUw92NSlSz68pRf8T2Ygr0G31lvvqoZqMK01d3u80gh3UH
ZQ4Ijv1j43BqHDQjuAgXvmi+2ZnFR4oZGcYaST/DcGyJHJq+9Io8s4/OUEzpj5RNlQUPzBjwn9Sd
VdpuExNSukXWZKKwtrgOiHzO9V25srfZe5W9t13OBnHui66HiSAh4EsYkDJx435AeK54DvdDTYUr
MImkQBydk48GEVHID0YL4Hvo1mA7AeIKOhauIEH1++nP3vO0bJ2HFSk/Jfqk+R5arJlMAFCSc/TQ
u5XNCRBtuCfOiJSA8TBrrixnQBDmAB/hjvXzXkc/hRQ+6Yu537IeW/l8V94AG+Uu/qyT3rKQRhV8
OdMldfIwFz5o+WWnU1NgTVY02GlTlHl1i+mz4cRiojohZ6B/AS4iUBfPGlYNLdUSn1A0DkfNfuIx
ZQxjcRqbfSPExZ+5OcshhoaxffE5XhZAMSC2Oq+o8D1sCKEJ0091MkZDYKxLCbttPUGxLzo6h48t
jbfm1LfS0MSkNbuBPFvlCBGpYvWr62oqKyjKwIAyfjZkWAUmP0dPPKlXzbmVOH/hbtv6adOVa7VI
cfRO3hNGzzAimwRJeamgrhO80D+MMcMmmVgYfNsnGTGQJwfV9bP6mie9IeeQMMHTkVpJXGnGT+Sv
CogWLtX8rZ3GEofcBZLSQVsi2xGNDG/Bvgd0rCSZ+nlXMN5IKIR7rdOf75bFPC3EK8t3TrRtiG5G
4GbRW+uufv/xlyvHWQBYHzLoO9SNn/DHhnOYkGN4uLXPffW+/JQyh5xd8YbJp0L9/J06okCvbtU+
zIOr2R9aXyg5DIMjTfmMmjosPvSu9xP3HEkIhd5pLedNRcj7yHGBbrLv7lBrQ4o8TIXUX4w8NZAE
eZS/a6GZEuE/ahdeVGJDpPyqk01lxVPCcs/srq+R8LpaAa68ekB5Sx8xJu92pitFsZ9VfEHwS8BP
A3jzeAYXPKPTw+R2XgZlWzgkrs16WSEfDdIGf2bSuQxwcmpxrtTeQ6pQm+5b72TQH5cB/IrK20Bw
wwRRnwUiR+J8AYg/AVMg+6pctaLdle/9c9E3aEq2Js93sFuHuUDsIZuFUUZmX4OH1ycUvXlWOyt9
02E6ra4llrh0kh24zBiXf9COhKBuR+RHObh+otL5wuiuu9XBMF0G6HXeqvbjFaKcbSzFKzsFqYpe
vLblrCxgkMz0vfADq2LyNyKdKdNZ+44bAaXoTBxLqFXRZn71oC+Wib2WHWCMdN4ZWbnKXXA46bhL
+cnElMuMgImoMQ7TZeXDEdzAPsi8r90DFJHrR1a6zTF7+tIUoJy0BCDhaNdLEWAE5ccNer6c+r16
OImchcTNXJUTD4chUHBUTavTDJPBNMKDhrptB94cCUktzuy5CezZcCubMxEXhw9PhflLID/JEFht
BR3ne9cUYOwGpZ1KAjx/Fs6Zur++BAuPDrjU/y/pzUNBfwKCXzoVPM4nO+7ZVCjPaHP7i0wGD4JK
RFCfug0axX/A8CvmVCA3XvD5Mc0v8YCp4pWh1U5OcScKcmlyfGc+yfMIPPJfO8Nm9wsyXZtwDcwm
xN+08/KjAO5wOOPBrmGEbBfRUkcNlHKrj/u7QFyd3zDyteEAN2QZ+jtaMAN4p+Y6nqqfb8mwdwNo
GJh6jOhZ3XxPPiaVYQvbCyH7lQQSy0azv0HuG0iBIsMyqaAjXe2h6Oo13imKaHhLp50SmEEi0boA
SLkJ5hp/VdO6ibslDc3EHNZaswzL5i5xvWqsgrte20GGfK5l/N/mEu+TUYVfYJHG2M+GjvqNchFR
bhCKcjpPtFZAhumVluYEMO7QtmG72MPfWizPKvXRBN0dduOptgs2lPMB243cUWYjDsfGqtQNWXKW
nRu9jqVnr5VZ8Zm6EIAHqc0i9gZVbpy3IofOgcvSRBSiJ8TSbvOTLIsBiOXLBxNK6v9zj7DAhjMG
TAxwW8TgE3hVJeXmOL+Z5Lfv8lG+/5o9B6/7aWHFGp0XcZI/MK1FdrwzUe++Z1MFAA0oBMPHkqfy
t4jnJdJL3vgjgDzn9Y4Os5oowLvuHyJXgvaCcSpr4yc0b5B9kcwQjyMHgifL4T8uq2aPzDNqhuG2
NKj5j1WLJA77+qW8r5nWxwhOFmF+CJcXh9AiA0+gCRrL8ANapVnQLf0N9MfQsfdjVVbT3o++Jdp6
2L/OLKPP+54ylb2e6RDq0tu3cMVxDgrPRvAMzbXuwcCuoFnqgqfCjGqjKx2tc5LPZkJKWEt1IAdG
O3yzdZjTLxbiZJ7Jh9S08ryAknm1n8LbMvKu5eeEUWoXueAJtcJa5M+AduvKdL5DwQquC/XqcYvU
HHE8+059fWYFhGDqJAVY/O+Mm3/e+PKFnhek+QtMZsncfvYhuu476PMN4EkaqPHj2CXEnn9E/+tT
pVPZ7+Y1BBCsfVOD4tl69tyvwb05oIIcmtGM15nQuIVW3NXndXi1tHWCMr00+QOOwZG61z0CTxF2
LZQfW81YyQlkqe8bphXfzMnYMAukQdBdutvKHLa4nlwn0qrfQg9kpyvTz66OERSd+36J6K812nVt
CUGiBqOHJReY3DV9B0700IKr74pBRTFWecqhGP2v+s3YQwJ5n1uw6Mmiqf3EbdNYRyLHUPACN8zj
+9fpQ6n4tMprNfHF1siA9Yv6GhEhConmE/8BQ0C7O5ZZnj2vWunGP0PzzN8qPIG4pnqIkdjn5IXE
Z1aEyDcEFGXqtSFHLpunMmn71DONPK48TkIGnpM2Z3PDwRc8UwbxcXhpHcfcF/CeBOhBz9pqGGyU
Lt2+eVXU8GLozNLIPR89ly3T+Cpa4sY8+gGHMWRH0o+ULl/YMZGugLeJHUYpKz4PpFHzyu3/ZjfN
ABhHb1yLK2Nx3IKdyK0Bxqy6hVYk3fbnpBIBcYsEQWJK1Zt5he9jHyLehN3s+lqEbDqaKgruR3Lt
x+YShMkvmUqPR/O1lF3FZ1pD5qG2auraWibNrppRjO+iqz8PUSC65NaSpQq/AG3z6UgXuTDZMTe3
U+WbWOsu97XBtPD71SC34PriLChD+S1dK2OdifMD65z2ZRZbaStn2vuSG368W8buBzGdOm7BXFQQ
9fH5jfEiJTLZFCiYdl77NYMiKe7mtJTwr7PBvlsaexqw1+/6DkcqLYZPK53g25QvwQMVAKaL9A4L
F+PdJX6rOMpCRV1TczE2ZGAqsEd1TXfR+5UnRDmzoqd5QUipx//PCYTWsLzu3AWDTvFfs/F3oNUV
uG2m/xWzrp5Ds3wlBNJa6N9zMHu/bl/aUfitILKaDkgvTduUlTv/SBrnO6P42j2kBMSGpX4O1kSz
K7d3tNtWrHTmdybxbJPTnVTUC9tbo6l2O00r8Tlro6IeTre0pkqcMfwy0rMIF9PwTdN0WgFQkYCU
hTY4jn/fsZKAzR45Pgi4JWeHbqtWZcrLpfp/LITF8OYGK+6n57f3xn/fokxRZAOliDN1UKpXOpeC
J9fbZrBm7E/nxBATjvN3epKEzQdC4f8bgNo1pPbnGWjQ1wIYBkBPfClrSUJDbOy/s0o3Sz27ofPZ
XEY/gB1wHxhs8chNnX5V7lhMy02uzxLuVwIVaRDaVAr2V3Or2Z59HW8OJeYRc9tQ1cBxXDJ3fT/f
koinz+LO1otfg9y12o1zRSHCxVlRsLHKrPp3eBjm4IVxVaKWCqxbWqL7v4m2rPCQY6JFbskCG17J
9Kw9WLyn81pplcvxt4/HQJchSmNvShHfMob7Jy3EocOcGbbiVvCIR5shRH74JoEiwOlZtiVn9ZmV
O9JdIvjdpxUnjYgK4S0Rel2sXmTj0yWEZGg1MXyi6joisxIUoW6csiTGdIMS3EHOmNa9cCH+pTW1
DnIIOXyMN5dHFSJMk6z1h4SJWroIrMmhga7lh41e2iZvY1I5U7QfKOpYqlhctKVHpWtvtKMrEqfw
1Zn8bnR7fzlcXlxtYxaI87WYdrJzt3OpGu+wskOniguBO6pCRGGrIsGaqwmYudKUC/eJ/lDL8v3w
InrNEGJ+bY625xydRwA582PDb53xzlbqUY8IgZLYBQgbehMXwG9dRQ34KEpu6Zs3A2TYyjM9ctws
V51skkRHW+sLWB8v3xzqucbk5/erAbkZCrkyBVvr1WTHGbhi4yFDot9FXMysCspRqa8VMo2j4+C2
R4HWsjfB7ioDcwCPUo49JuCq0SYogVkpaJhBgQUd+drvVfvwCoseWm665OWeFwt8wi5J1TkMhQMz
Es6pO23/l0kk1e+arD0rj4VCBNbpYA3renumeS6bRCew2jf6ntFI/JvZn5P3tMh/0wFNmdyPJQBS
Eqy63hPgFCC5C7FHsQq6te9zLnumvWWZkmZOEa9VKIwdtgs0K78cn3F9v8nTG/xXOP75Yyfr1tfo
ujEGABEPJPduvVRCCUXk2wP8+HLzwCwYMxUmnNuCRSxE7UA37+i28UMsfYumf5Qj6rQWqph4ZFSv
nFvC/jEmYo+9rT+Vf75wRBc5syv7ICBKBgZd/8/Rv6pKTHLYgqsUF7wJRxPpGLuyc64XzfH5Eyzh
zETJg6n70MrT7Ghq7XnLWdL02tGOFV/QwbXXNx+iqyIi/WYzzT4L/njn26lwAUYrjs/dG4hrivlw
yitbJCaQJmOMgEIO/DiiXkqRXhF0yCP8P7kO9xT+uBftBuOau+s756iBTan7DsuQgR8HmGtUkHgV
qf6y0HSDlcBA0bYNayyb60yfU/Py9PGwwIKY/OIV06WArnPKFlOJ4kOa8dWA4luT7xTr1ebXRcO6
3E/1dT7zlbj0BKKLETWedynPznpY1bzQwKOzDVb/bQbBcVhRND6QD4Apq4Heo5ZFf8J+ifVTNmVF
yRS/AZLHNcOM5dfUmSTXydvvqObhviC6A8GD5G9pdNxUX360djCD8ywoPR8mFamqU3AdwZYQYgzq
OvXX6Hz4ekV9pmyPw3UM8al+6RIN2BgTyypb9Uv3X7y5l72jQBFWluh8ZnqdMT/wJuyyc2noZLZE
dO+0glEU8seVF3Y8UMXQTKf9IIego+WmAIgYxWJBajdClGuwm0JSROg0B9G6aF5K7sorAOC9fMej
aUSSCJjoe8Z6X6i6mLl/MoAtZBMI0PgD/iUni2rGvswcmklranKhbbSJ7ZiZb+4U/PPenLVouvr5
e2IeI+IKKnfCj0o3lEdSk6YizIixjb4fFw88T4c09GtJNKp4917t7Tnn66LUQBYUZqmX1xdAr35w
+UNGRm4qIT1lUsWXki6k7SxYbAjj1LvGJzbY+IhXCnAAIg+IddpXzKHxFIRL+9kP025uxywh9Wv2
hYD7RTmKWmqr3I9vvTt7YZdfXBJlwQxMlUlUedyolC77Ng+pbzoLQIQoe9o/03cDOkrCnJ/nDtAH
UCZJjhsi/IQT1rNviwkcItBQkiIqhB60Pyq2KxEegUwcvlkDgUVi/GEnDwQX2N9TfAz7JEVD8BbQ
8PFcEGP9KRa0MCUldmlqQQ5GNM1op8RRdkxMYAMwylmxVn3VDGXwJMEmaezL+KZdVoY6bVqR/O7N
Jq+H9EE/wCXAo0o+mMxGhoT7jgMLskVdrhyQdsUUnsUFQCjgJGcTH0FBOL1SElUK8BmWYjH+LPpG
LiBT36qE6YsCJPbWSLw6BRZYrUijhGwDtbZDI2n6OlTIWOfYl2oQ8RuNSI8XFLIvx0W3vXyw469b
RhH5i031nAae+tchzO6KVgcfwCGMspbWRhNuC+DtECnWnrK/bUcliT3GS21IIGgdI6xvF/wpGo73
CTYZoIG48kS47IwZgmi0KrfztEvqlGX7lJZbNKDH/hl+1vmyrTWs07DCP2mZ8h16Pp3b1tpNHwWo
bK2tNzfiQrf4PCSCqOJBQ+z72ZDCRd/cZChNFPPxV1dW/ItVwCJ4Qrlz4uxOUm88CddHWWRQ1tkd
6w352zGpFRyckgKEUjr03fh1Qjl+cXamsV86hZJMyz54xLwReeG2VQg53Zu32T0q13RsFuTHIR5M
aaVFJl5swxQYgZURh3/pP/IqZI1Y+10k99Ug1zivlTgtKW44i9KQcmmZMTUJwwAPwGsuPsVfIiLT
aDuP5v3KkCBQr0duELSWSIXXegbJ0XK/28OBkU30WH4RUY65EfWjy9C+NUEKW06SJefMwffn1tb3
vwuncT/NTZIG77IKLVj3boYqAslskY252ZH7tC2GqythemWbO7ZhTTWkOiVdyughJYYwLUiNlgEB
WDzJkEvCz4TVNaTgkSomwTC/At7IzRuBVe1f1Yomb+oEylcSA/dYz3E0MQvYWfsjVaiOCvA/Wtg6
qyVV64X4j7O9RRJlcICVvqW8l1ehjaFHKUaALUC6h8DDuKiPbWsPPt5ctwgJCSr8/4rryHsuY7Fz
xqJWh15BjgkJbqvSKsraJYZXM62ThuFUNoNFBsdhqNjrMKmQHn1dBoe2E+bhcAXp9+/RN6GDCdOE
YAqnrbYF8fqJlmJIjLZV6/Z9EGCJbOFQfXoklo8Bb0AEowsJL7KLj3o/vvZktfwegrel4Afl9FtW
Z1Gb4JVqJ3Hx0NKvHl/G0xNIAkPjJjHJXYdJIAcCjsPnQRVO4DEI+Ku8IpBGQAL3tgGwdRpsM31K
bxOCOz0waStYO/WCmMgoOH73JRCG3ztjYZlR/oQ7ETsmbLVf6IVvsd9b492FMcv3x+7SC4Vo8T0a
zMKLl0AIeV4jN7qpNxWM5MKS6asGY3ElL1EkPvGn2Y1tsv/nqoAACa6XpOt1hvFDq3eNtgbxCzQd
jDNJuhvrkFRD8sbfAeTsxSWkP6NvOImI5cKyXNQHxZ7VBtM5DIrNostJ1G8gxoqcwBHseC50/J3A
a3GXAm0p7GjeA8aGwYzIvJNDKfatRAnb4uUl6GvoW1HaYYK3wpl0lUT8nIzdX+/qc9LEh6ieHrf2
x9AjzQqYpSegxyTtZvr5Z96KUcP0XOaEnWUOSiKbhv4J7jS9OJnN8mxihUBiZL3WZ2fpAehkMgrC
GSAg4tgIDdHfYvcJSScP8wHcpF4hIwco5q8/GUdiwg18J7lsDUmjTGvPFTQqVWKwfHTZmWMlykjo
9wvoXT3W7BvNIIPCEcP39dixnXj02KA+rZ+T31RWsSWgapYdvmSEChkRJutqO11PjffNfxwC02KF
u+Gm8pkCt0VpBtedMh0J+EiIJzzCmxHvd9DOuFY4TehptqK/6rcw1zEv2OZ6qmT/pZAZFuyRKYt7
Z8uNpf3sAyg4N+9n7WYfdLF4Frdy9XwM6/yZD336ShcjKtCiYmqH/BVZZfijz3daODYt3aDnQAEc
/Cr3T858C5H97Dm5FuoUkc5Zwvek1x3oqYYMSYlND4aV6gVcdAZeeDAO8DSIhaJWqQOR6dE1I3An
q4k2MGLlpBh4Q4bQL2kAfaX3Nh7KvZmkljhoL1pRO8XkErpS+lBkYHMb24Q9imjN2LWCVHgzHGfK
z9N4dm+AL3GniddYuHQ6Rol2g8Y8Hq475FvRRVfg2q85Kg+/WB4oZnC7G0nLXpk5hSrjeNw42nJn
WS8yb3ZfX6ezBtDhLJHktU+ZjEudMuEGHvMI0E6MOyWqYlAtGgBcZopSkgy3GExg5Izpjli8iiuG
weHt0wuy3jurHVLlU6gItQiCQH14XXNLH5NtKzhN5212lF6rgQga6608WOEtDY8GEiM980ACFycm
Ie883XYyeWf1iLLIb6L4hfApSYjTadeXjhdltVdslHIP+CHwC+xLuoK59W2DNqJAEowZ5y3rdAmv
xOggvsPVhjwwvHytuZUDJr34AGTzDSO2Pv9XFGcBcGZ1/9hTDGCt2+OPyNC2I3pd8h7mrZ3CGO9s
kLGa1qfnIbOuDitcf5vHQ5qjlnvOSyJDbxNqBi0AXahT20VypIgAisl75to/+y6s0kz6faWV13tQ
e0zFOvDMSr3o2lW1b4Xh/qJZDgeBQktYsHW5Yy1bpqOLvK3HGoD823Ibs7sLJvHO0RZ67CvDxPdC
U/Bzkg/IvPDvmtPzUGWAAD9gBAt4C62m6FcwbodrptNqcJWc3CATp7BVhqeH97SOYuLqFt9jD8YL
dJqRNUds+JKOv0xkUJtkQNmyzbsq91gixLAWOBLEyHJltgnNRrtu/y5IqPinbWcp0HEG+XPaPpgf
EJRJwfOPIu/lDH7iRBMRTPFSkQrLdhzjUfx1zWBpXRaD3COsuClY/zSzdzR3um7Jm8IbmEJzlywO
Xat/8hhkcDgl9jLbTSHc01JM2ZLYKiLkf9UrZRogkcF++f+RVCt+ZZtWqkVwQu2oObg9fX3qEOSh
sCu/bNb+Dg1Cc8z/PC0aVpcfu7uvI0bkpJRJU4xnWHWUCWO7UG5kdipDLih+uMGEn/hLpHJq6ddh
pNPuypiU2Ar7oqtEGLotS/fBsHLWsuNqbo6FQRuHykQ1/Szwj/z86Mguig/orrpEbbKWOysIPt/W
vzcuN5P6Tm5Kd8dz0p8QTvbTCg2rkpx5BGlKIYkjfF6/kcUDutmcsehgDIu/V57xU1K1dJ7uwD5P
ecHS5B2kTVYmN4Olh/3Bb3kl6jN0WJlhRGDXo56W0fmJkSgS1GewullZGSowyM2dUtKkhPMriXrZ
W8MNCbdIhTmhBy8D/NvUkiBU1niDrlkMIgwpaK9XUOn4rvyopRtlCGfFPFz6B+VXx6Y070mhSLxB
pcX+rs0oiee7vS2dEbAx6J7jPJH3NPa9xC0FglFyUh6UJXdj549DvUEw5bOxUHUrOkSoh6Z62va8
/7UTd4j2DyE52fdoIC1c02xisMgQfpqiv0LuaOIGvbgF7pshe4NOJE744WGgaa+0x7sOzc8ahH3q
poW7rx0ylbQBJ81LdC1FLGB+TTMQpWWJkkfDhupGyXxIIS8bntiQv9JFseXZWdVvu0/9ps3fac3P
9Q6U3zpmwuk1x+YG0TDgtCoBBi7wAKhKlEy6tEMSFE3Dxz7HzXQqxoQP2+4HZ78W5TEMNdIdFwS3
vS71mYhuLJyAOc7v5w6VwfnxKp1lm7dg8ySsYBaKE9fxcD8W5neUuXplfaVbNF5WBh/iXul+P5le
ohW/ZMQzFl/mjUEmZq1kJ4PydF+dXDJqPSXtTIY++AkydZ9OmbcpxIV4w+VVkibtVKWCSvtQ4n0a
HFsjduXJDxrj9mFXQP59+4xN67/+wNOpn6+6UowSsCRZf3yKy+OsgZXOeuSvPtv56ipfMKMt33/v
WuLrR1RPXEsGB613tNlKhrJ8G4pKTgQsWB0kMQcEscoT4xZLQkotSXq2vhVN2lprk5RyNadc/LVV
wErFk3t8dU4HodO2OL4VejXgVr4xtfiyFnWANhOassZ2eur7GvsLDsONaIKPrLS3riR0Xe+NKaok
AhRpCdFIj0vtnCumYDQK2dHQwzZsQRtC4P8/UHLb9tVYje4NjZeQq1f8bT24O9dhjxXGt/2f2zDD
rVNJOyPlE/48I9+tbFpVNmjcHMaAQElmRL4iNp8060a9yLwYUkcXqSxoLHaJLyvYXUPuS1FC1ckQ
Queesp8IrW/L+hF/J9JXtZLI4weVfA7Uqe5CqIhqVrK5rify7nPFKJ3/7U1fXfdBqVoKYTJ+mEZj
ELvp6gB+X35//5UesuZscSELYBlJC0e3rWI/U3dWvO2fS0b1jEkgFK9Nd5vUuU/yuVTwba840vzK
ODh+VfbHfVjuMKXXN1DmZpFLQXsruTEHvxtFgXfWbkFMXMadtfnDwoZc9eWKX2shW4rOPv8kMjlO
0/X4ViYsv61Qs9YwOAWSfR3fV7UnW3129t3GybcmCEVkoltQNuOdB+jPPn0+kGoV40vmOpDXhxtv
22FFmfoIi4tVbWDXbp0MkHwaRTKihWCaygk4MV4hI40U0qgbcBnfoRrTVK32tA5QTrHQXkCpmm34
QXODoB9Dy+1HmusZXvTXkcapdBtKADMAXpqsq2grBtlyf1c5GTgdW7G2JmPKELXC4S62Cz0ymO9Q
CeqSlpCMLqCDwzKfQ9tY1BcsTg5dcVvtXAqnehRnziMzkpGIFy4kx5U6SkGugZI9WqdsMFBuJeBV
Gd2j2tBVFPkPMcT7WiJ568wQ5QLJmF3bAGoX4gaJ1H5ha5RX7ECGmt4bS9PW5ln02mATGD2xY4JH
0AWCgdpABUMEag8bLisshCQ7iIYZtyOpieDUTKZRNUIZZG9yuX7Up483YBbmeJQzw5hyfe5IUULI
n243c0RfqmgQ24MIbReU2is4zvHNlci/Iv+rCTAQImggMw8mSehZv2L0XDWDDfPUFvS4Xy/wYhOm
UpIRVCoH2Femcm8FFzbJJydRTCYUqZGO7Zvt5GYC/42l64KuVWXFtFprzSmOoVKWbCQaHYrgXTs2
I5ndSVwaitxvPXSnD6w1BUP4yvFMcBqkpyRCV2Bn+CIztRBitJYsPqeLZjSUuYABewMsLyO64DDg
IHzkEqijtN6OjJ5OiV53uh6roF+C7rV5J6hZjXx5g5ahFS0k5hfL5JXGJeBCt1w1tvwe/ecge9np
ZhmSWm/h60JG2v0m5UREO7KNua9YURjmxMmMxlj0QqfJk9IE7OnWFUFg9ZXHRRliKjS+6Quwmf64
J2EAafJd4uBq536oNpS21YEu9XYp+YCjdz9IcdQpPVqHdkPukDNECY87nhovOFvMGJ8mfQ1DgudU
Tx1wFPLuUSq+tWtbTeTVdxxZEv8fjP6kWd78cAqyrsdoo9R2z6TwTCZ9rnCR03mczj0ZT1sq/7en
cznN7BDwxsGhgdRJhp37/Td4dFIpHDMKh8nRvTXnCj38UFxLVZwB02PMiLTlixs9Gkl+/Egre3q/
7YXqGEamyODcQYcJeGhyjJbmKrpg+dj8re67TmSlt3msYHckUwPRpke96+zA4HwF8wmGT2eNsZyu
+AhEvUkAEMqjnF29JskeVMsG7GUqzqWUBGs5DNpbf1rOczoaxSgQk6At/L0fHWEovhmMiFJtumAc
GiaI03SKCpN/jIiiJt/8O37alJNuBQcyg2Anqw7iQs1LWp7k89yVbZmKy1xE5idb8mljN891uVo+
t7jXG+U04eSKLoBGMcA6TDUOeV+lSXOzdCBIwhWVcYdogggofL4uso3DCMmW6Atf8Cl6e6wTQapv
AEiQx6ql+jWnxXyQi/srkBh4rG4a4UU6+Ui5GV34ZWfzwz4BPnJFsFqeeMYn9zcEIoDqeuNtL3+C
KpYS79u25MeO+O1iHLhJD+RDRoAluKjF34tzf2abvOyUP0PlCKj87ovCJCDZt3N5hdrfJrGqgfQw
dqToOmlBP1lfqt8P+KhmwaE6juXph3Hq9oD+0Z2RPKUEv17Ea+MdUwowHolOZugSfN9V/UL5mXgu
hWp2rWPjiveIRMFh19/hhAp5Rqt5XixWxM+4SgSl72L189vKpPWa4fBAszgKGqMiPSyOuDFP6eSC
tkQiT18TJICzesd7Pi1yImPwYuekcL0NQ5L2P7zsVtEy+rf6tqVKfg4XXmdhvgLHIiKee7CNp7DH
4Zv+dCr6ibdygYYk6x2bDdSr5ti0r5PCxPyXBEaw+2Oka5QCM2Mwe7jMc4etjApWpAJHff3i7+5P
SyDIcOCVxRTlamw7Z/PFDUANNC/5tPup5vDAninpQ/8UDkQCdRkXeZlzfnp2uvax6rFxSgUZsJuZ
kMwhJmOxXMGLMs5PMIs6cRcoMCwfyxm5VLZwsSOYQQm2Eofyeh0lGjfP9BhS9DTcIuSHLE2B+ZJX
O5qOOy75pmYpXbxe8hN+rAaz4Dw4LPozYMREvsrO7gQsO6ASCGOMcynLoqXaJ43Hp4C+EhwTspS5
l7gQY5tEjxnIG+8enO0xzrloLbfGla6OTDYbctlPF1fMseA8NaQbqfGyxJjYQ50dY0f2V0tYSnsN
M5tXtsBOKh7p4VQ6EX0Ujitc9GqRkge7JXyQ2O0oSAUZJdm3A4j7XclGcwuavWWa+zTRksQM2Kfl
mgsMXtRWnsf3ySZ3e7CJmc/3OMVH0tDxc6pMC1xWJvH7c8rTpSSIf6OYPJwIukIwcp3rdhqJPr38
2LZK0VejheOMWEEbDa8A0AsJHG2DYpzbQbvq6uy7CtZLxnOX2HeMbd5h1vtJF37LQPeKh01FXFA/
8DyRQVuD5bhsFt/o6oD2cM7optZpaMbwHcFA+GjAnMibstLtLvf5XblycXyA8yyeW3Q86f2sqr4m
fjUVW3TLlJpFbfnTdHtyIAA8sDPdPxdRMQZHBitLMfyW4sxlGQx3fJcLoZytc9/9MFZB+q1QYMc1
o7psdK3pBAwWrAlAjAeiyLrYf1JYFN4OzjIKt/sqNTmlZ0eZZAi2gXUi1NafUgBrrnF87vXqjRf8
TFCdh9BbrahWQ/xDnRDmesNQcPjfwM3TMvVkUxBRo+psMdznZiwNHo0LSWp6uKXHvJQaphm/BVJB
MxviEqQa7lTgoXqjztt+gsmPBWgL+vAOmAsRB+/rJF1Fnkk4v79UQi/DhrJt92evGmKIxZjv8YLO
xNWQosBHTx/JvLmDKeJ+3eGSIcjVuG4wTwdmbnfLp4LabfQfPkGbT0k6iDUeiCfJF6fNBtTRFtH0
n/PBB7WmkjsiM2UD8P9lmMT7UhurMay66AruRl5/Ju/97oJn2xe1q6r3l8s1cRc05PL160JDjmI7
+5pn/rVf5hBlrf6HPfurQFmjbtjytEzu1xzNlYGlcCdiZ6vMhseKQN8Ex2WmQ0ICJiFlA1Juk9QO
fe8DHdD0oYmidNXigEL8RJWgKsqaI5Jg46Zr5PoyrPYOljkrpbBU3FiYLRLYWDjXc/MkD4nNbzlo
6uqbD87aJhBZ62nb+6jNVQskIbjP+ujnz9SU0JkmqniQvaNuu9Cdl2ztiYCo08jj3WuDsuctkEsZ
LMRBY6zpwXQ3NkkHMs7QzI7EgP9Hyb6VbwUNINWzcV89s5BmiXgzMsX3ZL7/Akjv1JDKowoaf1Bv
bcfFOLhsp9tSj3XkNcO9D/+MHu3Qwxz5Kc5kITRdYslZY3XNDidv5g3bu3d9L+fqIsk3eJBzH8G9
QMGAddqYKKG17WkrTvz89Bz5QSOgApYtkCyT/1T810VFvqJvaqTMb0wZSOteaKY3mlyV4FeamD1u
KwwbjQkVvXYs/Tow3L/9TKdKrizjGi27wZ+Pq9+nHNBi8JVIjYjOALzyDi5ElDctBerhXgfMP4a6
ExybFu6ZK6B4P/v1pWHOiBmt4ZWHjgc5E7ansj64xZbWNsAzHpTCBDVPh+39l5bP/US4mHrDpI2p
xfLyNy+DzKGg8jPSUA+0/E3fVcKz1upIEC18B3+RFXrpiBr9K1agJn3f43t00Yqu6DYqcLzBn1pc
LbQdAPR1kh2AyZhqzfiTAd0+3gYLIaZh8NZpOxTO0ZEYh/7rKLssy23YwpSltXc9L9rFwNDkl2pM
oac6w2DVFDqTO6cqofhlIBMMAjbtiQSbEs5x00ouxLzexlrDlvN0bNJ3edwr+alwpX91TdsqZ8OU
nb7e/L7UAUo+/WsTRGxcVLKNmbwBPIWp9/+vLjfY3pPcjY9dAuzgPaB/85MXLDfVi2JsJ5WNu+Az
JVLh7L87DKcwCmEyQG8JTNL0aEHH3XrwSKEReRoiFvxkkIwHCW8/ZgXUWfgO4LqjXzVKkjQ45vOt
4XvlooKiZGVyqwFzhFaDnsQp6FdabEiojBxeXYBby94pcDsmdKvzYXSN56d1uw4N5ALqNx8LIlk2
uvCRqzwohfCsVnoYXitb50k65eh2h2fuZxF4cXIRt3ZqMj7NOfcD5tojHmk8+B8XrvoA1fA3qV8t
8rfUWz8mc0GF3Rfvzxavw//P9Aa5vXPL95Bsvxf0hjlnL6cc3q/dy6RTTYn24W0841T00Y7w+yqs
kO615HTAW4Yo5qmbO+jqmNthZH4KZBMR6rpdHYLfEKP970NMdnYtjgv8eSB9kHwTsioIUPKGnGHu
ugIotxLZQFkO4lHDgdSV0ohZSSoh4HjMZp/Ff0opfki/OgTAsxE32pulXOVtrQou/OdlXEbRWNZC
0B0ITLc2oYiRrPlH3Z+C/iyJH3Ujuu4DRKdzlc7rn1EX1GN1YpTZluvYiD4P6PP9BlN5Dx/EuhPU
CJeePYse3nRaOlTsWtifxLAtE1PzvrCn/Q702wq8t/iy/I8ik/Dma0TUqfODBNyemes0dET/iT+Z
+XSLJ8vIS8MiVA3MbjodCmMwShYrnRaLfDSLE0VUoRW6R6opSinKJh5SFgRmXxw1M0K/EPeWX4ZC
isyk/hvXLQnjBk/9wvVu1BWXh1EFsaAiTRCR3myKdah0LZmtoOzDbe235aezU3eHof4TMVelkqlg
O2qPm8b/YcyMZrgI8IjmSwAGv/KET14k7eop8KiP2n7/6ThmMiOOGLR+C0qdI3kG43dO6ephsUKk
8A2skBD/OzKeR+xiEAIbaQ16vfASIB9UGJK+bd58t0/aeCW1zMEy7fvDS5a5f0Wy5don+yMYOVap
+Cgfzvn4z3pLabNRwW1WUmq8f6VuR+PXy0fwsBgWAxrhNpoZL30Z8lvskr4cIv6mhzd8XAgbuViO
TRdOax9wETQnNJusAza/cm1y/fZy6x/wGak7ZC5kr4o7nlD2Tlm2ktF3dit3qZk481Z2kBbnqnWY
A7ZygdZCjrW3K86IxYm7ZczN9NpTSFkA2DW2aKdItYXDVVUWbwVuXrT9Pd4B
`protect end_protected
