`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ajag644NzV7eeOwulANUHnHIVncRO63vIG5BRUvWG/0kb06bmkkKUJcCsFof3TjMNb5WRe/rkxdi
mGP9s+Uf6w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QffREl8WoD4LFXyaQ8XN2eQXUU3ddTTkmU1ymk79MZ9ydJNyBEu/FBcgSKzXd5L3FinrARCxtwfZ
6kU+bPGfomWbShgSpgmc9kxxD+K1m91r4L/vJjH3ScGeghwCaym7WCQtA+0ohXYoV/g5AuTBE9rx
STtdwBiHYJlEUBzsWVc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wGE0Jlu6IFxO41XYcvFUrqPFpuNRffttCy1JM6cn3D6ym0CHP+2DD3iGjBGVJzLUV5PyIsMo4KJD
mGY3ay59kv4yi/j8rCCBPp5r0/UEO7J/DRmmrnbhSOTtWl0V8eDCfMkp73RyQnzIjOGotVFA9bcz
F5XveZbUqf3PNPrJXaqFNFuJTVIp/1sNsoJ4hxjZCcyzmk4gKS+mLzc24LBSPsDRICtw9eaE9lEd
D8ly4nqWbVnxdfeWs/0tRIwtPwtLs3PSSjnUtXbXcglm7bCJIvAd2D+PDB1UWsQQBhHxgJHFci5y
tVvdDl593ti8j1dWfoXG+In04f98FWhtyNGXKQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xqodx2rIG2zIju0kkIhuk93mdi/APUQrNKC+dbiLThBr2WbvPkP4HZDP+c0EA+/xNdPP0KSEKDqB
752DUTvelefgGY1rc7vJQZeB4ZmurIIYYvyBgPU86UxtnB7FJ8nlL7Z+CYPd+rZkixUtfDf/0oAZ
4kdV/rtPi/1JHL1vKCI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dKRS8i8xlok3XBetuJG3cEuVp01RE28DyBPkNoFDdgCKnyFFSQU4b+7qbPGftDKDLMXwU43fwX1I
BeS2CF30SRoOfD1U8tYYOPNh+Ke4HxA+iVrfk9XGcktGyXtMZIM0Do5rSKO5ujzHxmoX0E/MTjKW
JiufEYp/RPMgeDHrPB0OEc/pCrlY2yTq5j6Myked8WHzYSRpjQGeNDgm+lSx+Fz6iTt5lvlDGGgr
dDkm10pFZjJG5Jk7JhND9MMWTXff40WJztWydFgKnNAC9U9ycULV4EBQkn086cnIOWLNVcXtzZ/1
AnLr30QESDPyOUFk+6fqeg/BcJkeVpiM4DqHhQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 34944)
`protect data_block
DTCw9bR2WyQiGuWo64yph0M9CBWOsrMZs4Ft1dAalhwJtkDcTeLrWMN8d8dXg3u1maMM5zM0SmMp
u0LP6hHxz/DnPyDml6YHdDN8Jneox9jZk5sjAAwumpdoi5HdSWEvkOaISoB90lOEJj8NmUGGSQJ5
W+GIEBpL2mFT5KJX3q23wTzWyfMAh9jVoP11h9z/g4hsMHTgsKD8B5Z3fouzdV1ynKu+sig2Jjsq
MCNNsgRWk1Erblv2NhwfztgaVRuvakKL98WLEMB2/Ht3aJ5ObhoCH5bUHmGtl9Y9IzknMI4vTXys
MQyR9Y3AOd3F4toybZdgRu5S+wTCu/GTK/SrMfPaSu3C94850D2Q54AQdNuIaL9gEemjwZD+sYHX
IVeJl1bvvAvia0yVuhEYV3PivMrWtyyYX4IaTd/NzQ7oniaNdOdfZkYMrTGZ/TYr1rCzUvKilAre
Nb/kSpzxToRd67lqRlR3oh1lxslhWlhQFkaxc1jODGagp2uyN5HR3K8+zrt7exmkxF2bnZF6QqYP
MOH3TLwVBH/3Jz2F7TSWcr/9ksVKx2NRXTT/ej5kbu3BJ/p8pmI73suLANwylT8Ej1TB5lo0hkEG
+wnW14At52iGke5xZMYDWoNA5uFE1MhiBrs7P80PubZa66V+nGygKM+87O/AVIeYDrdkUTnZmkdx
bWeRSqXi9YT7vWAcasCcJpiZvNpBHl+kB+tS4zIToFSGW4o2GJ4vcFHeZG5HAI/6TMoBxsq28C3U
q7vaE0krcfrJ+eC0siXvAH2MgTvwcOjnuPrwfRNLtN0GaChmXzTcMUecJg0gQ6n9Iu1uCnOik+Y9
7Xv1QtPGDVmlKHKWoqgj5jrw36/kGn2JKMTqTJ39s4pFzMunAsMYtf8dj0g+uZdNdY5eEuSuEny4
G+KCFfbVA3eSVRorsDMw7v01tuAEBqzAoDdvaaDwPMoSXRyBn7/Mp3YFwHYEkpTzjQ4vnQiIw5PE
ppl9Y8YdILUtcku8v+mUnP9DxCPlsI3d7jCOdGCIKRVYpWwGYPPB6VHtOytGLKLWjkuDXC4bS4tS
peJ3QSskKSgB+KPguRwhDFfYAaTTGckkYMakqQ4fxqR1lOiwXz75qTVsFzVtfLcSvHzKI+w3dAbK
rMv7M3j0Gu+wE5AR9WuDKEW3v2v2Oa3k5yatxzWshl7g5U6j8go7tQWVaH410Wryfm/lJFOblLmO
M5sLu5k4ZxribH8yls5wzpmdQzZ93pmOrWH4qHJDJt26ShVay3Dnxar7a7SRTlxxtJpiE9tq+kJY
IgfWcPrSvq/Fh+Fm70SHRkFLCTX6qzxzWV1VxAGSDWkahX7PhkHmxJmyQKT5KqF1a2a7lp/Lwzrv
XLv2bD0sDBgg4CXRJWedL+bG0zU6fUwHRWrEUXAbW+qhDq8//Us3feuHGHaDYTx7w58goodMGYZJ
heFKW0hXwnbG0VHtNK9/UBlTs213ZN9IF61lpGZ2ggB12JgL19LSDIcKRt7vLt1qMgzkduqQLP6I
+PSm3+NkLuAlIHoLdZjn0rm+obaTSbXz1rOlBcyVpFDxPdHwiCRL+TLonPpUwry0ZJigNO6HJ92j
/s41iEhMxn38S2siomug47PglhwkY2pdzm98onNgr0Ps4Xx0NmYBhqYvAee/XCPijw6M4V4HhznU
2Wyheve+Gm8QuuzyJAGEZzE4u7/p2JAwzykwnWYdAZCmiqdXmYYwtsLpucTutcDqVAVYYe6tOARF
ge5y0ZFwsL1HX954XUadPL44OZIYWv9Oj81Nl9u5+4LogTvvu8qPF6NCTpbJfRIoR90muCSev7i6
nFT5iTA+HFMTy+2pQ0NzQkgII0IbO5MDyM5X7dmLO0OG7Sqq370P0TF82xAB3OygMGb8Jwto4a8z
vtloLE6uLmXh4hXZJF3/jzT2pGoWnuR3YCyeTMy6D4SYStECkXI7cE7IaiwKnsw3eT6u0QrzcJor
1d9n0+Q4rWZvQzD88ik3CcL6gV7nlFQX2t7PYeAcMvHmbAMjnB4MtkTO5J42jlxWz6g3N3bCeL2D
X2LoOWQYOgILjJlAGeYbE8cg54K29hLgzxj/7XEu1c45U3eSYERiyIE7/rarzwCMsfpUyBCYgH3d
H2wXO4rtFxqbEAfk2Ie7bIkpqlCP38vcV6nj73W/4Uw0Wgiw4urVkSybtHmKiEWD7RKTJzgZSbp+
hay2nBrfOA7PINln7RhFBBS8ajBSI8vpnubdzzbL6KDfAZGUH96caJ3hSo0vaSOHUgtFxJaTG9l9
+jX/dPbjiWR2h4nO2E+R6nHNMB6JWrsxXC2zJ+SJt4fhMclaODaMNYoL0Ruq+m2O98FrvLgLTNuh
3RVa8k+9gsLdDNuUZOWUaN5gK2oS2gTUzbNW/HuV6QNH59LLuov5JYLuowTKey7Mub+CjC2puIsM
h/MtvLzBSUHPSAKgD02OQMtjBt1ZKEw9Lxq971j8fDwH/bbqL7vgXOVFdhnFRzJVqRxpId2YHDUm
obR6ja/3DXxDAZDNTYnFS0rmzma2xcs1j/oTJFto4Dl0pjjsRNE6WZDv/kOtFhUWDWR5bpeXqZ2z
mAlzoHlaY5f/HBgsglQ0yP88kILpAAByWmK5JfR98dycL5/ScQtb9kS6tOYbI0e+1SxaJIgcT5xH
Hi1prphKTK1lLSkS3wyEBCfH4OyRd0zhHFR54C6f3JN8JB7ueCQe2aGLSLizlhZ7dqR1WZWn+oTI
yOQS2yED2wjGUMhVMTxdftl+wP6+Tjs41YdSl2bURrwsvHh3dt5BbAYqZd1dfY/zGUsOFVQ8GrlY
8EhdrBYFl5sAefE+ZNAVa3Z98meCltbSaK6qcdN6+9Cw3XfAWD8kZSyAs3o9cfu46UZrsIn0vlRw
F+i8RSEAXklIXaNit2wX4YzyymBY4uASSBjkPLq1nDowN06dHzSXZoWZiC+GR8+9OewTe73cgBnZ
9HyopMJBlvRo5XwvUBkEYRTc1iB8++3WN2cZB9Pq1gVVgN6G7Mw6oUBbnrHRwvF/Tz9RIml9Wqf7
5LDPoxtWDh0WN7J5cxpXO2jvKb5EIjEvbcjctAHXLdwcSrEoN+ADtyanR08/tePe1NHIwBUWJi/A
HJKu1yHHst4IF44N2ypcKTahUXoTjmAMmRKWss5PAMkEnwvj1LfdolR5sYO6jz0Fn83QDJ/MoXpO
54ksJL/+b7qJUPMlPOgymwPoe1r49kBNAqzrYlGd1F21XQ5AXqCpWIdmnCJQhecDZrvIBLX5XmQ0
YrKx/LjLmH3WgBMKZkNnSBEIkZ4gR5zpsWVsmA3+UL8NOXq9FDfbGTKfTxsBrw2HhQ1fv7N5R8zU
o1mf9no2TpqtrpdEgg5GC/456K2XMoJngp2+v/qvK+Y8BoZDS2yzBuACr4V6qthcFTQX/0+X14zy
b1ZDwSsEB4T6BhIjsEyNfEpOnkuP7cF1XYZbNG79zQYTXLOEZ6XRWRgQYEv0J+PigYUIHYO0s6Rf
rI0o40mEfKdkXupKat51e1CHOOSYprhx2H4qnmE2WkXHoJipwLVGnd7A/XGx9mMODXhCnay0qyZM
F2lyl+zZYXYmCtEymxc8Apxvh8bXmJk8g+juz8IfrRFnSqFPg3RJmO3wdxXFhImzN4qqIOGdiJJC
xcaRZ2m7IM2Ux5I0+a2xGcahRgyy9YTXDFyLYR3e/C9RNptX21aDJblUE3HUH9d+fbdQ2oTNLQBZ
UEjvx+WYBO5EIP2Xg0nOUhd55ab8p7RWXBNN6VKZ6ebFYVD7UtnAGPIdAbBHYbAACtksDLTa1Qyt
rsTm6toG3+m1LfNzNAvyK8Ln5j/CvrdznlDjIZ+OnF7eMwQQyax1mr8wuJD0PjYPaLi4CllTi6xj
U108XwiHNAj8ho1HzOO3FCkNehST+35k5xdgJiM2qfWMCH7ZpnA5oYdqjx+LnRrO5LnYd29yNoGW
SYfbqcefLmZ8ThwBqAl8VtRbuop3v36w760s/59ttBiSgrLFlcL+CqATD+qGh05PIyF3x8kGPLTl
VUE+gucDsxWiJPWVB3bDHn5Ww0QotRa7o1fsnaTBlMOm66aWNV/D9qPhhAbPTBz4yTTEyIBqK0rZ
6iJQe1/vbgfPCzVovvJHm4+duruV37EQxI37OIY0EDeOAjWoyzZx6JRE4qnT2m+EJn0nJByPPmNj
eiCCCpQiiq3nqBLRrb70+a7VsZCVWWpNgnw2w8Fp55umtm2IkdMMmkH8KXvMC3xJTmk+5Blzlmqx
OIhMXE7bv+pxPkty5GwGW9EbEsJcHGbPmv53IJJDxIswuDcbvYSGFXczmYx7BFwqGtl7YSBr6BzJ
b4Fw4ojCXCoZzi1yKVktNz0TaKzuxcNQprOL4ZAINhqhPizVL/HlTVXgAEmR9aQdp1KIbzve+tfg
t6I0ePKTTiNp07kSzqPGZ+ME0vMeRy4h4Dzdua1L9DYtdRYpFcrJSg8KbMWNMBS2pnq8rNJzAOuB
bD5KDWcC1UGrVL2Cjs+ley5Br9D/ah+sce9hlikbnSPPw2HJjoBO2Mu8R/AOKG7Z/3EsD5RLOCPA
PHmg25s14FPIkikbXTKnqeXzFv/33w79No2EK1jyMb2Yho5bvvjym6Oc/jPtwWCXUS0TS30lS60H
Ur8+8K06RwQJSn8MucXiH8t5q/EXkC4AA+X+mubEcZRSC56ljYeQJ0Y45izi5Aemd+9BoUBPjAMC
4Go/m2mf2By7pRQ15Vj9vUmEWTfKkjpkDsRS3P6LuasMZYH7w735IISNs8nzGyt892SewJQ5FDl4
cNQ6Iq6rIABRPn/KgHzxUOVvWq7ak9qTSrGiW/zetp75TU7SIBwKpBNXFOYVjnTSHJ9HUlk+F87A
vVKvQSCmJgGCaLBp+6udWLvdOwZRKDBmnB24ji5o73s+/iPaq3MiMmW7khJCq0Gy0axH2kw6p1Jj
LxkH1T1lrhkgx3TMYWHp0Ph9tdmnK35U5tfgGuV9zCkBM5vu5uwToX43oXMh6HoA/uq01oFQoDyY
TPwJZmxVJODf8ZzZacdSBXESNtDWNE/i4pEGgyHDA8zFl+TJBFBOY+AhEFG+7/uAFPnt5c4bTMlV
k9Xfxok84wUU6lqTZCnjn5giKTTSj/2g0pNsAIw/en7V3r89AiTYayqp3WGdVvlOlsFFVKvrA0A1
j+fqluZCmGsErbf73eaF4IDLz1UQsCL2HOfZG5ybuXFM4Z/bGH7RMgaIV5XXpnxtbP+fnDTkW0M8
FyLjMMyuYfqdq4NmK58baOV2hkUEU47dWcpMnMdFWRIeakt40mKBxBrzti9kQAqjlwx7omDX9dwc
5zvkj+d6E8qjhtlMMofhgDx7JRceUxEgaeVO0r4Qs1HM6WPP8ZCojsIJek/ZYyB57Q6O3lwR6Z2f
O7VxlMUJTNp9vlrdvwW/4hhhFGAKrvDkDBg9ERk9oz7LR4MION0eIHLETv77ctssYkWhs34Dr//G
DmU49EiSE/JX5Cg5FF4tvg/+IoZ3yUhfopPyvIa43BmpUPTGBzDzVwojLwsDlFqcKcmgWaksssxw
XcyleaDo5POXdZiY4VxXT45p8O7nOnp8zewYpzDOaFKs0Zq1wrcZfkYK+KLgE2vwEQ840yS0xeQq
PmKflHNPHipyNts+jc0L/dB0TPMri9JwP531PVMnNzh4zuoFLxjrsEbOHXTXacaLDs0G9V90n4VE
uB75q+2MKE5+WHsrwmY68o4ldZRt5grcR2wWLkbkZDLZDF+RPJ2/OfC91p/tHPRDaVXHcUTlw8lb
6KAyIjDW1ilGmmpBOBRM6KKqGVYwdV+VZbZWlV3oOfUmoWQo2e4ui8LN5voxijzvS4fOLZSTLMcE
QysLkvQIw0ooJky5yRve/Potd5UzyplLLC4Jq5qKR1a3/HiBJdsqvFIWjIR4YVaJ4E4GZWF0HzgW
q2UZpn3GVPwPCO46WBv+cq1pJ5k73jH82a2oUZ7IQUp2KhTuMfkzhUon9YMN/FyILcgHVSk+h1xB
uw33BcT7YAu3QipBkVD9PdAJ2ojl3nHn4dVYkAXCuXYsB31TE5fW1BHlxPvhId6TLig5CbqVY+CW
LmnLmRllGblOx5Ze5VkKl7XwX7j1uIDqZBKJGEN0IZX3lQTnziigh+4W52K77wBYolo497gr39xB
1PQ5QEZYAifAEe2A4WC4iZOw842gSG+Y1B9F2dSyylNZqHxil15OCNLsFlyaDj+N99NR0LCqIcbT
4+s25+ahcxgqEQMNQpjBIVAb8l1UCWhzw2PkKENndAENG1iYL+5WP9ACxewVf76JrcnhtQAec8s0
U0swrbKmhTbEJs9XwcWXfjv5iC7z5xX1QR9oFbvrLCktNWi88QxL7geuVQ3K+2PXvuS+xCjMvhD7
2/2jm96KN4pGn//AqSKKiUxuMA80x5fiwSHOuajfd0sXOsFeT4GhdtJurtKtzufhUlTHJT+HzsHZ
XUZf+k+Lb4HeONXslwBEDEAuE+bbQI+Dfri5DribVc4mN1kmm4/kjRa9wOiv2M30DwmOVbHSyMzt
GzuUFFXJgy6igj127dtbqeTbO8/k35gTKf1m5s2wzFwLajFf9q1/GVROhPEoi/Gi8EEl2zvHehPC
8Fowyg3xmdX0EA6JPJXOoqBLuaG1NYrQxjZRuDv2m6DqAAkfyvi4WwP0NT03GDIhfYz1cJrvrf9x
RuGW/Vv6GHNqETglPircHz1Ihh8DyMZMUn9Awow4M5TNM3yQg9rYyhnxkN5tKMJ9DomHPIlLNv7Q
JsNoJMLe50SHjQH1+F7I5In/mXRpZm27cM08oxI4bIu1CLfEt5zs4iAzaioUMqQNKTRmipM0ROYC
lPXFEKG6ceAV6dyUFSi2CQqKQUFI/PfKF0biYl76ZF5XFotatrueTQRcnJV5IIhfO41sdmhj9KlQ
xcA/iXZqzL3153wO4KHMw+3LCHzo2GKWEjU7W8CkgPE4sFEbyuUAYrZPddniRurpF/xy8rCy/cve
d/3zAvrXioznXy1DMH+yunTO5D2AJs7+CVq+cPQ1LuY3YtMmJ9qofmlrRik52HH34LLi4Zreo3Ao
u3jp/PvnlpYNSkQ26A5TFcIDAhhH0SGFTRRPsIc+9s62wvdxb/YLU/QMnDT/jcwNae3ljWvXebov
mnnaXBbJbMD7Od/DThy8OZ2FnXC+QqNCYBJetpdQTU5ZlUwH0djl5O0L2n5vQSSpY6VQyvk9q9Ea
5QsuT/LxyCu/2f/hXf2h0b35CgYHV13jmG+/7S9BJcE+Bd4PG29gxV2wTf3XsSpRDxLuB/QD3d+j
iYwuTMGy9KEmUo6kbWluixfW8f3p7kwekmE3VQaDHoLG7B2tsVn9xMaZZ479+W1N0L1IXAsQMiGY
sigZTOd5y0K9kQn7yKTPxdbqQfx40LESbzmfh0xHjmGNDS3iCh4IrkMEIv8VSknb+E0kiGZD6IX5
VvNs2So0m4fAgdRvMttBV9HZPt/EP+5rLR4scwx3QgXc3qsGYGNKag7UL8fx07v9FVwC7S/DYb0b
srJuplj5tz0d0E34iSgSX4Jqlv00YUKaXzlDwa7p1dWdAOXELvWDEJEw+QtQzu9edrDxaLeKuFIG
ScGMr03ZMrLL4hgyebFznt5vUXWIuVjgJ2VMWMNvP6SuVcYwQIJSOSJSG5BWZpnG8wsh6yOduiaM
OYGdGryzdJiSLVQMb4CPtTNCqVpSouHHgDpkJBZnhoOlzC1osCfxZkXn4aJRU1coxp15nd1iJU2X
AsR6MvtPqNjvKTunfqq9gCrwBgtiwHVmkGeWAzgSqaAQYHhh8ZRsQkHPxrE30f7NJO5kaDvb4v2m
lN4zk8LyxvszqSox939rq1SPEPmiOlJ/ZuKlPvF+JBYa8p8E2XFTLdp8n3VPulgKRHdRalpsLgJ7
ZUSP54syiBje7aVzmESWniJUWJEg3I7zW1jbjN9EbJRHBCzAqOIr4aKuF/LgV8AQN8uGANp6E2MZ
ep64MVkqZFZA37Fa0Xjgcz3JXHX1svqdvk/rd1yObL9yRvTkO/aCppRWQEFzrazms5Zcw7Y/dZ63
P4ewt3w0F3Ec0k74k9lq049H3R1hLzP5u20fhMYqTm8++ZNC6VDCeuko8sdgkwKUC76kWCP6Qc2Y
YRGDwxJ/mycmIvCmX4gGw7oMU578QR8qv7iSwA2xIoGhAlSKPOJ36+Y4/KoJrbICkoYvLM3RGd79
35sA7Jzk+amQNb1WZx1RoToBsXmfx2yPqlEBtxtpFFSWoq6dZVgq0Wj5P5DugT1qb+zpheWaGoMt
2dRnSb6xZYTgCSgW90rDiwVh6uNtZfNRrDGPNGFsiFhoxiATuLPDxWqmpFCrQDvbEHBk6/p6gRWY
AeCHPKdmn1Wb4+LvSx8F2IiPpll1J9bRfsjfsRGSnh0dz4mBtcQ8VkG2gBPLFOU2SWDpNRW4Tbry
i7Lu/nQUiMycPbBqp8oOTAX5U/Kifxbh9kaFOjiJsYkASsWJgGc2Pj8IXYskb1f7iXx+m8httBw/
8O0tIN+ihk2GGhUzown4Ow0R7QBvWNsdcasNgzL6WeoUU4sycDjO76xYYK8bBLwpYkJ0bOD3wePN
cGU9raVlCVR7T0npZVifA8hqlDi3cLXikTF2BscJeLk7u2O5N2B7Qzxu2Jm1+OMol16X9FGqzwlw
psvDaw/+yFQClNcndDvqJr1szCrGFhlixFm8nOMVSwVNgreeuN/rGYXIXf8WDty6fKmeqIfzSnHr
hvyzQW2qtntxq/VcR1CfY8moOf5dFNEJUDBKQRIh414e8dKVsqMhDTeYoy26HxsajCu4dgczc2rI
1wW2BO2N3MO4JBOPT03En0RSZ77aS/12RBRxFEFtajwCCwXcJq9jeZsSZW+hJ13DbhLxjCW7fElf
kbp4TvmLYWk96mVQcogvaCgN8Vw/hcHZqLvTc+ynsYDkjakpuWRFMK2JgN/XeU7vFiPfurZdYKBh
/QiWsagmWBomONKo+xaMvdtNo4Yb0AFUIi1Lv+nlL3vjFdFfvBoArNj0Jt5Z6R4J+Q3ZR2azRo3W
QxFCrqKw0LgpWbBdmiCd/Jh4ArZ1shPeCGfIQPgGchYl6gOwERaH9bf4+4z9LwsdUur6oOarbd7p
ONSqrYCaXmDObGojUKdM3XaVKb9DH3MYmn+yh0v/gvzxM39Jnglewx0eHVVKCOGZpwCFZSQaRtt7
yMuulyCoO/VJRMVFqs0tasXRfQbMeUYbvoI0oqiZV0S8MBRgEX65VA1RS7TXdjXi4uOaCVTlKrIh
EnabMDF2+gYrlqIEB4UK0pxmomgVaag1e7sh06BPpXYtKXKmlAi5whO8ECt9Kkm+wNb6rYO0fhEu
cBz+d8BLrDIaEF3TGotm1LWDv7r+R9ZjX8MiLt9FX0Vzw0xgZY0buVM0vKeXMBuXhHRFaBH9i5PG
FgXlsr43V2hCERjITPCEeMkgsvfTD1PBGC9ZN4UDr1PJtHFT3hgD9uDYyp9uT2+QhCl4pEK/FFLY
w+6e6CmkT3ezKUknugiJ9Q47Eo9PLSgbKvfuaav7FLIjfidJdw3auLV/GCncaV9pngenAenKfnsb
THUOu7B8ulOmozNov7SebkgZ093fGGiOZAtd5zD7HyOKjiZKXhHdhdI9yPrkr1qQmTrtiRmG1x01
Qy4CNrcnEbzWAMM6G2fLLj+Z1wEiyJn92sqrkNgQ5pJgpldcrNgFCh6S1CW8zuRf8KCipcBqtWkx
SSzANrq08f5iwGsHB/5nMIPcs/lgzPd9l8zLlZlnXsvCH1jnGCS6b6GXSz1oqSwWExa3ehjBQy20
hSs9/vZlgKMN3PRFKFiby1HQhSf2n6AfG6ppl2E1JaWHd0ex6+adZRU5tQ9Fw4itpuTllyoII0By
dkJjEX9MkFRTAARhM6vRwZpfZiPxk3Ep/NcB+PHaWlAWRsNdGFD9+C7Sq6kTzWzJ+LLUWuLQwRqz
GelGKRJsWaxUAvQ+Lm0jx5/EcfpC62FHDArbgerruAb+uQcD0TDxSrtDb/f5T7lNnypauUn+39t2
KUIXilBY1zhWRL3kRx8VlvKhGjFh8CfaNwmeGhpx3VU1ttoP7vOCFzT5A+ro8sXrZWz7UHF6rRhn
Nuxe+ou8vNJs39h/q8IAjxIY3LjvsTYsODewwrxBO/WgIkiW1grddWJOkBH8k1KvTNjbFnfb4x59
0AwflSbDMAipcTxDnKsNvIm17fkcX7WchJgpE6BNamgwf3EO211P0dXTcWXaMcPFaFr7oFovOLH3
4Y9SZTKyhZYQNpPZPytcdpc1k8PJwH0BewJzeswdQpruAAPpgN7z1LLhsUleUW9hC4Q3JQBtT9W2
As84ItR8F8u98uTd/Ate63R4DMaRrUB1YXT/eEDCDUSvrvIUhcV55B8Zq8ETTvKaGrS0W7eBEuhs
J3VtX3TImv1+7aGzFT4ZAFXvILl2RobEptGi3sP4067TWOEfBylJIeUXDG3cfYEHwc4jgc4YoaKk
0Muhas8eP7pG69kH6gpni/coqyyj+ZMMEkOlRguSZqBJCuSkhq9LPBUQILBxkn7uSRKABheJ3p/1
2HF2b+uWwS4b01OsfQ+cWXAFqO+xQDXLpJb2QoMplbL44oC4rWPhmpNuJF3fb2YDr6tsqR0Wtm4/
lDIBY0Q5KE/qZss/D9XbuPUSIkvD36GD4FuohZS2AS2ZrtEneaR2AUCgQ3p19ItLvxnJuYAVcmno
lY25LbU36sbLUC723srl+ETBTmy+9apzQbHrirtp8jw2YHyu0n6niqdDE5XyT3+ggMJ57j/0TvPt
cLvj0R//GEQ5ffy0Ji87HC/PAQw094SYxMBFHPC9l1d2Lp+hLV9bCpeymdwlaBVF/gknFwWV/02P
IkUuVMzLBeeZonYkAjmpmOhjVsE1pKtq28hMw1P5Bdwddc2nm2uH4avktLVcWlh0i5C3uShdtTzC
ZrTMxYTspdWRxsSQhxgjYnhAqWZ7mq6+Vzfacbl6xDT48rQyD2LabX6M79jzpXfn6am+pGy/hXge
4ria/w3dVcHqcR/3YO0FBtYAjBhlV9Zx9TEb+f/VlnIBslJCrev8OghdkQgfgRebszmqxwzJj9N8
VVz0BCbJzdu48HogQ0IQG76L8hc6Udmewu82f0617M3s4Suut+H3JjVKPZN/ZxGD6V8Mkv+PSOlF
xlLu6x0IU68r70KfAkZgtfd7My+5o4v5ha3NW4q40YHt/rNzqood57S2BnMt1k25/4u9rxONz3aK
r2LpsjBKdkSPOWz+PrLRG/W71e7GCy0kaGuW2e2k2ixNkvW3KngpfCCsJY483S/gVWCj0eComkBw
TgTKvJTXRjfmm/oapaABYSXHEQS1vTFAM0IhqLat3Y4vMmbQYy5rZEnRVp8LU7HMr6FGXP5oDooh
Yz1Q/ekowNsZyBQ3MluJpDEVMF17tyBj9wREUTjKLECuzVKNx5tCj7STFe40b8rMlifHj0WhGlhY
0JXZ9cZoQi/jkvXOUd5dktl8FeP/BV2YCtABh78mDDeJScgxAki9U3U5sJlmOwuKepLZNNHan4WG
+8c3pE65LqOLfTukc5YfAbLx8BeHmP4bEpe+UAYI2NVtfok3/Gabb8WbE5O23I5k5AfoHxlRypCG
ddj8FlKRlLgcG1jIm3tybey59rKlC6jIzh3YedzyDE7EO2LftPScNE6wU0d0I5e7clTS1luYBi/9
Rfq2/B1Xueqa/QWySWIE2tRsVTEx4cXAvbJhA4I5/4NXcXrmJRWKHIL2ZcAOEVToRhaexP5V4T7O
gTOXaw9LPpOhlw/Wq8YzjU9Jp8HdRkT7/KUEN04ec2eMJfGpur31nNvlB7orIpamEcWK3dsmxsv7
PgPxfBg7mxQOMq7dZRMSytMTEAD32sfm9ZGC1xWyTyQg8L0Uk0DKVnrd6Jn4S5R4yDY97uEcNkJ4
D4+dmFgG2ognmxXKmkDT+qxZ6GO9Rxo3nCe+lUHDUIQJ+gltmAmIDLQAHvNO40P+MLX9V3+H41eb
dnP1Zr6Wf2LA4L0Pbb5tZX4PRLt+9oy24ka95jrgM2V4WLbjyz5REBnI+wMtiRAgqExktbbDmWpF
PiBR9hTOh4C5qnTlW+JWW1UDD2DS2Lwd0pZhlbEj2lUviszkEx33OoWA6sAgIW5QU+5XcptyQ3rL
PdtZ5Z6E5J8Jo2OxcafKvghsidzmrug5KRcQZpg6o8KSJeJzpgnh3jtOprJFGQ85mBQFuGBdlMZk
j9ZixpEz+sQOxQDcNgMTUPcBxwM0gk5oTvpBxS6w8nreUFQsiW8mYMIQmoQ5zDlVWhR1VuBxZRE3
B1+1lUqpe14kGEmbt+b9p1bOKN9qQvH+OHSvpYUEUqHgFYKeCoAAJ5ZXJtDnFl3ZwhBElWsTbzi9
b66p9kciKA+M79aymfLpzXfa01FVxBGWFV8jnfHcI5i/W9BeA/SYVEJz6xRiXb07SdiFw/uC48YN
3cZuWlsx8BGz/1vEIk8sLO+u67fPEIEWGz7aKDwobB9wZh3tfCFj9iNqLdjERvxqYx6zF2ERWv6S
JUFX34riKtQKuUc4qhm7cCZfJEcX5TLmHFcTpPru1jrl3J4hMl8xP5/YOOdCfC/07j+hiwldo8NC
kvVY1oYpJ2EeMxz+Go0Kq2pHR5ovoOKC4NXng59vndIRPCDFY/o9ogJMT7fHhBUh0ZS3VUhrbgXI
1f4afHzF5FmcN/WMReQiWRAwxI6AvkR1bAhBnZTtaTc2SrCQlaMKwr40/jUeoBDLPQeNdYBCEXbu
7GuQP4RdaFZf5t6d1zepdm+ZRz0liJKn+8qJM4PNNgqP1GfKKeDw/vn7D+y6Miw0hJ7rEI56BmkZ
rsVeGYXfCY/HSyYXhjWrnPchHX+/s+dET4VKp6kcZ/ZaUY7mstFEKYD/XwuJQOhhrVnU2vzTkTwp
wki3kWIwXjHC0gt1MdNVqgZvgRKuNoLGqW0Efi8JedZnqm4Uj/zW2i4JcQ1eLdUYn0YBx2zmTyOU
bIl08iRmIKD7dkxLtUD+a2ssEMbM1zR2dpwJVqFT0DIdhcAHOQtF576njX2ssD9EzteZfBO14Mtn
7rzyRK07RLeVOmdZnfKrgS1WCNjBxMADr30twzG5c0uXF2xIRzkJxdFnoWePwSS8xFfYAqWPyME5
SaV1tU089ulSgoNEJOI9+7lKY9oVJblQkt9tsjk5p6xcxHai6XU/hLSTkKVWwZpM1wKn35ieRd+b
sgst8Dpg/KiXtWS3zdf7sTFM59Z8ErHebTAwviDwUY0vHi4liUwgAQfj6VTY3pNtM8HYWaNb7Cad
25FJjvt/Z/5iS2eS3OzGD00OI9qQsuBEj3NxdbDvFD4jaThvXlCbwziijvCUFiVIQVK0CSlkqHoT
VFQwTfjbMEN+LMMl8IP6vhLao3HfOmwtFon7gViIfezVw67iDlpvpP/8Wa56lXDbrbKm1yKV36Ok
YkcLDGlLNw67JU06edXuHkRrBjvHTSZOF9JcYorCr4Lpk7F+mFgKsO/X5oTig/Te5ePD1fn+QiUe
PfyUFYVC3TICFkVkkFj4iLNV7BwkzWqWoxtLZ8UZct4mE+36wKD2cyciYuJrVFhuipHrvg1DDbXO
PE1iOEbzXVIuNTJkvJqAhrZnpqDrRPcPYGPzfToqadT6BlTkpGBZE38M9+fHbMzARIyr+3JCjrKt
7uFCstXkDsL1i+60RQ7ko0anpjNY9OLew+gs0pdSjgp6J5IGIwKXxTGHrbFiW87wMUSx/nbyGOgN
qcPS5dTE/dDYy6tMqcfwyD7UgAfng0Za2nseKXo2GcxMCXau6d7W0p94xv1kJvS+sggwGo7PWP32
N9hTBRY7MGgT6GnC1G67udTuJJqJmkVlf6VuWb2dCwPm41rLL/e30V7hWcKzU3+vptwXoTls2OJF
3mocPJCEgf6Ja12szTFEZENk5dypOfXbnRWeuDKHgVQIT5e0zkI4xBGcLU0CX2UNbOX8gFvZ1IhX
uM2HMjyG8x0BUMzzQIO7WQNPUI/2DctzSQqpH/lKULvQ6lMwq7E4qRroc1jk8OxHQJiHhIVNw/gZ
n4gBIGj+lphcPWaxnp6BOHTRbJm2pQIzAzSP446lW6LV5Lo8tggR0gHC+cH0mssBxq6QSiS2v9hV
EBT+nJ6VkjMjWC+ulDaSaM5sOQlkBO1oyak1mGyGqgQcOqxi1Jl3rbOQoS2al5GCwdMM6isQ6DAh
yYisMnNJmHLCuAiL83A2xV9Ejp+tnrat7lcvDeDSBDmeSD0rddvAuOmSGrPaGWA6OIYq+LXhS1Vc
fLGftx0oLYdpiXa4+r9PHRUt19kzBHQ4x9yyzZkmqXp4YubqblMrcusPwPatAtm3NUuAbjECgrBb
u8JBW+9DE74YjA/pveSiyGhcEHDR3BrJVp4CWpYE6j71KC41AUVFr4QpjWHn9krIPGC207AtxY3c
I+DrzJmYROGwSL4STHmjOKzI4GagvWBVnw/4maEazsZEHPfUpn3h0cPH0KG6vSztr4ZbBMOx8zTv
pkZJIEjsfKwPLPuvIqg2iAZGpvOuYO04+7ZZPZmTEXQjJHSwHQRjKYuJV1M/4dNGhX0z1MZOOo9+
BK+M5tRG46yKcYE+oHg1o1pBZyRIV7elmr9CHd1tCtPOsozi8tcqSM1aaTEryeCjMcFy5dZ40c4b
PhNbTKrbe7HCqjPWnNYwUrv2SeOM68Et0TgoWlDE8hO4iZz95/U5JMd0E57rP/WBo2qf5jNQcROg
S+XWLfSGQ99G9Tm6oJad7Vnf7CyxuPjeHb3We+yRDdPi6NwTQl1UkRxrB4g5AP5DHxDShQ+R/5Ln
5TcqJD/6lOjJBIkdD1NUgRsHsnpTS3/pZDPvaCVwdMeFepBRo32dnS5GGDPbZvuv+e+lWnOByCzr
9Iho5UyZSZtGct5ibSLJu3WZE6OxV0qTkqUxj+gRkI/BTCG6ShShIYdmvrVBBvleDhflIQnxKQ88
Xuf8INvHxoc5iZ1vr5N5NDkOWr0h6nsKDA4z26s6D5Nlur/9swtxn4sAxFdTozlx1skLYCgMQGYx
Gw1Gvl3QLQvgiPduL/lrNgVDePHGocCR/+URy8rXKEz10N/kBLBB3LD0i2bRcLQYbF2a1nQhC3P9
14d/3+yH3PIzAy4qYqMhTzQbDWALgMkHm3uTODs1QTbCZsX/MVFcXi1xrKaGR0BDjqaWxciNo8xD
fo6JUQ6dS1Bl6WiGLPObGwhqz7Ef608IN6jBmVr48ij1bK4dPabBr6uW0KEr9DhOw6JvFS6am3Zn
LmXcP9erzxoYDhwLOe8hxbQ0SJTC6uGy7EEzqys6R2sNbCsdegDDuaKk3PIBkBhJlZzXkLLpfwhB
ulhPzmUCzkU08NmNuN2LRh68A36wFfRhv52ov+MY/qNOQEpnK5THDUP9gFMvGzQnY0GwO+g6Wg7R
+ZlTvs0bpVXsBFZdt9v3GakLkJm9W9HhLMSBNpZFJ83HClHXJpbpygk69JeJpT8hpVr6p35Glonq
YcmCQfRRKjLBsD1pupsCXfKCY6P+dCT3wXSqfGfTVvnBchp7NAMSwZ7+tmZCKeopvhr/sDiP8rhP
OTYjav75EWoF7ducF2Te2kB/ChJ6x8s2gNCscWkHIKEmSWoHapd+xG7YED5O/06jtweirUihwSTO
HTy6b5/ZEAD/135KXr62IHn5+ZWQqjE8cJAvvpMRchG+WgfWowBuhIduJGJZLwDu0N81XZtUQd6V
MhPhXuIydloKf9DbsneWGmU6aZ+PoS1fxY5fKy4xi+5BuAMIsCVqQWSzu0nidRbryK0YtKVoLG2Q
ZtHmguyoBM8VExlQUEbUvTTmR6x91JuctfTFssFTbDDti0S+ivmOTSz+vwx/TZVzuV1XJfSMKmdt
pDr7E42GSzGBekTtlFR4dqnGXngAijkSibcUXFkJOdFAzIXNLzrtJRtLQqw6Y3VkXkKIZpr8azPK
9Wy8ED5Iio2sInn08PKLM7GfWbq2Ouja4jVoWv1xm0Jr9lCZxrivTMbcnd0cjA3Ubk348L0VbpBL
ZUkEDm3VSn1hehA/tqAWQ9EkzMRWKPwHUkUnR37/5MiWKrLDRRUEO0eoRDfUA9ToD1Y735LePiR3
Vdr60JkaXZdUayVCQjQ/juA+acxHhr3CxFxaZQe5jATggv/FjldOFq6N76jv43eyTLUAjIuglz/w
ydXaMOVZ/AJ4d2J5iD5G61fJp1iM4WbPi/3SM5I2RwLtaRwtcz8tN+5IMWBqMsuBA/fxp9kzYr/S
r3sXGfXXUjWyoGYNiM3orUpR74K59xOt4QsIQnyAhNqD9MkVogxJVePv6RJLtGLMeYyfcPx04OHg
VIyKDxuQUWblbaAvFlBh6f8YMWxZZzHKJEKDUdYPl7uiOM+5txekHkFFfJdxznBswvrxOEIJIJtY
FMjDe0nYpyyvMv/vciK5JaccjtzB44py/5Qi5Mw5+yAnCDrCqFsHfcBq+bC6cmtJq4F9lzXH/qXl
osTB44ntJNbqnKdfXNuUdlIwBlF7pH5Wa8+klJqpWPgBchRL1jfiW1bto4gN0dXfuIx/vcDQvd0H
zK3JmZhvKDFqdltUIc07pqLsuhzFcGScbVQIL6uniLhVnT1/YryC2ar8zsVn4PNZPTYQ4bNg56hA
jNSQpglxxxcNuE1ty3GX1hrO98pbJ+McsCVWnpD7LyRR1KtJdmEb2begKGR7ukk4jNrAuxSX0p1d
xqsPpiC0EPPclpt96DGCvdop2ZXrLO2wD7a2AwKpWap/dB2FNBh1T2Hq1i8yg7DysllkJ/qKDLzf
DZhgdOn4CS+xK3FEoaILpWTtYGSjtdFDUddYxELAyFBKwDOOctQSN5u14+bu5nsvuKfeY5wX6W51
Ib7r+ierSQux4NdzYZ1GR5m3qt8bSv05A10dXS7cgoVg49o8V7L0q8qI5+UPmO7JPagWr7oVLd0c
lUNE7PcnXwIw4bU8F56+rIkZygCIJLr6q+PX6x7XLD651RDxiWFeV4cIUGCQbNi16Agq91VzydJf
FtP1U0yRSHqwQ10KZibL+vgpmW5VSbXJcbGgoiTAK1ncu1QrZM+7bIQh0KUxRWLAByu6wLki6Lkm
0OMEa5seqgMWX1maZZboDno5gdtvqGno5pw1toPB3KitiL8GWdS4iEnJTeakvVRZw/QbwH80yxJF
rvk6IWNOEW61YSAp/1nRNIkgqY3AqNduJDJgmR7KQ6c6dCIA3OUc1MIfnm5umWZZzjOFT9DX7PGz
3X9nraBmjvnoSaak6jEXdLVGUJijrD2JoGJL8W146AX1u7moVc4zk8vzEqpzOT0KECptiH3uj3et
+XUZQQ/CJk9rIFNUYgd47ArXWHMMtS3Tzb8aV9/HaxK6yrl+oPBWKi0nF8yE9NFF8QRgKxZDgCwu
DbtkWw1XEEf974LNvZtCL6NYVp3H50ru+jTxcJL+iyr4yZFajJspx6RjDPJSL3MepE1tTp6BjQWI
NcY8LfFlGWlPI1tjU2LWNRxM5UyH6XPC08Wcsa/nYt7sM4ao4CsTm5S6q+zHdblfRGXOZTmr2NmG
gvPaZe1MCdahUbQiT+nyxe5FmEeZg4CPQyoVisGB/H/UfIScveUc1M0842Z5M9vpvwADVcWu263Z
Fk63JZUi7J8XQNlHiLVk37yz04To2gWaKKLBREu4+cluGszemYchHdnQLrggpX0boxrQLrhkJ9kY
1UFiJQ/lfWAB8Q8xO2PqtgSsvyVLkAXmwIXM45b2ETwHa1KCUEXViAHXvGdKS/eHPnG2AW0orn4B
ziG83PAo+csvv9Sb5spzg5w0QhZKyPWh+wQNUXhpATv3WTjfx8BXUKyAHVVWDKVr+cv/caEUGu4o
AW5XE2HCSkrZutKQw6/vg9SblYOdvalK17O99KBsvu9dncq+s9RJxbrsWEfUG5GARr/08OKcP6JN
JXydWYM4ylE95Qd/2bjG6YNN/NS4h+uR+7YCxZhola2u5hIKr4GuGiH/9fnzj/R79YUD27sf+q7n
Int+DIcocTd8XMn5o032Zlg6lff6hgQdKkyK/8mjXJyPdRn5Ai/rbEkYvyUmGgjBhzSKTDDWG64y
N57ExfiHaZgcVswclBZLpsgosdR7PXotcckGdT9uk9V4UF4DycSlUn6ReWLLNdtxaD6nY55wxz1t
hgHX0S1kRRDSGm7TmXF80xrJruI65kJYFWRc1RF1jIuld7Npph9gXXnY1/mv9+Rs8LOoBGnxloLU
ZiIo5i+emlApz1EJWk9MF01zWnF9AUdtO4LZL1xxMR1dR6vHZ2nWu0qHJhGKzeBBJnoMnLvzD9+y
6X5LKHzDy2vb/uuIrcTeaIAZv2IxyiERcbcWAeeAfljnioROSHoISGh29Tm6LgfE7frYvppEr1ww
TQh6Ec8CPwaeavgXP0LFy7joOP5ax0ksHshssqYHeLZ8711nyM8IhDYaf97k9E1Kqyj2xeoqENTW
mfX4POV41ARJArWXpiTJ+hw17xywOog/XE5SGpTu9lxPwsHF9jE005xP92dDW+3ieBCSeRgpdCor
Bxve4dHzBnWJJuC9YlJPxu+pvnUPKhpWsMGbCMgjYz4h41amuWNH+QFg7cmPXnWx0L0zyUKss36R
wBva+AWi3PvE544HuDPMvgV3Ew/UhTK1JIUhT3Fy0RhvyI8wtEjc/tw9pDvevbWbmL4n58hiQn1L
r97vfkZ+l12A0SGZMZMNC2Tw/wMH6As7S+dNJ5j5yHqkAKGjRN1Ku5c6cyrGVGzTx3rQKefzhJd2
CYbZjDoNCKs23hsy8bwPfd5KAX5hkRkmOfxvOF7pQyaQKn9F/vNLeoTKItZmV8B6rJ5/oSuWiMGu
e7IHO5PUTdlPPl350GWEMFe6BwEV/PpGOPwE5q/LQXLMgY+FGnM0zSI9HVjQWuj7oqfSnLr/Qp/c
aYvQXFM081dlquh8lswpBvArcjVdSL0uRFSnMZwghAxrKu49XIOI5qCyOJIrrJkOO/g5o1SHeGCw
0oY/bUUfcksfsVmXTRqUKpXkiz2bj1JIIchA80XYPspnhsMHDAGOeLTVzY6OarQt6kPId0yFoRue
TqazL/dtZ3f/p+yovUMTJqvN7zpyFefPBfpc1PqbDNGmE/u4lrHtkWuKod9/o4cm1XdNFswrtIkc
lO3e1Swf4K5wUl6LihxFB15UYNMjHDs4qKfXmgJF0ED+UMJQgrLkevVyrbwpCHHbhCtjGm8PS2os
NR3ryDQ5WNJUE/mc4XbF4SF4A5OIzcgfg6xoIayGacQU+EkbAxvzZB71HBW2j0NM1GZACVTJx9/9
8IMSDBilqhOefOojBX60ufQNBG7u/jy53LNdhkS+ECFEsd9HnkBvG3Nna5h85ex6iJt7a8vqDDKn
OgIKU++qr+iSKAQKc/MkHjJIv7oIzlakk2zakgmqqvHaPGz56n0e+cwaY3ynmdixftFZJcK8P41w
zYrFqWIE5QgOT8JgFZCs+Wq+RwtxFSsGAOs5dicjND7AFvbp66G5cYvE2d+JN3nv4VEwVBZEFVWH
mkjMnBASPNoOpVP7CHS+RuIEjA0hoTFiNKfmaxyEbBlwB8oqzfyppiKMjuBCm0YrUsO7cOdQi1ui
DHXnntZAOyTaNdzvaY+pkIVnAnVAGR4K4pKPgY9P6vO1WSnhsPzie58MgaUp69IQ3E4PWYsiL0AC
b6YZ5nX92MyvfmJj/IIym50B3iZ03MkjZF3mO1ihO3Ge4t9xwbUOZNhgQ4L0gE5/luYCbXH0U6YA
V3IfI0YHxJnwDxmBxZgWJ1XeTFzYruOBtXoCRX9zXFFRG9ifXePLmFKJzq/fOAhW3QZ9hjmR+6ZF
+YAQ4B0C3nMAn4anNulyavLEiYPmu5YP5Xes7YXllwjUU2czCeoKKT1Xv2YW2OJfyHJV0D/uvq85
ohHRZmm0aQU+gIbiC8zYEEOjSc2c9/ztgnWuBCM31nD6diZcuV0Szcdyj1QZ3oYKEBT+kZRTfGoQ
PdRKp4yD3pPL81M1cgK7hFDjMhpJ1MI2HlqRfrpwOo8sSfrJNM5VINbKpmt0GqvuvW5lq7gmW0JY
316MibLGxzFE99KY6VPd5reNy155HEgFRRKyiy40HNgbeBbaJGSvz9Hk/FLQphqRPW82nvtMShBV
yHQR3P/kSHexRUw5xvbNVHmCmTpXg6sachjdCZ5RwURdi8cuzc+e08R05kWHgW1KoFj0mQTSKASB
DsRbT/BRz27W1N17z4uzC82xHn2iKEZ47duZpa5G7CQY2njmUPCdXeUyrUduekuoG6C+Z3wmV1tb
xEHZaRSh9GEAxwU0us7MPeRhFoYy++GMhb7q0Wglk/CBjy+NDoztzjriCozsdkXMyJEbZAQL5Tcz
UBlFuLgip3yBOy19N0nny32LEopyqh28AomyHj17ih2wtWfA4x+D6mxggHShw6kksAKvyX+fCYbk
8KDUZJN/IrtjdzvHNKSGSAyKlTzOtbbJMAguquyjokcyf8+v4sbr1ZawRCAODnZj7CpSzGtLIkkr
JA1cDGdiss3OhSh8A9SX8yeTQ38TT0MlbxXcfok4LC7rHfk+L6emdjr8h0RjemIZ336v9K67zZDV
F6QLTlxeq4tF5rYApsre7gKVMUhTBDHs6lqhsrgXALfeDAD6K9U5VSa4dRfnXjfSqBTavK8NG9CY
JW60Z7xYDG7St593hfEvgqMsv+3MTFFc6KlvaYzkQHPLk/32wPeq4cRUXAmEfs/xzrIlcqa/9xft
TiUY4IuSHuphh52AJ4uhgrpM3MPOkyH06TjcWTCGhEjxuW9yxfrmxhQe6tYyr5CqpVvm7sOZFhHG
plpsK7DWRnv+8+CyhtigR+gbpZt6+WI6ZSVHRADbULmbzC2VJooMJpMbgmB2kQsSJWyexxbyVNxq
uX8YwK7Zx0TrxIvQ6wHHxMj3pM80YuAqqAKlEn2QJeseHg/0sYG04EiPInblvjWQ2bhnE0J5Pis9
zrvKDjozSx8JkvJoJFrKgKQ0vQgGTaRewIteFkhVCinC6st9zZ3PMM8xD+1ZUXYNRMToQTkfaYWj
uE3+lSEynb763oGoYxSAfYa56goq/Kp3O0qY2jHObeeU68T6s/Q5PjOdYEn54VxpUzaKoMFrCPch
gr/6O7EbGSi8a2fbipoo0io8dtrciNe14STUqyITBLQ33dAgmuYF+aoSNnqzSk5H3T29IK54cvuD
b6XQJBNhVzxRh5F2pqTA+MdBBQI8SHaUEV3HjOu8Nm0KSmnYLFtpe8alRcx/uDR2hYNfvvOzc9EQ
1haysJOChfvY+d1n7ospvQMQ3XKPs83ZiL2YUD1DkRn8Q9ap7x2PJXBWqCHvnjfgbtDkeZZsBmdu
rNARo1aAKt2paY70ofIQtarL12nbAFA6qSxIUcNy4k41u3J4Ij6yNENecY4SQla2lQCG/BX5pL+E
4YAQe3owj+svMF+6W3+jm/ltKvOUZBI9fXUQlTw7+oMBLKDf7ezq/G3P2HGsvXs4gKmn8yeRu0ga
p2mJs3puKzzt38QeALJ7x5GywCq4cQQ+Of5ks144Z3qZ7MStNBhWxkUrp+RNeul5zvHT0wPI/Nb+
2IROxNCvEsk7Ae1dq8ao3t4o1TeYJv76en8lqu8VTGwLMsrphelBSwgaGfiXmPWEuTolHx3cvvWk
0G4z2wjYEKInOLBZwRBJlx6jqymiUeyK90K/gznnfn15sZ+ihL4oeisza1SCu5464FLQkiUoxdhH
Cgp+4uSHrBuhBinJCIkFA6y0/9hZL3vOkOoh1rPSO6X3/lZT4pxQvIBc7ITxjpr/rJHgEvYPI7hg
ft/9fH3qk4Jei904atTx+4qoS3Dp/WtAHsg3Dm4Xok7qmsrhCwISWOwAa7ScxDXfIK7sJxgJgqss
bJKB98DYigkU+3zwSfJvIihwgls2VfJU8AMoBHYpPfd/ODoSdFpeM739Ey2e7+aadTK4Un8tZkU4
ba51sEY9xbJcnA+r7RucaX8v59P6bISRnkvFCs2Y9wnkLel/W1qP53y989oM5tR9eC97mq22XTa0
g18QAmeZsNJjc03fQ8jxGLIjD0/LZrLGGOYcXw4yhyubBRgeMvsxIaLnWsF7edHo/Y7vFWrX58dC
FXLhLPEdpF2+eG6qzRXGkHKYbdUw8Mw5v4IQXvaeU3Yl83O6ekw5k2mpUo1N4JwAfmJwywtX0+SN
LVvcr6jqNnDnI/j/3l5JWIypsMIRelvlbX1Y9fzFs74gFo/2d+IRvuzOZlubwBoOKzmS2XtgmyB/
dCkctoXFzwKtKSCzcJrJeAjXiTEN8vy+0yjQrmAK4KdvF0sXgrZDEi/qr+pVvm/sQwsV7+J+QAQa
NPpYd1NjzYYk3PvDRr1cFBvk/H3igXO+4yf6z+jsiqTr7+06+mJ6CgXJcN+ALe7nMpFs9ETcAFFs
KrrCuTOyXlfwrB2v+ROS7jMRqUfW8EvpS2ATMhecSf40/JulwHoX3MB/CGC2OV7gOdGcVQesEyRr
lrqp2nSJBkshCQOm9L4AqvWEeNz8rrxuDyjCKC2c6nGQNH+veKtBMM7/Cibmg3e5ZSfgiIyaW+k/
V1lB9z5nh6nER0MvMWb4VO1fpJhVS/kF3qebRNIVk39AytbljKcuGVmkkrScFwqMAPeu09CXyw7X
XrIkupHbEpBSAVjgl7yeCEttJM9/2R+qqH2VP5E4ziSugXNdaybo0ROdCuBwECsMVzqlVuk41KAv
n79L8JqQ9GNrOnBIMg7ht0XfYHz7k9QFyBwob431XR98ts5OuPeqz8KhhPxaectfzv0IwWv1jZmm
ASB1JHt99pD9Zfv7zN+/V3spSV9VSPcwU7QJ+4dFNgCI3YUhDvN4tfy1P5TazwkWPs+ceOxVDzIp
SnuGIvVuPDwqoTRe67+rnAfNx1tRPegadJDBYi9cw1l1fpzrB397CjTc8eeTZdjA4r5MBMPMIgnF
UnPe5R99fFLMau0AC3iCEjrFESdDWh8LH2w0PjWhmE9XSyp6S2R/cBF9WB9Gg+dA/ClbsVn8TyxC
EhOIBxaPo717GOTZ8X9hBh206FWqo/DjXToMyjmuJHexPGY4T7BXZZ3SKKniUvJ+PlDaDsP/8sxD
txRaF8xpIxwe04o4yTdPORbVjbeYTG9LANfxuJL6i0T2/TNRKfjvoXexVC+aXbU8ewGvqf8GcUlw
dOHXiE1BFmwYyV+55Ozg7Q+6JqIVyy3iBjT+36ykuCK6d5x4R37CQEsMlo/+S7A/57lpYQfvgdRD
ifcyqh5dgZ7aurQhnbj9olkLlSk4ZtUzWItNG7H5zCtn87pNgqgXmIC7pitL+KgIjGHdpfTMRowc
YOCAG74bwlkRw5BWC3w9l8U05wmPlEHKWHuPpAw8MrQwMcJLQYkQs8ebCuSW1utMYO25dsXVb2G8
wjww9xL4PNIVZxpf0R3Krmyk7vA1evDyYm+rsPtXx6n21FH/dXluh8tF4dTmUW8GMAZYu5zLAqCC
QW2TGPQDoYJvM1lV77p3vQBUfTP2prfiWvM59XJHrS+2ILulv0HqtaxWN4LuyMkDg86OKkr17Tsa
0ja4uBh8CNZeZ6FfeQLeWnzogS9kYp0IOwhIppOcxtg1AlMyGBJF6WNVVteiuAcn6tfzLNMJE6/9
nqTrYrSdEs24btSrfyVzs/2EToNP4fz2nY11bSMKBu7caGs/b/maRx2c94PhQYr5bUsbI+o6i8hj
wiYc9PoA4ijzyRnx2APOuvpLpodVnAxnYgGmVcatkp1PiaCdMn/BI7y2xfZ1Im2I7yHPa+uKFZot
Yppb54JqQpdLPWSfAjxEwLGrxSj3P6zsfPQ97ywsbPMq7Ci1VGwZRCuQeWILD6vxNSEwcMa8qe9J
M3BzLpeLn/M7jcd+g3TP5DrR3pr3nsrbnRWy3iwbxMoxW7GHBukDbqUXXZ85i3umpDY75SDQrlF8
9eUI0ZZK+8ujjGBjuuEQc/AQoHy9aSdj8mWzz/XGfrbAoG0XcRE+FOvlO0eOdQdAPX8yWf92/COV
EHuAqg8jrGpz0jhvoq9M5zksnQGjKK4/fScuQvsaU+e9StZ2DANF0SV+dFNfVq8FU/oYrRTK0oxX
t+L+K84EtLpT9ht359/zeyxzkRbZDk1ax/CQQt5qGUTFn8NF6jFVsdc28QAvNaexhhvIKjUwosi/
FIrgJN6lnWEpg5B/ZahL05jnmMIAYGNMe4qczn2Hyr+TK9P8wdVvJA40FGFjNLjCDDbGYLB1aZ2J
PPZuRR4VG4D8jnc5/lUsrmUyrksIzF2/XqoMAnpTORwt8TX5SjAmSQ9AmKKuR5N4CzTcKzo6VDhP
keryh53VglCVJqvfGDSTVXrPD/mKTRrq40CNeh/OKLanUeqfFuOvHxV4fNaCXUSsV72GX/jEllwc
sG+Sfbr12XUGHDQLotBTj3SGcyHiKEJsHQ5vkzodQwr1vfBT3X0ZyLAklH/rAi6D4uAvjBwBERGK
wNhIXf4wElDEJmgwC1p+PCy3vJEtPdXbNDrr9YKmoBflcoHDfasTQNXetIp+d8HXuezM4aswaUXr
orjQFmrDYZcMD5YdoX1pcGHGnQyMkmnpXEiCpmF6X086AMZO0vwGzYPFscY0XmfU/4kLv2JK+ihi
RZGRz6DddIRUXb/T9DDuJQu+n2XrKMz4pE/WRq8JaKdAGzvHqL5gW+F2dgb0ZHM/PxG0Q95ZX1aX
odQ2e/843WgiQiEXZRzvD82SvSGm+GtFuoyuFQTgrlLsm6SBXUEK1KHL4Dv5c0LpnIQdsIkO5ZK0
wWdtnoATX+/rRKamSjTNDH8/h+8epziQKO5RPQCxPkqOS0wNellkrddeDY/7RvBAreAMb1tfX1Wl
c8mYJbty2Kp7pKI0CU2Fpmeu9hPjGvWnmObFiJA7tBtRdeiITEPbnQwWkR94krt9qg+HvkEAIxiN
HaxX8jvQJYDK3OQQwesLnIC3ynGSruiYJaMCfsl94F0mp4QBnlnNOstJB2ds0saiLWzldITuJZnL
ScEguWlfeSD0pCURPN+viNOvIgTI3XEhNcZ4u35P7XmU81BPRvAJmXFgtcXZgisyURB6UIEKks/q
Qy5ZXKsOrjn+ZkP0Dohujs38fA9vPoBKdXnx7PlTmPnvx8uu/rutwe9U0fM2W3qDgjfAMpmspk4o
M6s4UAhQVFTpfg46T/k+OoXjxLAdeg+l3TFZpZK4UAii2qTFC/4ucAC0oCeuakLo7/z4UxCE0tLY
wP+oN6o1UDnhuCgk0BRTkakUEkGjB6AoKcxRtJMZzL3LkjgrKwm7Par09H3V/yz/87lzdYI/3asK
ZJHHPQ7/GDUCKunF+h/+h5oWh2YbaXOxBoUEKFd+C28KtT5/fJ4aoOQJdX0QRgnp9dELC4vHZaWZ
dhN6faXgBYD/yY+Rv8Omk+ZcNCXpN2Us60twOJxYnEZg4yPezdleiALtkkW3EEdJfgz6jlkjW7vx
CgHkei3qAgR0TWVkT8dJOJJyeBYk+GWiS8rCIb/C2kZlhSIJXVPyHv6VntvuryxSQCsXP42hTJVR
PZsZfde6bmg2RDCNpdaG3nduaH6/FZaCd7q1KgxhjrVI8AnTTTOFX9kRh5v3DTJ81BkIUMPWuCSt
L5JE53ywYmRh12z9plF+7gAIf5ylx6mlDsTm2yDCNAl2ijikn8uiGi1bEgICWR9gX1scyLN6RX6D
KoGYHs02xVifu1i3KyKyqfXfP459ZPu0Ej+DA5ctb8Okk4thUhXksFKpIQ/MENd0k+bmjIO2eWCv
zXFSIQtV+MNVN+g3FzdW5hnvBGpuWuUuFwlptLESyymVBb7j1qz3AYo6Zq6rcZeQGz17xKOSCe1w
HZmJj/Zw4ct+tnn/vSAYQZTMSyh7RjbJDvzzYk9mSozqMV88Kdmcfu03+07CLtIAID0r5Q7JGj49
wY7m1wfPyu0XpChhP3/jANZYzzFRHaTD60SI5b2/lK6MtmwuatRvIHyTomaWaiEiMuRiek/sr0tr
m++ccuXohCbZrK0pOCUVJf6v1W7BOcVBgq89kim5zsSqoea74GYrMoo3+hPa8OiQAekWrqXe7ZMD
UMZxHd+GvyMqK1nhhAbc5h0o1uFXnRfXQdYwZ7/N4UrbfRKhPYN5lHrrh8YfzdiPNyKysJSBH0yQ
Gy3C4Yq8cqav0e8NFag+FVt1tbT3kaSltyYN3psqeUyJg/GZF5+k6Qmr6c8utuNca3wcNq0xquDa
urKE6FbLT8KNmLHzI0kVoWdtsg1Vd49+x56NEaf9LCBg26uxf9dDPM2r9jwELdyHiWAov33LSaH+
gqrjzxmuENRQ6IpLZV04FqMs8X3HEJr6mbzvM5Wtqxq4YB7ELgyUHNLDGFCRYkx8Fg8saIuJs3u3
i8txBVCBRksQ4DuPpX0kVkSdRYwlVmGuDFC1+cSqANOEzAsKyAkLp+PvMzDcq+M5XdzdY9QqpsT3
5tKbiwXpA/YMY87A3U4QSD13iMtEoeRwlv/pCi4M7DETQEEuhP9bMMkSEcTC9WoaB9Ml2/t77D9a
0rFrzPLInOpAq+mbHuN8a7BDtLMxFdOIrCcTwqslg2Bdox61s49B93ixSwb/VDsnVvTCfyjs6OUd
4bjoFRTXYz3n7sEruZP8Mlsa4Zx7OIvLTlPxJtLwjfJxsRw7zBD9h8CTuzdRWNEWGgrC06QQgtAE
2ulwG5UpAi2K3ilQCZGcLFADcVG7sCy7kHHBqYoP9+tj45haKfibm+xZFmyXOCOIYcEwOYRWmn06
d/z95oy1EOlNP4GRE8NVKfK2fO1HwxcNknBiZfcNsl+m+5V39+8r7jyhqqlRGewA3wVlyTG8vfsQ
c0mP5jjpnQrxX94UGpEBT4ePS7jn8cO0JDgU3XWUJynJVuZh396+VErVrpqRg0JJk5xYhXSpUzzV
IS3Ol8UfWb43/MHbokrf+w2PJC8rbNIAzaPWr4uMwcMl12CfVp1pdlx5IEOYRXa3HZBTDtBudYOD
UgokkCsd79mqYN3zOSZl/lwNyt/ksKXo0jxg2DbunMZSGXRMX/hyjiiiur8WlVe4owbU7OsFK/Gs
QeMG1h2I+E6FygCAvmln197YxaSjLjC2lsPiKJ9ildt7A+ELWRvGoqw9u0EgVmFHI1cHAY/0s9nM
Od9hqCisF1ANXZ8LtDbnJBmdnxDpfY5qmfy03+00vovnsSA5Ue6gjdd1vFvVRP9K8s4teKwlG5Fn
g/3WDdyAfsjGdP1Pzxo0JI8m4h0CWjg1diHnMg4VIJkv7rvtgvO46qyVi4/6Wpg3i8HSn3htmR0E
YnzZb5TP2MD6V9r2JlxMZnwum95aJXIpiXKP1Uawlof+BukNCQ184K1RW9VpnhNNkp83ycEVtJBy
OXm51Z6qOEkWLAAXnw+DRFHqvqXteu3QzmBgrBBRWjRkquDzlwB/2MZA2y+OXjHd30B7VrCRv7Jx
5KVToeFcBloE38gGDmSLFqM8+nz9CCN70wvqDI8vfuYceH8ZbwmHp4Vr5xyzH6ywV7ADvW/f+czW
n50UTQZJurJARj8acDePxUMv3Aw+lCNC7y1tc/QtUBBZzGSffPnKJSvstQQTX+xc0jTcysRljEEP
BARdKqZUDNepPdBjQjvEGZwB0EHfWjAzHlT4OQiEWwmZoosg0bzo/Y1+mblTikmuhms79Q04XShx
lD3iAxM07bOJUGLOWpqQAqSkG1ceR96Wa23qdfkm3Al09wi8ITR8+rTe8aQz+sYOKMNfJEp+CGGt
X+ISCLsLVPcMvmQ8kY8wOfjIspkfdUJdpEyiGgbl/hxQKtDb6pjsSbVyzD2c4Ig2NDWp9kaNGqt8
RHmu2UjMxwILcPdePmRptHXUMOyZhmNtBbE9x+m5k6Ox6cSFtNXG6PtqZ8VH4RDCXIbZd0FJvbqK
H1ky4pw518Qwa4ESWYrC938Mo5THa/ReA2I4zbCvggsfDQOK2vxvr2mgGY/7jnBd5odTcn63uRXZ
wMzlPfTZgE2sGhGS/SV1EzIIiIrn5ydD0hCTi72MOVRbbw0StYUwoRydbYtLeGQSErSQ1VCW2MFd
HsaD87g8K1de5VJNZq/VGe2+38m5xgyDa1jngC8xS/Aeqvrhhc0BEpVGHbN3R0eDf1s650ruHOH9
Orh+WOpUP2bab9JWbIG3/p3CZWuSftBM/DST+kAZWDd+OBly+3fGkYc7wRbUXMdoUMXPMQeaJr6A
qnLgNdZk1aSdXanRUS/mlWbHFzthAktpfaiXrjM9ndzK4E1zn/ouOGLECdszOAC0VJV6QkMHcDLD
ZKbOm1LinfqMLOn2wHmnPXMgBytps7iFsC9pEnPjgHZIIYL9xx0M0icC/5j34v3cZIidDHvCI8EL
6TwArsvxzTduhLhUjJIjcvzlC3JD0MyAVfVLDZ9VBEGsnj5PxExjTl88TOjksqEeJCQp3AHA3kZ9
iE+T0E2cOYrT0I6xINVa1nA6OohxHwz4lNuPFwUTOT97raMLrP1fXs+gHWPuxTqtUuitF5tsyiiW
6bwovteZ1JkO3ssBfxMjrO7WmHc0eY6CoUURUwSbV0SHKkkIKy42I06RYJhwwbx6V2jX8yXsKDmM
300gPJP/UuOD30T+nH6xcttmlC2VonEEjJ3j8bVovc6k5Kgjza8tDwBdRXpDeHM0UTpf5wvUdk9W
k0nNMBR/QBE4n05AKEW/VYPYpc6AxafCyDMBvzkZheJ3W1M6RMqpTQ9FxAVQZQ4Qeh6Ohw1EVn51
jnem1Qd+D+j+QCAus6BIBJzwntSndMNZGqdaeSjbpQv7EQ6gnRMn0govsbBK7xeBZpq6B8MBdfvH
A3TcSXI2eHPweqepkjP3OVSVNSx0wNMmFmRJL3mKsx6/ywLfQj1qIbwHXvUeQOYCfpM0Nj79BEq/
J1ov4jPAetQ0eAmhH3s0lsuzWT7NNG2vj5ykHzgeeUSq5GyXEZMaiztzZ8hm2QFT3/yidLoxp0E1
9+dHea5P0Gp1RIrmMTX2+2O1SEhhxcThjfcdBRpL6r12ERFnI89ome0iuXE2bNtqiC/jheRpuYzt
2nLm4GHP3syRKe5I1x4/jS+a7tk+Z8587pP8Ux83pvIGpPaL9Azpmum9AB/fQGlC6l+CsnB96iKn
275gAQBJDLkza+nFVhbwickTW8014LoEhPQFJHRgbQjElcvWydGghHbKEaIUSmQZgPHEGw0guqj6
yQ1DukRgui7Ib3TzIlGdveOzCoXucqumPyuuMNfUmQC3evODZRHoLXWa1Rc49snjn7AMkszRguUA
UPBlmH7sxpzlU9yUSyni701f2GKBwKA9i/5ZKW2o7KsFt7kYB4xnJuRVJ4OEvBeiyH93qqH12eof
jQ6fMfaSXB+4UhTCM1zE04yrsQVaMAN6Hw3f9VoNDk4JxPYDmK3Bn0IlvMvdLhBAJSKdzOHu0kf1
C/fZ03AA0Tygrrk9Seq9YN0g3ZRMWsj/8CWeMyZ2QcItbPws9zPYcGBMxnASf8DzSWH7oSNzrSrd
eXcY5Y+SONRBn20bUFPAYzxcQQmPIHkCOj6gbh2qvZar71t8F2tUnId00g6M7cQbC2ZDo79ErCl7
K/9cRNiZSWbiyGTfNyKrc2PtUM0UemNBqESFOK2mSS1gkphBk+tpgcJKPIchf6lrn5RHXRrxkGf+
AlHM+F0yictRPJXfA7jFpf6dJHGEo1yHmJNaptzUGCWz29+0VcNDcAek36MMFVKKumtqstBubGpy
nJTzVXvxZJZ7V6ECyEXKx1HVxfC6DtFy99M3VPVf0nuPNggJDXl3u+UOlYYCalWWN2XCH2y9TqLQ
YCb+e/kWSBz4NVyIKb40goQd7yIq4ihmp/NsdujbULTFRFgdNhu8NWRhfyKzL7Q83jb5DNaogcxy
Y07TXZNK2ohUjia9ReB+/PsK1qDv6wkTHimhSP6yK12scz33rTFXevSz2xkR42yHpgI/6VCh7nYj
brPxyW157lpz8vxzY7NXLKVNI9mF8meNBCV6U+ughIrhstqU48RfZM/KbQYJVU9j4sBWxKE+kRjS
LKZnRJBF6vv1Kl9ksBoWZLLeJmKbw0WvlBJYguvCHEffGNti/PNr9lbwcPb/5rgdrYMJtNxrgdQT
DgLKzV9r/UaJZHR7pO4bf7+WcmvgwRWJXyPWnCplQlKftoRAWOIwVjuMS1KgK0ZBalYcUJqDE0cf
D4YwVL2rWRvXS9TAgyFPyarf+qT8j0z7+iLCq6FQEnJDTqujI0yYGL5FKG9sRDCFbXAfUtMvDkbL
GglD7qOBfonAuHCX41pCEdMwzZ3S29LZdp0SIQkl3ekTw8Y0wSu7Ik4muQY2h+Rud4gbl7Su1XqH
+nBvNoBJVTItx02HnidYSj5Qum38SCTXaMsYLUlSGWzDhCE9zlstKTlF/L4ldD80mSuKwjnl616w
MXoYPNEmksB4aQe9uPLT3NjqLZZCK0HAp6k8xx9ClDmCWWi3NfHPn/s2z7bl28qNE+huRvPy56AH
aut1dVqMWJB0BDPTP55U5VMfl36dkQiLnsxefPo+qaWi0GDwqOSUGIRrrzR93uKKT+QuiPfs1ZAs
ecsy6YAx+FGeO7SI1C/Vpb23gDA7hx4z3FXAo8gj0wG/82NJWNGvusoupJSbwzaOziyBKFrgpMlD
FQS4YvJbyeqtwaMBHMVbNITTprRsUCrr34kR4KpoHWGN20JmJVOhUpx4OBs4BAsEr4gAamhKssKW
7CLoaHDNeOl0fRUi1qiNpNM/xCdkNVtvtAhOza1dqqROFWPlQma3ZOBDQ+VL95b5AboTVW89ptdR
dQ2WKEuD/VxF8AXvtA/pldOVFydOPYKQY6RRqLJLTpxte93ZPQg8ZemTz0NkdOrtcKnfdH55lgtp
BhcR7w/5nB0BaAlUGKh+3zIxsTj8kB0/fw26g2BARJXKAEfhjJjmaWYJWJXZEtRVr1UiAMP6jt2A
9i04VgMODLhBIg5xxzpzhMqAK4MyN4kIV9zOmeytUnTr1CjiIQms6mFI/s23HXzkRo7G3r3t2Trw
vQPeb+KuD9/Egq5lyZXKyu9E+SCK8GaVdS5VAj2UnFfsM5XrnPLmSHcRQM21skeg4sqf8zwQe1bX
S0J02podPi6rNzM0l6uu0ZoVYkSsRhTkgFIdVEDYrlWiPRSz30JtnG9sWV+CHLrAZt50KxoaU8Mk
rGMu20v1ZEfnOq/L/50v777dCqbAMRy4VZnASU6v8jiFe6oUIb8XQmsPMKXR2uuV4vyla7gnQsDN
cQGz780qUoeRlBNzXkUADh5MMX3wNhGYWFmLqXky0EmlyTOAJJmMTNHSbFkvzJJCGk6FzOwd6M4L
ycq5dF0LjuwJW5eWP9l9f3WOrCk6+vJUOAPZFMC67O1J/ncRFohCiKhbdqfpNFq1gMuN8fUeeznP
c9KeX0y8INpbzCMsJt2Xs6Q8mSRyoqReb+XAOcn99g2p2fSmbs/Yav8aDjPSIHyVCHALvNeSzoKm
5RNA0Re/fLmwjo0F2+KGUXSJJ+IClmIpVwZx8Dm0LbJMANCV/65YO4wVGZcebjZXckb2XiBH9Pi+
GetvOjtpwG+N+XmbwaMMrkQB2DSfC6PUCK4x6SG31Nk77Apdza7sdEYqHVFMgmO5uGl3NbxSyUQK
+yIIml3HypHvEqWAmmCeBiRyiFfw7dhuBsfnR+viD5PlEGwuGdjHmMlit/akU8NClF26I2B6IMib
YPMnhR0F7GWv/LORvMYhoy+PRdlJ4F+W51rdnfs8mfKmT/e7+AabZFUYetm5GKRR6UEYspPS9UPe
IeLuVAykoSWyl+yvxIbsC0SX1T7x2DFLWo3b62RsF2Nk2RQeT041VH4bZNH3eVa2VSOBlaTPypXn
AknaQWF8F0Swuwc0VDeW5VD9da5LsRKln5GSVI/iazvJ4QGgMhQXOlhVVVTDjDXVwQChyq/mB9jd
59XG1VIarZoAooV/C95fT5P3YLgWzDHbYXTq3/88xEV+gX8Ww9BuCRgAnfuvtmor6agKAB0H+7Ti
o/OZrKHUcd/YKkekugu5vbfZ9Cg8fDf5PRBSFaIqt+SFC1uFslosezDkWs5sEiRnkzXiHnyMzt2s
GivkZTBc8uKbRO9NUc9i4udq/IelT7zNQZE7hT6EmFGWNyJ2f0Nl2yLrw3R3IcpvnAdYyFXL6U4q
MfwqbZ3jbIhaGBruF2/j2QJZqYqvanBtyPqoMqeC+ZaYC9JX2gm7Ts0YmxVmmegg549CT8Z3A2dT
EAnLQ6K1m1SNpWpDuNbIKM8Pnl0xAiyUpHIPdOh5y6DII1jes1KECzdh1N2bLrtln0L1ZIMtWhpX
2EsxF+sL/8xpbpd39q2NS/sYKO7xWZOYwwZLZEYrN5tL6pOecJf7Zyb+6E7TpKtxTJVzg6L/PIAZ
pviA2ahZNsOJyJrHHqOAkjb+sf+DnwJeUfkAvGzby/xVQArH+GJ67hZpkoTST2d+u1O5JF5lYANB
ASKzprGWX+NplD54v2BJu5fSUWqqfBKiYWGg/vu8wEG0rDavKmbKGMhbbFE0eO9oUNeT6Lsty9YC
yqSwV/3wYeWilHvgU2SpIKbVO8Kx0+fJm7epx481eg35NtK/B6C4BiDus/Wmk/u2ciPJ3XhnSObQ
HcGSO07QSZFNPh9RgbFKdZihu0704PEyWz/tDPcmdPXN+dNkjtWvZoG0xThOeA0s0zA3rbG+DsGP
LVVM2V1/RmeG8YVVbTu1opHfdGkyJpmKlGLR4H9wRo/Ujy+Kb4fU5EOko6UBmUBx/IizcblkVPKN
pB1HSKSs13dQMwrCdxxjRwOHSReQltNphsjrsG8moPK0IsH5mVznLykoeAduoKeKSkQ89jiH56KL
cxH4vBC3x9pSUvRUaJy/YKe7VWWv+RJxR9NrrLTdzuezoWm02PSSOLu30OFYUHDTwVLO9iVX0z+7
o8nlsCw/79UPAGSMu9vBEoEx9GNmXwxlpc/sxrMryPgKTtKm4upeFi36xyXieCDwRKgXBKNMpDmf
TWjKVv5GKMfC7WzLESZ81pIIrSdRhtLy47O36O435OfXyMJbd1nKvNQx1Zdw6kj5biVIbM3OKav+
dI6CPgfhmd7fxcJ9jNwMDES/ngnls5g4+JBl9G6ix7k4XMlnXqrsfRmlq9I0V4ShHAfezOad/nis
DqVM2lhBQLzbgvjw+xYCPCFM00d21pkN/dtMnfKqDxjMikJ3Tj5FikIOwgW7KgNnM8ZSeh9D3JKJ
gorSUG9OeaTPBV6FH8kpz5i+blNXAAHwM7ZYz8hHvpeXFRtubzbvdzc5CSfi5SgpVox4geAeCcgt
sUAekdJTJgwm18TxeeMlhdYplxoTKhyb4fotBGO33NT3rSA4qeSiyjGJHF5OcGRWjNUOtAlwqiZX
EwbSJEFK5Kn06khSgvI5gLYn5YAdRl/j1UfUPbnJzenN3ETyT1LSnIoa1VTtNThr/6NMLDZeLWgA
02VTHGYJftkxpRw33b2PpzVXmnWVsq4JS/aRsLE/oMWcnLu35tShQ1GfmM31/WNAgB9fQ0imfvQ5
Q7ikixtpqErk+0TvnHrRNXXOIWIZzh5PvgHjsQAciohLqBWyH2R3HKC9x9GS589CA+MSAzcMtJXJ
CQM9roVwSoshiTMTPBUVgFEsL4cW1J9nPetnffA66hi2iMkEr+FcfS/I9cJl5lOxH8P4mDkQjzMC
YVoLiZ65A8vgzBQvRn3F5W5Dl9tWSCWizQP8FxGIIHkEmx+hHJMKVFkPe55WreoIsFIcA3zcinjP
oDOEKtEzsY4B6wJ4WMfg9D8oas2XSOxgbYG7rADziKMiDxxZOsY3Z/7lzr+scB6zZN9Bi468ZKcO
qXqzFtYNvaYFqK3ew6jEtMFA3lO3zkW/8CVzumqpNF66jO8/1jEVMXaqIVwuAqJQN0idPokdXXyi
193VccsOCLbxdWMpaHj8fgN/QG7nhQwN7YS6CCk1n/Z/ikfzFzfEW4qhqg62A7InR8Jz4Hvi97kX
NGUH7QtALyUNsHHDATEVj27ty+K3ixllUKXqnXEONuEDzrHVhEmh9XeL9YB9ZIsJ/9fIFGcSdxUN
jt9nm+2pTxJftLLmZYzWiNGFM3U4793sfEXq+HXBpkO8/3s5AhDz/EdUxa9faeOwTq925piI7AyH
IgeFYaDuYca6AYlOk5miBWSvWsygzNpZHk6FbsjjQcA/WYAeAIyF2Pr0Yn9eeFHiN+NLMq37gUI/
+xfn+dRR+IV6qmwWdhqgpX7++fsPk8cs8GUVusYbJi2nX561TsGHpuhFS8qFkQs2Me+UHtdht3NQ
EhmsqM++pDxe4JWWrbV/Y/m88pSDkWoWxTCdaUQqmerXCQgevk9pSILp17eOPg00jNGBjRSXLyRz
0/OWhzDFKQD2I+BskZpbVHTvysUpQiyb6Xqfzftnr8HEnW+6m8HGapCAKuoGZHyYo+NDhkD2MiSZ
IkYQ+28tAR1CR41cUMtmDCXKyJ7R7atseiLpnvwJRJLBTXmryG+/LipKJvR2+v6MecQ/oeYtyOgU
OnWQBSRBgIbOnpp8VVmWl971ko1WYV3MmX3xYZ+zwfMhUwuwepVQW3X3ugjyn64gpjkLGHwakR//
ufZLdy3mtkvsRo2iWIwdg/Jfm5nasQ3siRF9ZTaYky5seWEaaOXQDAXhXQ29ttwcpuuazdBf2B8l
qkb8SAciufmEKIXlTRF1LIb/YBWN9+8zvYW3nV8HpQ/v7qNV9UsCnmht6vHFMI01EKiFG1k3wNuL
tm6uKNIzeSaZI75AU5nRwSlKPG4r8wjZ3GW6EcnqqPej5nAfhtK+f01OHcFgmMOJgLHayHZQ5HI0
Ko5b5aU+pvTX693fQp/VCAVQ4AMfNtEYAkt7YFpTJi/V9z3k0BQ7i1wmU/aBGtfeHWp48CvFioJK
bNOFeyZiHz2DcrtrXsYeNBDXHt5gbW/w8pn1/FPAQs2LPzIcRKgYh1fjwpzRti9qDp8jpaWyUTSB
klYErFNGU9pdffvhoerdNTQifnWren90ayXLy8dT804ay4ifnYm+vsDCAMUsHn6UCE0UIOoAI7sl
wNGBxKSfeT/V6j2jM0I0zg3SbXnzIhN8F+803l6w8R9UQruuVzU/QL/s8ZfBlifVpiX32ZRg/22A
iemVytfMLx8vCvDq1qDv0+LqWeS+W64IH5Wwx+KV2Ip5kcg2rLzCYZIuAO47NB/+ZKHFZ22wC8su
lXj5X9+eKaEYxAGdrnUjFtfK2TCSrQitoaiiWU8lbJfzdv0a3XgLidGCFoCj/Tu8sM8bQqjTACj5
sCJGkBFGb92VzFJtemQQ0LT/Fdnu7SVDF7Z/4yBki9aq8PFFgmGYogD+qIJmbZ398nHtaCFkR4JU
UHhRm5xy74xxjCn6tOiRuKadMdALWIA/Y9SrjD3RlIauNtNnk0iBNrKGrQjequEx+9nKbR4tfZlx
07xEEvkarPrY2kuBh+WZjUWKtF8H55ymFq7lUCusvYmcH9xr2eKs/pr2/p57OxwMgmdtaM2R+IYn
OzbsU7HlQmWLBTrngLWEYTPrWf0SjVy2n2NOVhVgkAdvT5j+tCRPn/bkXBljHhOlgT0CidT99adA
/GgLAdeuRVNHuoHoWnAWCSQpGcTsojCZwCZ0H3ulF5s9lGhI04pENdUMPEnkRvlQDKy+DCBP+WPh
f74Y1ApEj/n55bmzOTS6mUtDnT7pJPboWh0sr6+Tj4ca/eMi1VVM8Vbd0A9bml2urjo1Kl0mEb7E
ugBGygHmfQTn5iimjOy10VNYBFRQr5KbaybjW9kE97g1kKQl8vh+xnRJc+aGA8JS4mL8zQMtNZO2
LqCXkTsUjyPqVkxJTPYMzJfMXoZ0+2rDj9VLZE8nuV1tpP79Q2XE4YCOVQn08SNypMODIO9jcX3P
K3gLA5CiEB2l+nLwyBSZVs+01ASR9XKsOudOQRTJG56sQ03CPqcBaR/eVJzD4QNsp6pG7qMxo5pt
xd3mHkWAQnb+dyidytfmpJOg5uRQ5LdB9rF7iRp1mMFSWUEwzmQxHcMjWVi3D5yF/N0SCRZKcmM7
VlItwulsvlMG7m44ZkWiuTM2SucHXhHcWmttLLYXMPMmJBpv2IZojJYPNrlFV0+djG0grNDYTlY6
qmNTUAcp0Cla3hNax2xXQqxFL9qNLPgSoSCywuj3UbGIxT1op9GasEubWJwkwObhp4z+w6pHIuBi
0jMvVvlcprv+/JvMVKtqd0yYvZN2s9e/ot5PkDNHbJ4uSxCRVbJ5p2tVcXCvyED7mrEQ8JkuSIJ+
6feiJ7rbp2iqLI1MHLMLXKvie7KGicUPVqm0vUcOL7FBdzqshXVpqop3WwesRpa6NlgmdDahYlU1
GSAyzSXPiJSjZPkWfUx7fBuSjcsxX2VRwlU4Qw7ixeiQz2Hf8lqhjbv1FNd99VU6TOwKEd0ICqLh
FrMp/SQ8QntnosdXnJ8rGS/naqtO86aGw3M6dQunEbfYDAleYmdEMtCBoZt/v2BtcJN0POIPziqX
tilM1I2e+UtNHX9qS6dNGcBwMS89mTgLr+GZ6WTDVX06YxG06wRDO/7lV3juL4VVz3Q5AnOluK+J
1jEcx4cenqoWRQTCqUUbXeOxwuICwT8EYSKJ5FsEGY85U3De0x1KjTIijH/VziJwPE6o4XSui3+C
v4m++72Gx/M3+/hy7sclMaOSkjFTv8sbkUZXx6at6K1QaJcQOqJhkWpbVQFFif7cK6jdOlvc/Sbj
Qln4WbWTs/v+Wm2rG/N2/+CK90FF0/374DIZDPdnXFlIRRWRbC0a8/B8x0lHkH0a+fI8Ts+vnXmi
tit95ZXGqcAFQM2Ge/Tx2QgiWwzzSb/iVrVtDYTCJwWl3qK+PYf9LXshtSL/RX1TIZIZqa9/HQIx
lJCtwYW19WZkmpQC/G4wIlFl2FN+TbFrJEXeqr8g6p0WEXBDOQJYH8ZE76gbnljkgLmTXp9/JSR7
pBMYwk9KcUxpxMfwouZtQjegOQu0Ku/qv11MennQ9O0nGtGZuXwUW/z/bx5lUD6c87t2jNFz46VF
b9by3Nog3bx1NFsWj6M+8nuZ+GHqjHUcF0J3+6L97rkqmgj5RgJdPvt/2sXGK46AqYxZeTLF3WQv
t1Jt7JdHzlFNJ4l2EgqBLSjkw1sDrLiH8KXdd9Q5rHRSr/dTy0SMKhmaiSufkqMT2e/RI6vYF/pT
Vm1MxeWRkz2h/lEOOYVWNcLrTZmlG5Z7wg2ysKuTrTv2pz1bOSFuyarS+0B5g0tTnXpnCJbWv9bB
/D9J2WSX3ln1NVURl0sWVK0ncheYppSAUquIBl1QEtcnF2NNEB3BwyJoZeJVgH48yeK9D0hxZuPT
Qjkll3uUaAv4jTkRx6IRkKWdICipRhltLvOLD7McFPUK7fkXk5M4jj5c03FvE2cIHbuTaKMhv1nT
0YemorBtyAU+Ibi99jtDwYwshLGb1wor55w6nBN9993krGp4fHF8sjdhMLguFSgotxw49yQall2g
M2ifV8yttXP/D73wRtGMOGP4ZRkaIQiXfg9jOdqqDgi5s/LeOfObDxoo78FX79n/158k8tEip7G/
DH4hW+HSGozB1KgJVpKfSmEVRk8qEZHjJzns9SQnyymOgDeSqd+G+GkccZ8tTv3+pV55kZ5peJp+
Wp1ri55CecXsbZmIqrWc5lyRzIFncN72jQLSNh5TLkmy0kM9/yvsA+qjqqEE3yEKAB93NqF+whHp
UE5/MT7jk75dt1bMMycE00XEdi45rDJaAfRleaHA7I7F2PP/ytj3p2TS13M6RbR/FZ+b7OVLXoyX
DuHPDyvFkVmOMMRqQOCQFbL/Ot3HMc4R1YgSAWG3fy6K3pkUhXtCyUGORoajm+s46yWHJYjYZ2JU
JPfDZWp1iwyXD7u/E2MYL4elkUJ0C4VRE4UXuQYPu1cPclFn1V6uGBR1I7G8eXBthx26UW19BaCH
Bie90tDmrHSgJoIr9GSNQHnn2wrxFweHeePYh7MyQmi4tBiXv4/KHoXJkKNieuSgdoBjMaRMSwkG
oQAvxXSlsF/0BH/yf5uB7cUz0aXZ6VBaiZ8cin8bsiBfKinkvzCZTMry9oE6rdbYy/LqPVjGfBTs
upe/DOazFm9sIgYhvPH+8MAX6HXsiH/uuih4A7SFnwvWM7medsgccPb5OYGQMmauaSyopoTy4Qe0
AyyXvcoPvWCwm8rJ2ggGP+3n89Sk4cTJK8akQUgQARQzvtrX7eAbr0obpygfYo4S7oNsypfbwZBq
xCo2HASUzE9lQJGmAgbEt3U1kYFTpQo+FY/srHwjop358XkQVpTeg73Z+TqKv9mrtwh0B+qQ5Zmx
/T5DnktebXllNkPT4w5Tpv5TsFBHuznVVhf+F0grO15GJlS8WhFdsuHw1T08jaCYQxWouEvXfFE5
FlECbGK4mEVaTVE5GB3I3/oPXBgc3xP3A/1PCBeEiNebOGfQp3DeEFwyq2BGb6X+o8uYTkq8VVuj
71W/2y30runIsa8eoAUv5JxRTXrK1vyTq0R3IM/+PYiouzJhD6TEFQoo3c5U9PSUpIBvZqvDTfc9
kmvZc1+FPvDg/7PuOPZgC0ITsAcQaZ87lllb/ac1FGoHdxJVUEcWcENOg6zKtqspbDn02Des6QWz
bBhU6dID7B5SULkPiPHk0N4pApgKND5mpLndswE7/Z1ISBhdDewXltJEsWMxaXPOg8q8KvOD1sLN
/CrA99v1sg5qdnBU7LBSqFswd/yFjQjR4m7Daj9z2eX0cZEGtiWpZuOYLt4m1et/MwopYN0ZOUh1
YL0uOn8vw4QhWvN9QrLCdiBmTQAi/6HqtgagMVfcLEZ7x/LJ/dCbz30j9flQNOkwWDEVOONz0dPJ
T0NS60XNcr7d+GIsEAuDAZPbjRwnegxOi8dxQMrqVnT8/IeKpyZolmGZYjE3k4mFOvjYTfvZNBBc
KkqIxaxJEiSxc6Ee5rGRjy/jM2qTz/n0Ucp84JICD4egSP6iS3ARZfDQMeszd4q5TkRKUenYCDx0
jI32cy3FCfPON3wMXP5zeM9Rp3fRdWqw/89VLRPzon5RuNDhOZ3BXq8dtC9A0iuERnTjXzJ4ztZs
dDZ2gMlbiWr+yNXhG4WLDQMruDwuVYCv5tADJ4U/acvOp52VNaAWhVGJqupVJ6+VjRisUGKbj9b6
C23/85B2DAN2qEy96CPYjsDPZYEJp4Mm1pIefrhI+6fFMYEqsSHMwRMIDE7yjlgEevrnp/ZZnVWm
nD8JSOBR1vKwy+pgppLm1V4nKxvhsJYk9zmMRbsMoRkNfFJnK0oNKRnU3CtojeQgPXSjPBOqpQv8
arNnrclsu9X5PE+lqq6BiTXuejLS5EMU18kYx2XaximySMmSf8LTtMEssXClc70TmulRw99LTo4B
RN5YTQw4eQdtDRt3BwoxArDjHVJuaHVabgFL6QYUhA4u6KE/H5wInbwSSZnk9y6RsXr6RY1MFBqW
HzQA9Vr/KtQVdM268a1CCswxulu6j5ZIARqzOAl4eac/8X9mmjgxzWzRKK/SPV4xS488DOR9ZR+3
4WHm2i1JC/gBAZtvAFds4/OqhZO2e6nHT1SwfCRqpDhmbRYRBeJsziflQSy4i1HCdf2TytEP2Kbw
36s9hZ6ZWdxgS6o9yqZGQS2Ee+JzfKLyGa2UYNR6NOINpi8U9kfngWA+nfIrEuBbaeFd8dVrPDhs
RVrNLj4uGMWbjb7CwJody0CXjKisKynWvpa6JKHt3+m4XYEF5U/P11PvHh7i9tahGpfe9wyeTPUe
I4LKdIjs9C7OS7SuqaxYxUO/7pvQGygDL67DO0+XrvIn/PG0jgVlJ81Z3oYR/htVwO4LwpqsdoOj
5bmNU7iTYF/N0jqeUgyOP2MRuEjyChUzIbTltaBsg8WorX9rgw1hhxuE5cEIf9B24kpO2SQIArhV
rR90m94J4XlzQVEb0mzZ2/A+vG4jBOFUUM4lmOWJkdgK4Pom52C3+67QMFvjlMbKOFLt1suqRTVb
IAPGNeQ23Gj5Z5MiIPWQkqfOBaNJo1tEut1aVft4iV3EYlEEfO+JYj7PdA+bKz59KQ0v6eZMdgfO
m1KVmJnGKzM7pwr2iNhSi1pphsEcUHr3axntIDdn4hcAGFUzkA3R8RyL0PfnPXDZPx5I8/SlgQJJ
UlzQcRxQ91yBt21nnVR6XGiTkfOdt3Q8DQHk/EmTbzyszOgnMT6DeMq7gCAwzPvDZIjFwWWII0Vf
GykyXAsXXWZdZ9Kp7zlNs6skb+qM7+vVnmmqD/bQbip7aGifYcAC+5c/q7i/qYWOMYeqo+XoARK7
9uAhh+dN08CbeQKaHDKNKp1vbTCkUwIPoL8byT+qpMk8+lv26Euw/wyMfdEgMNkVBQ1/Bt0MQwWO
TGDQr6Ft3nfloYh4DS9K/yLKuQbM2Tlw6bU6EY6PhqtwEtzjNXiJB6z2TD2mrMjXlu5lAnIj4s0X
jpl5ZYBiqFANEEVwehVDSgCDqLuI6a6Do1tKKjbd+stAy0w1rdg1tzrRv6LplEAPjvxVHiQ2g504
OYmNOtXoXJmr3vhIs1hwbHro6UMx98K6kMmj8Per0fUIfJ19lwN79pHmWYrQkMiIq2EI10t0uIto
moptW6K8NeSAwYxk+7LeCybviVxRchDM2dPVHs3M2kLzgBaxuS2pdp3m6y3p6ewi9qov21dPiM+L
XDoUbteRdfqdDmn+IAG02YxPBvQchV6Brn+H7CM4kXnMaguAK3sfRdtXgTFsx6+RcDJQ7DI2z4SB
DONHpQ3xkv3T4X4+VRJ+IGKiLXiatqcId0WNDlpS3/LoBv07+JWW/PHUxsSRZXc7wCTZ5dJ+PtBU
CEShKi9Q32k8Wob5841FiyK/M1K5ojOydxkpe/A/mVxcSrGBJ4cWJK2/6OmWAcTkD2iAaN70QZlB
9mXHuEQdHcoGWbQpVzrNQSuIUpQwP9qSRdRFPW1N7t36S9GCoHIxO7Qe/QBGxdOi3kekQEK23eBc
SY3aQ5Uq9v7XDZ0mlN4TWS20uLA+FJX4Cxueg32IXKeOfg6Re3lhz4Itb/mHT08vI78RNoKP6/jo
5oYsD6KUKSGCD/IvNZ/PuNZSfGqbN9MZPZSPjq0HfhfXmGQNWIz2ENLQfA6UOopLxK2HEjksDr3e
G4rGUQrTQ11HItLCL2QPslogRPXxMgm9+TzjeMZcMQGJdusEbwliSStmUPvXLCdawq4JmD+ejEmf
tdLBB8aIC4zvtkWSZavAiqsQf83a31o9WXQsPe1Q/+rOqen+AylINq6C6W5c+MWKw2S/tVTzvD6S
TmoXLJW9Ts1BpJCRTK76vW2IpkKynUVYUpnPEem4jq63yof/tK2T/g/hrtY7pdCzxI24ch8w0ZP5
lJj9f9QVTccRtu/lLshNfDgZ8fkNuGhwrlkZaRf8rvcKO1ljztLj+aq2rdg1kHJ6YS+QBXhP9H0B
Pp5T2JbMds9Ipb43y7zKQ6cB/fN9dRrseqIrZisGMnhjlSN+pct9V7L314kWhpeaURD2pIoWAiuq
zGYj6+F2bDertkN7gzZIRgQdRm9lY2WjxH3QYIuFS2OWYTtOBfozg9I0e6/UC3VRUNd7oBhskZ1h
5ZShGzE0MYNHKFnslQyl/yuGI+KyuO7OLGSogUS59s/FYCOSv5nFvySab8NG1o2sVKMwGKq+y5Q+
47TcTvSDy8IWNuGvHqOM8THzC2lqgrbEgEN1sAQbvKJfWpdIvvATdYNy7CrD+qCtVeHulXNeoAsU
GqXwRkiAPGTPg9zw7ezaHvZOp1GdHnDLCRUtXZcc2BF8t54SK6Mm12OtC+ZLROzIMIAj3OGky+eL
6NxthS13xzkXNUduHdchPmVZXlt1B99CqnL9J6dutaSp22+8QlptGsIdKL1gcSsqLoTk0EWGBhvG
5Pk0oKEWOeFdcz1r28CfAVZyxF4J497pJtfHzkfjuK+do4BxJKJxdxBkpWIqf1PTbIPLNcTxMVxJ
KP4v+p97fjDLdu75h36sADY2eRxMeOpilC4QpeGnpADZCHPOv8Zb/3VVRcGhzHqH+oHWpiN3JBIx
FoN1KVHKLwGjKlPeXdxTn6B2ea4TAta1Z6oDMu3FnPW01hI9wfJo+fY2F5+Q/JTuvfEHZd6AtyRy
KXOtbzGd0wajrflRXnya7WyyCM5H4bvxOhMUyn9D99JhQFy+lFv23KF0PA1Csz2KspcVyQgqSQQk
zomYp6njb29ilzXxVYNjOh7lpKZk+B2PLa1QR6DXz9mj07ad/ISgDEbRrY/QzWrRypC8X2UTOOAM
g9vKhnB3G7090UDkqeCbCMWBxp1vrjwDVPqDNH0z2cx0m4aIXh9AzB9RH7A6EJBcPkbphF3K4bsv
4cdLgChlRKND7bXrIufACdyhesTjRU6fMscUTR0zZ2XLrN0hC4FFugpEDpBhs/N7aKWE68mAZ8FE
QWLEjWdtIrL2bjuRtIaiXGJdIxZMqBaa2erbuBnrAy8D4qW+rQEHoGHAmzrCwr92I4QhLs47vN0v
HjkEDNWiuB5rnrNqMsjtHB0YG1c2qxoIZiqm/N11TYsAH2mOCCqz8QGO3W9IpGvfqvu4jKCfE/Ro
CRJj1r7+nKeKuSIMQrPSX3qd4QVwH6dAwUu2y94Ey6R8xlRgfuyWm+m3T2uIPxZTvOU9N4t/h3tD
nDkBLiBHWMyPwgNPWqtzfKDCT4bPyn5pEHtpguq+WbLQTg08P/kWonIe7ArxRcRmM/055haOk/TQ
5sihXflI3ol/GKNXewqCu4IgtECKIssBLXsBf/BIGK4cUxiTPDyO/O2Xg1+/i1b6dDXNwwBcHacX
z7NDGxsHP/IsW6AlYZQA7qPJw5+gVtYk11gmhAh0vuNXLQWjDWVlxs9B1pJDgFnoOA6CSjw+1wjM
woWhNT3Z4fWdos6w6k9e+xwRA1kWSUFUT2h4TAaMVET6NimDz9VfSRIMCzzf5hyKJVM1+KQG2ouO
UCl59THuajYNYu9ZPKzj1cIasDNVB23XMcDu7SfNqVQldYEAUbFMoQBF/2RiCH4YbgJx3RcxM/AU
Lyvrq/sxieBEBLYIMtm1qOzwoh5yZDDTI/hYftSZlJZ9mSFRAO0cVjyI5XsMj9EdBb8aVkoY+PxO
dVHuTd3ju28/P3nKQvO17czVwaQf4l0fYGXH5q5xhMX0Xr6KnvwQLWJc/SVl5UU1JvWYbX9lVBNI
jfhJxprGO5+eIYh+tRGsVelwqVmwaLYhuJ5HvcYQbrgzAuMGj6kIi3RI6VxB/zT4QGh6QHrluNoU
EAHCBbGHjOWhTk4TM76o3NAjRMEHyB3h/71TvIoZEEptR4ZzWMCYJ10X0jVrC7ilN1JQzQWib8hO
GujZepMvHUTkcIkwas8y9RQjFh8nagBqrSD/cdENm5kw2Kza7Zkne8ZhLkQwY4Drx2zsz3AzoFPJ
vsTljc1w2GwlFs0jBPYiALlG0yn1pSdwg/DqpHHs9kXZURJR/xf4yMmtGrbA2UyLnPbxQtAVtDEL
sK8p5MSnIOUtj7mfTzc6Vdhyeow1bCWnRl/dv4QxAIlktDo7taTrJieAUAJuwEUk0BevV3b5XJs7
Py5MjmZOkaxv+CRjz6a+mlNBf/ggSZaht1aw0xOV47RjS5LZrpnTjmfZhuPh7igBOaoOa1gyQZz/
TsN1Wu7AGTDzFUI+aH96gDMBL/eoFuZ1loTbU9YXdkSZQ7oV2vii6+PuhfSn4aralajNDKLibly5
xp4B3zq68sc7EQmL1aTmuuRPgtKWzQO9W8cBQS/f8Tc6D++/u7SgDkjQqDj9+ynAe72zu5n1K+W/
nhgCMw96aLXVZhvY4vYFUEiL+uyx99tsFog/rERwjKC5ByMMnIcQr8C5k/zXFj1Z93a4VvBC18aq
/NUMLrtj+8wYLxHqOq/6XXgSQgThkx53QOmy5jwm8v71NBU7qgT+SNWC6EjNqvnj4PgyNWpRDR2X
t63ekVPoJW3+HHeLv557GOZTZUSHzPzGb/Lsdiah81iT6D+K4xVaafq5d70vPR4klyhg7+gUps2G
Uw3iLAAEbz0s/Pj06nDtwwgyzUDGifVYh2Lco2PBvfJ5v17beKXEf2tBRw6pbQNjKp2lzpLjevNV
8Z0EfkPXDcGpf3XvdScD5/KhsyG71qU9XXDSFJLiPm3GXhQojppJ4rZ0yf118OTCGKOg95owNhom
vfPnI1je8ix5DO3R2K2XbW64QevyfbqxT6Olz9pgTT/jNHfD0zYxeMBWtqo+UKFxmuWgNi8qyAGa
65RjddqlYJCCmQVDIxPbxdEkGgEeIGBc+uv0Az8n8sx9c9rHq7DBsKZKNG3WqiGi66m1XnboBgNN
8K6KrscaqcVBjvxn4avAVzG39VzZsjRkarnPh86NZLiy/115qCLF9pSS9H3xYd+2Vcz/LZ3POFwy
yAVn5wB6sJ9g7I36tJFHFmZ2heQXHibsuCMRxgdOsZaz3QXlelxG7nQBhfbFVEQPkld2AIfGoj+W
4xUQ70ux+z3Jtcgm7W40v0Jl/2mZ9Kc1X8eMyoF1vV4YVH1e/sM0Y89k6XRk+QjRwVe+jz9QcWGx
kliNVT95TswOPndl+OA/cKCb7yBr30QC3SomDrJSpnRGRvg4PFRIQwf4/6Y/kGQnfrf/ZCcEbc20
N1nmrV4vGekTb04BX9gGgZYv7cAo+Cfv+naycnVfsrVJNVZ2S8UYWLcJw/ysp+t6tRLR6372Se4f
CnlNjo4JKFUeRG3Q5G8Cq5AkwxLRW/BY9xr0fkf8XUJNnW7LLGdIPTnfxfHkud1WRIoad365HyGo
yE19AWHyxgBLUHvZPF+2uo/VbZh4ircCNVl2mGSKdlgPLtHcRvS7KBoBMfKmyRyh+dN8+ED01IUU
kpgkd87Aap9qXIrEqmE9NeCYK/oRPRAsZ0PKMAsaY0hZTuAgaKBI3rjPQze72Qp8XrtbwL8s3GsQ
3QkKhwlRTPU8qmN+KSW2rMzu6mG7mDOhpYl7IcsQXDLE6YwG+oaWrfm5Xo9TmJhXPHolYhG66jjE
aRa/vZb3GP0f96MNYzgvrOmgikz9Je2yILNFVHJlJlo/y9hpHHpxT3vUCUWpdLmdghy4SE5psXGc
t99w6+XdsAQ5DcC1rUBNJMPpMVtb8AjjBr1/xtdAvQnccdmzNVSyy3fG8RFm0EDbbZHHte75V4su
2nRbKz5lW1N9xgXShJakSrnxy8GGSgSn2yie5kPGYWXvvn9JBEIU3RhNH3jVRioTE1O4iNAPsxVH
IF46ETq47cgZa9/PCMjhHd8xjbEKyV+9UU1uJ6c5VYo3hemebtEgYcj+iY9EQuzm78Wg6SCgWL+8
Sm/GoHD7dYifcGcqbgAItfumAi89u0EysyjXlKVnLvPWFGtqDpXTiE/ZQiuGYxJSmikTvKE2g8DY
XZQPcESC9mjg7eSzla5IraOc6/MbF9Hfhd4tj62a+RBRdjU6A3MgVkQxeGlY7z//Rj9FKLPS+2fl
QDLLuwJxn2MUEz5EqUFn+vnpw7sYROGk+85HhltXTuIR4ey5xQ5AwlQFgnazux7ax2UE9Q7mapzc
ax1J72J/omL2pG4N2uc0kh+GXHIMzLBJbAoyRT5xFiVwnfZGqn5OEblpQIi0eB5wBeEWbMye/TV0
Fp2x1VuuNnztj8JGXUpWojdLGXmwFTZv4Udtym6nDbj2Tol1L9dmmEQvgk5k+O2fMk0P9DDanhIz
fl01EQvr3WmEa6a3ZD7kUhEY2QSsqSN5Kto7lVVihgWkm7v6WFfjdSEKddcYC4KJm7aBvl7xFDaW
Yi1TYcSxuTeazUxfBVtj8RyL7lqMRvYC7t6EKlnASmpNTwq2tB7D93UbcsYTpg0CePdlGl5gK80i
mc1hQipYnRfXFAJFKj6TXaoC5yjHuJfJvAu6xRlRbOybEloJRI8o8/ylwe9x0CMXe/pFyxkMLtio
p1bWV5qfPSSlwLQvdp7OlVJcMoqurvhrs4BFeQSA7Si1ejHDEcFP5tBO1MDGg02zIODz/91xGkYz
rvQpImf5IKCcCQaq5iGzvZYeyjgBvNZkHClCUTMwj5RY3y4fXBeUxQ1ePaaYvKqY/Jx5YMxsf2bE
LonX8gup7eLaUsVNLpFPLxnfi08/aLifoC4JUBTCxrEivivdoBfCAagnRKmUTkMGFp02tbqTWZzc
FWTO5fmVzHx1JY5aEury6aYM8sK1TAzi8QzjKCRCYCdsLCGHhs3gZbTk5offtEVwt4i6Em+tAn+2
q5lMq001STnL96RJiipALyKSQAGqKHDKlmfSSabqKBum7Y7UjbAYSfzUTy93hsA/X3zpl87tV9AG
uZevgVgW+u01Mij3oIjHWxTKvUdQDc0ZBOsheKPnwG1D3fha21aoT8fF3vm7C1+qjOLb0K2eC92h
HyATkcxIBBl6u9+APgZHtDHjZSL4CHwUy+dkT/Im9Qz6nm+DXj1QRRoEfxY9F+1f7rNGnVWMX2Kz
yfzl/C+rHJJzqrbCjq0WbDheV/CZLQ/YdIZz+OM4lfJDxsrF/LmQZ1Na15WgB56Fsw11LbBYGvBx
a0dhW252HDBnC81vCgL3l5/ORbMILIp/+wFFNCdq2IEaq2hEGC8RpPZoGRLbXf4UWXV5No437tr0
GteS
`protect end_protected
