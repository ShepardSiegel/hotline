`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IQV//2+5pfH9WCAXExDpXIL0NQT7rg5A8IG6JHIFViVB4NA0BerayKuMh6dL5DVnwyOLTxA3O5It
/7AjkZcQAg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Zm+whkx5esy/za7S+8PSLxDtP0QwgdMkcUCPenuTKhzuf0/SoPl8mkesANA7Z9se0AhR7OZDRe6S
jw1CMN1Jups9fzeERrr4SvziR9+pt8k0jFBGhWv3KGYExVr+HMDWuDa9YA0WNWx3xf7RNx1bdj9r
i4mMFUjgTLU2kX8vMtI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WZSFXLWV79DDTQ6z/Y5XAF859Q/MzZGhi20bTcknTDQlQyX5fVjqBSBS1mPr3dt39QpJeSPw9qC6
MbJS3ZO8Gxm3yaHHdLmihEiAGAMHkLRKDyViSFHils02Sm4kw2EeKoX3MQk7uMQsN5KFSypHN9Nz
X//Rrn7VLTgIf/SPwLf+bzn2+Mhs8U/8X71ASSKiLC5aO76OYE31+NRa8xwIFqWQk01mWt6HeLD2
fBAojTWRTkHzA74wLwQ2s1ZR3ia8Xe53XTP2E8uiWm/GochuqQL7+9gC3cMPPzhABUHOyr8av8Mf
hoSYbFNWP45lW/SerYwuAysAvaY9ofv1DVZEYQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
rmPrgCmGgKbCb6IXLSOYy5uvjVTox3bkIQGq7WeJhqh0ybaY+hFc6wE1pksyvcVLLhxlrTI9lyZ/
iiKLnq8UEhMFkau90lwzmKgkY9Xf4EPr1v6YwmLViNbuXM3pFH40FEPMj0m52IKV9opYocif2Ojn
jpI9nYzPYIjw2yPaddI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Xldv6pyBxAX9XAh7r3qBBup2a5MP/PpyHroccDut+y+H1XyrMJ7leMt7RCOLIOz9AofYD92fA5mu
Gu36O+Im4RWNeKRb1hmjDsLszSV1hFeDrJQ7aqivTEpqtVfZv2uTXGTt6zRVH9ey4TTejgzgg8BS
iLTQGHGIh37XoqX4sg2YGWGEE5C4Jn+XtEDEJVTG2NNx06H5PtBvA+fpwVraSe+5UGIcZj51U7DB
WEZsrOb0f5EGvjqZPVqDzHSRqdF24n7TRZjVLr/KWEHPwmnMKkfRbaZqZzLMm+JWRv3GgdputcT4
iVi8UK0Kf3cAMYNTApEaRdrBnmYwNw5YBS9DFg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 42768)
`protect data_block
M2hOAA51rWE9n9nvUXFrQkLaX2qnaeOAdhSPkPlbw5LVL08uI2wCNUmFdUQ2ehadvvokaU1pOKjO
kbRz0su2cHKe0pAeIlm8JUUIB+TDT0Ay2EQv/NatMaNfHoUYBh0FXGnLAgDW1G5PL/P+AFYoxiTF
ewXbHtZV3/vPhTCdbnDzQq47Bs4E8nwFELyDRA3Rw3R1hamrCW3S9dRoaYM+2mMDAg+F4i0cUpML
maIzorODuDF5ZeqevSqCgXWihD30fOqQcVRMfAFtu3tpueSXLyH2EP3lo6pmjUFNcUCUhooo0QSC
3jEo+1Yqz9qo1qcylW6sPCCFRDNhP4krE9FDzvivmQ4i2g5WWww3JNuvUZsaMFFGVGQJW/uE6pHB
ae1VDwZviyUm+bsUeXt8fCkogB5O2GiPu3IADjS72uaslT+dSKhUhOFWHqlm+6lHoV200qAE1IpL
nnDQ3l5ftFrV4efvgq4V+0BKTq7WmvZHRZUzaSkxkjVWbrt1t/nKUNcUwarKX1W6EBD+dcg1MXqF
0rcqo+MbUG1t9bo5NiFkhN/WxkEBnxbXmKHttaSOM4SKp8krZqcMyDhXcy17N4+IGRFLZ7Iz56Pz
GhNUZW6bEVsUaPkl5oNwpFRA9A9b6daMTQ19LJ8Tj0c3u36PRnnb8sHIR866aeabOEAyXtVUJYiZ
VqXS3iDRSr38qVx0JmB+M6+rvnhdIwajndWNvze+NM5LbWzjs4DIsig5hP4QS1K5PKjIQ7Q90Al8
UJBeOAhzeN99utcwVKQrgD5sXh8t2B7UyqiveJ2rVOtJEdu2/rlepMcHPwBccGpQzJ4HeVvcKvov
gzwOmTQCQKy/+RtRthPgt20z++ex+nYWx2DjmhF7ThnYWoCZ1AY8DCOBwFRMjxwgVqD2ylUi+/Qx
eXixoEWemU4YG1eor/zHfRU1YkYMwKIp5OrA9rlyDMwDZI0cgTdUBC+bEShpU0g9++eFKAKFqYaq
fTf9tEYVEMrNTnhbxUfLnLEwaV4nuvW5VJlFm2yG9PBmE5rWyj7gKyVdnewXpjOv14ZznmOQdYq+
Cq/0U6dfPDsXJCJ3mF+v0ar3vQCjMd8I0ZoC82pBk7jWMYBDgQlYvQXZMfRB7e+tkOGTk9y6kVSw
8piWr7qY6gqSE8SeAihns/OgOrIlbx87PtLGEhZvhVVijYjqQfuVbJ+FU7pgWE8fDcZOhMFwvHkP
G/Pv45foVQvQrOPpV83yefM3NM/nzAHUMFn666REciaFY24HgjUxzWL5nOypb4RPHaC6E00mLZD0
FY4TRM6KEJHF2eiSpIMrcxqkx0rhGQxqA0WynTYu32cGnNT855vlffJTVga/GqhKuNyaW37ldVHS
8aViXI92W+iUlQSfyb0Jlc/wZvASpGvKXTaZ9QmsOJjXW1u/aDQ77UkuqeW6GHvJAtdwFhqdNIr1
edYO6AbInWHM9e2LCyqq4iUex5G/Z++SZ2v4A0jzpTfTrA9snKa43hetKVPKg0DzslVsvb1LHGt/
yZn70S4hrZYCWlswOEMYHoVrfKPht2IRrEt4r3JqOisCJN5gEPrmPUcpfvs/nF224zmYliMr9Gv4
kfZODaWR0wF3hz9N2qv9wLadbc6ssq/o380bJkGbMtTXhnf9fGJhQy/wGYD/rrymifc1ZPbox3Ce
NAnLP4YiGEGCOSv0WVE7icduhD6Skd7LL2XcqLyUSH1y+ABQt9hQbx8GMRylKF2uw8dGzFOCTD1Y
yNsIIgjI3kwWAm+4pgnl63g1o7mXnThbaGft7MbnuU/eBOmK7qBX4YJ7jsMjuhKx9rudEgdQgtjO
/iTeW7BISEaBz5VvfcGmzV2bqcfq0klz6P6u+vGKtV7BknXWOzpSSZF9aLq3Tk57MV0kru30udWz
u86FqHYfKh8U/+UqgePEXovHbBemCIe2JeJxuESMtKhjMIqd4k9reOmquvdhNgrWz86Li1NeFyZk
vXym5DeV9+AHI1zo722lNivWEzfVcCraldBi/PynPqr64i4ngpszYTgwf93RgW/Cm0a4bw+r1iYQ
TAgsLfKVMUd0Qqs/vi988MHT/sGp1SNY4CEsFGVQQ5H1l0UPoQs/05VVqT4ZAV6WNsinTN7eDVg6
TFAqbBR2cway+TKJmsG7vaPM9ePU2V5QkEfKsUKpefd9/m+pyClWkduo0gbnzIdfVY9owXR0fgwg
rU7qcU7LUlcnqp9EQQhllzEHWRFf7ndf+hyK1tznWIeFAZ2whIYGG2ld29sE9/6Rco4XJgQONUKQ
/LHYsNzfllypgJ4V7i9PIn1OL9Z5X0FdGgym0GNgDfeaVCNKGwctioTxx9BaKZDGBUiP3/tynSa5
KE6zS7bYTob9tmjowM51YA1nF2Rsn4rjWp1C6KLtcxMVBifBJzsSGwAJNY2pjLgNJGEofe188W2r
nRIGci+OoRxLSPkiCcYFPMbc0Rlp/IPMvUJqyL0SLSQEICMDhd3rgZRtwdd1gnuZHIj2cUvYjKP2
gG3hTjB2g0SVmIQ4tJaEqIclMyG53hJWOZ5aXk1Pywfh6VIWUlRa8HupoQLy9HIpzarnJje+Rajt
5Sn6fO69Sfal4bMnVJeWF8UnZ2mvECwIv2FkEWEr+c/NGqonvIOcoBlp+Nj7q+3RrnMMx21NFGuN
pv6DISYVOumab4WHz1aWgVsNmA8ZNhEbpvLpelATySP/CE4jhUsMv+6njhIawewAtA7qO11rao6R
4074WCqA/CK6J5lCclhIevgeABztfPJDQNBlQmAfef5nuVtRtp+XdjCntDClbQUozxPYMvmcBY4c
O/TLkhVtw49wG4C6DLisAcEZuoqzsDkdUC6QbNExDOXoGlBiZT5qEcr9lnS/n82DZP7GHRkWHIFg
3R4RfiXJzt4x18NIyq54S4/UJ2OqwPK9F5BVfOFM5tqdwP5jZt0lhljxYiEavxfskSIDtcAfDRDy
kI+PjyuA0PXUtmNObprWBQWhmpHeoMDZQmwxl42ckvKHE51mYlYhY8bfgYzBXFnkdyjQNw0qfOeZ
6kQEH2fzxqbmXPFAcCLigx1MEmOP8pEVSgYHPJX5GxNjhihRLp1KMsOi7yZetX/F/b2vusUgilwn
fplpPcGrDuvE8UR7jcHQT1mWf0jQu4x/tXm8aqBqqCH6raDB64jUJYijNrL/ZRsOeYvSgfV6YBpP
ojMvGOnGPwFnDj1Bu5tCIz9eTRLcC3h0HBYJy8UKhITuatmvXOs7utihZAZy17Bf4YND5SEBonA2
oF6Bc/uKyWpNsrNAw9eNpLWSLOJqD9Oh+IUw2AFVmR8TWA87c4hVdyuyVzm0q7UZEJZPmEsQgHAa
zp6yTZBiWKolsF0IHWxbH3tvKooBTwFEh1SAB6F4NuVbAkYQ2sNp7/0FxRlIK5kJVlJE0TSWlkVf
bwbWkqiTk4a53OxXj/0hKhO3UkML/Z6UPgqTEdXkgLRx/6FFuIrIL0BOO1Sm8uKC+aEreUActjPv
FfIRkx1ZdVcQF6OoE9N/WpjizTY+hsvCA/i/5H4qf3ie9S/pksq1aoCp8+q+hmyzwmMzTg/qmNfs
JymAu8UA8qQrz5k5nyngm1vr5oUXqy38v8sZLkp9Zl8NslchgN0RR27ALRMAdZnwzXJVEGWLCobi
8bZuasSmm1TFfRQKANWedduGieKv6hQwCttLcHZ0U/uSYOOrKWMmJ1kvg+yOPFxJT+tDGcRiR6/0
6ZfBw5zQO8eusFhbKR7HmPnUi0J7q4J/YAjUbq6yIuDp1wvZ+K97j2ZDhbE0baoIpG4DDSeEWW4e
+bUyqpnvfYf98NWCYUagqgOOB0/zo0NaVGtnB0wTIN+CuRPTug61FOTVg1dT0/8fgZULHCl3w5Pz
H+wOyQ3jTPcP60Qmx1K7y5FKQQ2N/1WMUMO6X3/t1zccZaUQe+UAFFaxNWLcEf/prGFs+9Mgj3eb
QzFbJcqcK2jC3qJly+m1uuBVW0H6BuQcMwed0MbRmLjkWjP9VSCtay0r9pVlFHTxlDkXAihLP2u4
nbO2Gz4y8/F0QMb6jkKM059VKcsrffIODT8dP3RUKdvYQ30dADBuBlh+OzHtKzrfAgc08u2Z4+sP
zpcRiqP96aC/F+fhfuhmgbJCcF7X0Xch82l3NKSNU6lu8pWZ5PxVIhy1rMZbH7EcJgjgEPl7rha4
QUTlhb4fPyYNuEbVb+xThQGfN4an6wWS6cN8JuCYxlXrovKLnGVi6Wq3CGjpDxCrLdEPmuRQ8pJo
eO3aQ7kTvcotVp7quHUldm5GLm7NXSoaem8lajBC5Jm693JXV9xBkVUDr88/RlJgWOzyiWfEAVTK
FO2F1Lh4Uvv6EC+BeGKfPf1TeIaCveuLaRA2nWLrw+TqFR2fS9IJnCJ7ja2AVEmGZui9vhx5Lj1U
GFCqkmD9gcfpt90sIo6R/rW0FKnQx1dSjBce/yHqH8iKQxjFE9qdiTWXydpihxmfImsulbZKTZRB
ilAnzokqu6qRMEsvH8u10F4EuLtpxsyXPVZEfy6PiBnyTMvGZh443YEcQv+ivjEJhn5PUC8q1cjb
DHu5P89atHNO658k3+JVNXHXKPxPdYmkSfDZJthDFa5Sd6oNSuxvEQTCOn+I3WfvG47WrBLZoV4N
EE5gCcd/kSqKqd4hyFJD5PDa4sufH8xETZg4MgMOvBtl1HlVf/f8Q6IeYC1z/lH9HR3wsWKiYQ7e
6V5CosHHXu33apDOxn5t+qfFOrl3zZbwLKl436XoGpANUDxm1bEEBnB5Hl8k7e1zf0ifW+ESa1EE
ZD2exbYmFGr5j8LDqwB50rnGqtrD7A1Di12nxnqtWa2J3krBATTGfJqkboOhzHpb9sITbdIJDguG
1OL9I8bNmxX3HiJjw8ee5Niv+8w/mqQpvTmFCrDLPBmNjk7b/PgVk8KHzj7KiMpR6FTkR0qyTHpI
6LZidSZ3lGgIgpW+CE1n6tCSAHjAZR68yFDYwkK1hA0/jyqMpc3kY2exZ0PgNtMmmVnuvUQmY7Xr
ItuIvOENkHqnLhCTv0gKIt4p82cpCqLLSWU+PscRLnryUG/gh/DrF2b/gZh/AquOnCOM6mAYXalF
TxGEibX3n0h0l9+94aIli1ggPzcglX1E8x+pfJXq/gPGM7FRxTGa8dOuLw1f1n2KW+OyzkKocExk
qSjca36w8D5J7K5C2DTDc3lOuN02k7tra64lyUIO1GjPGEXsvwryOlcKLRxMOlA+wbBXq0TK5M2x
3fPi6NKpB0KT7wRX7iJDZ1pcMlOEa02J5TJ9binMvCWZGpT8gTn9lRRBbMODFUxvQ5FgNB7z19ZD
Ddqg2UEeaxaZVdMVfIhF2Km2iMuj/dhPregHv02rn98XZny0FOWd+sEmEggve4VAB5QaSQAJq4hs
KC8YD+vdkR3X6AW6HCyYf6gxDnVHL2cKowgANoLs0aGEPwqTjV4DEs9REN5ktzb1RzqXixd6dJ7l
c3AJo+wTzkhPOsIivF79c2uRSpTChYH1cqu+R2zLd0viz6QBjcUWACRGhGdPIOghq0DSItEfOiOZ
o+xg09Lc75I5RP83WxpD4tlqu14tEvghbr663cO5ZC2LJ20dSH1azJN6VCaXKhoW8a5QkFVGhM/Q
EOoKuD8OUFLjS2rdhtkyfFurrOWkLy6JkLUpMu3ObMUDWSkFUj+JVEYRXRQ27W3yKku+14oMqvOM
N9sMyKbt3hMa8jUplj8riPUU20y9lFz96zZzH4vQ/FVP7FOYRyhWWfjAtVC+okzXM0vJMusgqYTn
lA2+DABeou12PggyuQ8IxEpTUtMR4XkdDUIh0ihHwyqX6OP8+9zM6uXmWbtoU7NukagypFumo0lU
GG2lspICtbVv3uoA6KsegbWpPWzuj1PoT+6ZfUeYi3qyjcOoMabC9Baaxw585I/9dAep0lbbE/kJ
4b3YOtt0uzCHba5zfBJzO4Mr6b2zGFXDb/J1v5LUyF9S8ng9yONT1z1HcVHZ235kVf2kQq/0xVDT
lzI5UjLkXFRMxVqj6LYxv7tvPnsdJ0nb0Wj0fiZkBv8nPc5WIUsIJlnt94OPCKJenl6HlpfkR/iK
8i2i9i9pktBNlMKUGkh6wNNOVpA/4gPGGTPOm0n9KJPbOKY9iz4dPIKFMS0xknVKUJUk60Fa4QxS
a70i4VripgZlouz1UiHqRyPHQsSCNYZL0FfMf5ZRXarWJkMMddePy05N3Jw4nTIC8stNxEX1gz0T
C0M+tbyO3r/PUGVplb8Cvporlo7ixpe7evnBI67gnnEAcYymYYksk8YSG9jSPIbSmrO+JnE/vfKf
/ZrjobF3x6vnKor6CsqEw952VZN1/xxN3Jwnk1NHJnxCAAtVULoamqn8s/+LftlWKRfDmGSViiUj
31Nh1VvwZH7TU+QlYfsm+N7SsJ+QUpoyJmdSW86WeLdQSx3+RGRK5ubwz2YQ1smAm+7fkDz0M/1P
TukGj83L9HbozreXQaRctxDTf58MLZzFI4sLLlM7plXnqFwcZX9GiIqvqwPapiYATZ/Fo6SvELA9
06/c7qFrh6457ZI6jU0owmHv5XFbSMzM+aCiW4xqaBr0V/Z5HCpOjOsjw4pJFXGABwGgiDeH8MPe
H44RYnmEiHU703NJsu5yS1tXFMwKcXosR2Wqef3+uGCzBXIOAWjH6Ie444EWnT3PFqXSrmR8dkeU
pQDy8fGK76JcRsXHhDR52zIQpbr7cyLTd3qbXDoMSsJ7yvFXE/5NMPZ+U0YKgHkwgglFdxuia9h6
2v7phs5CC5WMwh8DSUwgeCvExisrLwbb7FN+buptyWBPG7dN6FRRNu1rL5edpC566LqlaDRrzlyR
N7EKsvFSmaQv/YKicGCXJkeXzv5q5njH6qUMJclxpCadBvS5G0dc8b7+KfPk3YBNtpP2oqYX0se+
Ac2PvCSY1dIFTq0nYkIgd8Bmy4Jubvd+EGtFFVhm34qf0z6hrWQI3V2W7oi78ul8emVI9FiV99hi
QNefk61FM2E/KVJ61bsBAIBuu8BXBBYbymdObTdoWlxZuS90Y2s1di5t513P/4WMisrIZGDkvUYS
SBXOb10Cqurlwy4vpOKgW7dWeR9WzUdqna0g7NZMEPv+Ai3XDndpaGlDUXiolCr847Uu9VdHTsIe
9ga+VlbH3xnHlMGXZ0Jvmqm6I714xu2Q4SE4/knPHHiGYHeoOC+Y1iqLgz1Yi0oU8Z9JuB3zlLFh
3aPXjkA4ufdgSgUwZy0uqwXgPexgPe1WXtFQs7GMll+l8jWxPnXgbF0tmr85Ac1FP+GWpkxWcI38
BZpuZS0DvXP1jMN3R39xPxASADYndCk6oxW297Mh/Yom+EZ/D34zF80L6S8UHQcFK1nAH6Cr4MFZ
TkypNSh67+8W5Qd3jDahlLSlLinMg23kr4HSXtIlKvk3fPGojqpjhae1m9yhmdaHKInVMadkKx14
gn919LrjEKrdj4r8t0Cg+lv8497BgMys+wsNpfGzthlSBC0tgaHo9mBCNWHOglWoIn6DS2BL66zs
d2Y8LW638rdEELc8HLAp18HuHp24pC6oBeyp2FfFuIHYEc6yH0aiNoiv7+WQeCENgjBJfyYPrfDA
nFcrPFXg88+npePy5VSEwttgmwOK4p3VgK+5zwKmXYvRO35udX/ImnodPk2Oxmpmxtqn304V3Cq1
GZpE9bqySk4JRy5PTIoF2UZrqUgn2Pr7CcZaAne1VjN8jCkLzEsN3amB53szN0Xx4mTXeNVMqn0F
KzXBdpfpm52pwcnKaWT15q8CI40YWUYN+4Kv78GX8/ZmYfunIyYHKdd3F6KSxiGIctYb6GvkmBW+
Ll44Xbf//Um+dlWcvH9AYBSYtI8z/+seevhJ8UYcQK/ugruBFV/bzmBYW2PuY0fPiQBgoT7d3mwP
YExcKB6mnMLPEZI1y7y0pbicpWVqxBNkUFzfK9AaExeojbu8zFuXdRbtF9YgmsVrMfF2SHLiD5pF
AXuScsTWjvXYZiiT6SPObCJhFCevPDhhDt9lNDS5UHuaRePdf6qRkXDOSkpXhureDUMR4YgdYSuc
jZgdyITFg0LO4r+X0KlBO9q8VLP1H5v5OQdPlYIKmw74cpmLpSV2j9BHij2XgXfvnsbfQOPzyQq0
VXXJ+39zn2u+Pt/mLuttUGAKY41YT64unAe7QuSeq2ZQ6UGcqORsMBeN20QFTPgZyXcKNxiuvABo
livVLAiYIh+3QaRxSg2uqUf6qXzmb0LL+McaDKrTn7xgIvdQW82ft2loT68/HEtU4SKe+NI4Y8QW
Xr02SQyZ14/Q8kH50t7RmEMMmbZ36brupH3qM3INxyjIimw4qk1qTqEsTjGT8nTbWwwst7aOn6BZ
UKYyaKiizcWdZPefYhf475HERizibWOxdr+i98PPRTuEpmXf3XMYVOOlLmnBdGSDDccK8X9dmUNh
wgTtTTiaeszNJa8VfIDLo+CUlOlrsJUIFu3KsVqAoHH60TYZgCvInJS1r5D8PmpP8KnAaXoJ/MSp
Mhedn8eisNvrXjMAlFHgeYcaWSE2QitKZRyW6T3HIL2zgYxIAROgnObw4jufwIDdVyJK7f0IABe8
A16Hi5DzjnkD4M2BcpUOM+Uo3aTU01Yi8ytYQCK178zYKlTHxYidaJQGHMYHT/qh7ykbuWVd/Q8p
HALJmrGmTq7hs/FDyq21t2NdMAJxn0HDMgUWNAOSfBDWecAfUydjIBva68WWou4DSKvApvKmjtF/
7KKHsKuUKvaFS2s+s/OUVMhFIt6FMmUxnTGkvy6Q/7/12CAMKQhDiqxYh6ynVxGdMaCASpjZRuA5
7k/dnf136a/S7whfSZBDAs6QRFpif363vgpUxc0WsYiQhfguPSMzJrsA4e7zpT60cS+zJfl6PrhQ
UQMIHMLwyS/Wy3FhOWgfE4klZPx0IpnoWp+drHoxLpYo2VDRk0OXZIsgFabzql/FBHIKJiacX38a
9//29t6UWms2qbSRgpX81G0V2mwEwmfHaqv9Zh3LZNx89fbs6L0P/Kn14SbfDTrnEtcYCD71Gxif
2zVu6IWozITNbu+z/HMu68R1+Ah3WtmayD4NWZVxotWud+wYk/BRLpv5Xzohus7rLnrogzPZUcao
TYd4bRlr/36TAuLsgwKaBs9Z/M45yCc6rlTMfWhG3jsGYveUB0cO7L1lM0x8bYcBUNl2MAwFoSjk
HYA9X7yEtKrm7zx5Eu5NL6T5OmtIHuZUA5XDNr3u6FvCWE6iqRUU/CPfUthSvKUftmm9pKMq9jIR
KuGg3/694AFz7WvNrm9B7jaElmv2Yv0QoHGoA5znqZKkUbyb1Mz6D2Thw5rwczfxUE4eAkc3RcQl
MCitXKg+24+N6gCyzJOsgv3DoFmfQfuAPMvcF0fM1d5bPaQCfUlyeOoMFM4ZzbsuUYr+/PqVUOoO
70l+3JspJ3hEwSYKGD+R2uZM3gzHcPwx2b3LkfBPTNdxaSw8QxKQv1NykGDRXcfPxzbDzzPyMXfH
lDKIWg1BTa1/zKXNziGT+NIk6ZjAjYALtYgFvt02TG1HFIS2Jrp7IqbulQEOSFOHE2Cna/KjebCJ
i0vIl/bWESJQU0f8Qm1aAF37M2esy2wQLEfbIkmfNxYJg2F6/oK3kmJdLQA1506Jz7jXls1hfVVv
9I15yZgOQs99Tx1IfpScjNE2p3QuKlDYfaOL/Iv7xBKzbAinULW6o/YVsn6QHwKOdgh6Ng06gFs7
eCQu3xdrx7bNU0ISEbntB4VgUeG1Xak8/r3jeSGcsIMGhdZBvYAgZtBvyk4YcRWPuPRGJLsI7+PQ
4VXVajWlhe293u8eoPsSd9G2T6wipjAcBVHgV1ouodUGSGrTDK8uz2VhvcChiytvqVOygTt27Laq
uQvsl6hAZGodnowJwQXJXYF0fypntvQu+TkYHwr9wDvpda+2H2XaLZzA3NFtHXldS1iPhQCKDnnj
HL7S9nj2yMQZDmisrLKQe+HByb5uA1UX3aoDtOFkPhBv+/+tGI2JQS81eDXUa8XmrdBuaFrwF9Lh
lnP8yD803kRaQ09m2YSiJzgv4SNHlM7WDJ8clxbiAX5FCxBGlebBxXhSLZFU4gYVrNMkAQaIB7+1
VHFdqe3FN7O/+Q+lRpORsCM6SDvGmVsP2KeGpLrczMeYHMfBEoiUmAldfbS4GY2LONKHpWtqQBQ+
Kz/Si7L7GaKZG96EZadsA3poWXocKGUEr2nvwQCou9+8m39YrXr5PWlUbMo5Rjlshxx+2TD+c+QB
TTf2ykIXNcVJOm9BFz77accrSTyBGGGF7V5iEakZOI8FDvoWzegSXElEIovxiPSxmQPvKLxUihyE
aKmOp1ea4IUsNMmtk57C3rcVWNLqjMXUTYDqcOqPF0BK7K2PwrW4xwqpgp3ZswZu/1LdfVFK+sXx
QhiwWiffuGHaBht64HEDb/x5XI7UjJrDONKElATv8A/Gcowf3aE6lqtHU27J1XayRB/Gz+XuCZKU
e63zqGdxbH4zJrICi27YntE4NoUP8k/vIfvHFQI1obE5R61geztqeEDf5lQm3YWZjjQ+0mRKeF0e
Snbup+XjDha5vyG9VUj3MJSNe7ZO+D3VyzmUjYeICoSo/sThZCU9kFbHvsU01gqYjbbCefFsQ59c
qxXFUdL2LeFP+2j039uga+GZp8XeDJWE5xbota5sqOEKFT0IGp/QLZ0aExZlsuad6BR3skApYKQu
qZmywVna05m0RdyaX5vzD/1we+t0mgwkNRn8h6Wd5tYw9O0nb8KH4/DkLnsrlVMURccfEyOscvw8
15/FY1tS8LqMta6ABwotTprPpEWw63gc1gMV5deSzRz/kP3XZiFDIlehfjV6P41ullJ1rgU0/WvU
X+Bwk0lpFCt9cDrkPk2jZf0NRYuwdCPYLIUORwZ3+psNjsYdjtYjRXzaom3D5I/bMcSHiorgB63l
9/UbYSh1QQevzVaaNb+z9G0FfOG+fgflTfaj8WG3dsut44MG8xv0VBg0BqTGpznA1ECUaSPF//pV
NE4OIIfteU6PgYjW0vCCXpx/aNrN2PUmPYgbd4iwZdRftVLji/q+0GtMuqxwCps2tavK0LTG0/lH
tPbz4FsHGKYvMxZqmYxVPXhFOJjXR3wkeAW2785INbLt4YPBG3Y9FwWJDZ3U83PgQ/Xq+uztJvGd
lYhf4o4ka75SJFihP/FYIdNLa3eVzgNjMk9pAbpRKekKfkmuAUoBTQX543kAnTZMEOkwE7nN+Qo2
65MNFBM+wN27kEIsifqHDV+O/uNhAWllkqkU+3ApOom8oper1x1c9aC0X1f+6nCIfjnuSvDdqo2k
aZRQO83CMowZkubqr5W/QCi7v3e8HD4P3Hy5q5LET4AlGhDxerNIMsjhoVPgxYCLxLvKoVUJTa8B
pjg2/srL7bnH77jllkK/ncZmJtOnmhoAaCPpSdVYsWjCe79kKV3zKcXz8ValjGABmiVX6QquG2ss
s+jb/d+7CH2iZ4fo7KzanU3j8IgCAKJbjeM63PsOrkZVnwjj9Ros83JF+M89s8bHaR1iE7EnAVPg
txVpi+hjd2q3Rnv0kazzkCAj34nUONK7MLA8VJO9d5svnPs6KMZndN2HP/cAJYPEDPnXx48D2NXl
KkiUDn21+idTtynaGA2jhihltrlsMqRJ878Xa1ThtW1rY//lZUU64sYk4/Zb8VPXdyirySGmLAc8
g87CTAg6fHPkt89c6Hi4ZDALBEm6Bx6ecLtbXKkKgGrQ2CUwDbTczxOLs+ACAHkrPRVEw7EEtQzU
UZ4FJslI/tTXl8noy/48BtAY9ecxGMY5xC+W602cNaBoEuj52fc4JWsnf4enkcBrF/dmLNAzu1wP
1jwL077zA/P41qIS8Bztu7JUFMPi3xg8ce95FdbYV+qLBL48QCSnFxF7wIh9RRHiL2WbZsA+mduQ
/3NfAilqwa4+XeUzXayfCwKsKV7RUvDe5s7WkdAesBY7UyMMuGG6P0MpNCPcQWN8WTZNlrBATr+K
VKbHVzovBCvkP1a8KtUCNltHkNX9EfXFBVkTbnYZrmO4lBtsPEVRHn1uMRD9gpy/Y6FKJ34esA8j
wHaYDr/i5BLd824FDez8EVA1UoYxdBeMnVKlAAIGEWDYu9g3hgp9g55KIzmWkMdJa+RuzOC1tI4S
woRE4WWcLQzzzOm4Sfwxd8NhQ5yZ7nMV+Wf+lNY9b8o46mCtp7rb6y06vRU9Y/bMi9plt/yV1Hse
jCEWrntFg370lR3JiNWufRXrSDw+9YDBdMu+o9flxvVT/wOjh1i42s0EsKCIgKE6GzmbutyrL6Z1
XeoqGkhaIYLvf4G+vBA40xNsqiJhgq6s74E/0E0IaBdkdm1SJD0JafoPQFM8oQ90sW7oJQeKMS1i
e587rVSPZu2g2aLaL/p0WH7J98QRvriug1vkwH4ai/jfIYXwMwRTdtQWJav3CPraElvidfZWe5YE
wXZS51jd4WIzW8g/KXUIiY03Tg4mHbBYYcQDBpoBsE4Mw0TkbiPjiHSoKgCL5U2ehjIlObOUskDR
OETlRZT+GNh+Fe/onCfe/6C2+CDIt/14fYg88I4H1doTWOWZbpq7orFLmt7BI3vCOOJSQRaDSq4M
cgupjx4ijqehhVvRuZyOIv1o94xQskCyCCITqrAb6SJ80pwDyFM1cafXuNO1BaOm8GW6hMQQMrSy
8FbT3mgrWni44LWliaaAYqZeyNltGthQNrO1ubwIKFRiWMopWnrWOJ2Cs9wOxZTwuhGL8omi0AMo
gV7nHl49XmvQ4SuUizI5Ye2uo9ay27RZqmqXoThU7OSfrkfX8YlNDcHwqLPJTxjTZcVhaBq5YQ3w
TzDRIy9e/BesEPJCZKYZhni9ieN43HmiU6L5r9IMCEDfyK40mTXTsuThAzKsCeJFP2UVciM2ge9G
HrjFnuQhxSX73MFYeKt2qR8h2w3idbPeCbjhHhQYnm/XMId4dRAj6ZL2gme9leBWwIkG3G4QrM6x
mgyhdTEIpe7Vm1tNV7TvvG8+Thpx/iXUvcJ1NsrnL36+7eqPhTXoE+Vf9ralK8WfNpB03DIufj5p
HlIXhPIlueiMjp8fH1Uj/9e3kFDHpfYmY7Yi6d8kajiGjDW9WazcG+8GVwwysCF1zOUs6Cm8ajl8
/yFP5FpgVaerLmyGWIBBtSNmViNSb6WdC7mmxMnK4hg+Il8WiDSXW8g2d5BvsO8TYRDrvk1ns64z
jav23xSSdtbPpuwZMPghxqT7n989sgRZeE82lA8M4VExRtRW1GmTzGc+4TKCMA7bXVl4W0HPX1em
8jpv4xaBxI6GqhaR2utNP+qm55lANaa+uWKLJcsvXJCY+/jM89XKvdbUYbrQDnJJX1l0FbtjhH8/
ebxWCYXILbnETVQUibpRlUwkAGMbFkBLrq9rvw/hZWwgY+3h4qRxjJei7Kkx1E5MJNfFIE7lZukH
6HYfiPWwNHIyFI/qKWK4X47FqWhzPfTFML06YSz1vP9dHkrgq1qF0tjR/OUSzmGmlvVjhYtZoqPG
fdlbFxG0HMn3ex0CI0oxZeO5Ebj+jtQfRZOVk4JTSyYC7X2K+EO1xu4jU0tngmvJXdFLPC/7ffzO
P5ymUz3pW1YBLwjBvh3IS4PZ6lpgNZrZJOpsZpcsRg/bvHgAwcFzT9uSp88Gvt8rEOJ/7VKo1EzK
ZAbPSxdC1MoUWsiIGa2h1GkYxUMjVnbOKfFzNeTIJFjqvqJGpP20Y3Y7Ceb0u3SziERZDcyNvavt
/ZuM8ZPB3BC9NraCtUMxDI9QBdHa1uqX434Om+oXQIYFiVsesOxOFIpOMiUYuroqLALp0gBN2CIm
N0m5C7p9TyO1gg6DnfXN/veXHVrb/7yFEvRXzUsGUsRd691npmB6PdqsTGRNPyJlAVHSD9qlbS1T
chGbohii/V6FYv6e1d7+pv5QQoz/2GnaIFLSucImGjHtAWQPOyl0X0Ea+J5JCQNfUgsOwJxFBSmJ
3f40Uvs3nNHHEmIcWfkb6RNPwLviHSUQd7CNpytLao3UJtKEUHeaCH7wHgrSVuRvd4cGlPf88V92
HuD6MhvVqAo9RSG0fUJpSR+3+iinnscZ88qQ/DiphKNKgkujIJ1Ly+0UDnoh/mNSJmMP72DHXK4k
w33dxe4Y+QY1bFA5kAppVWjdaKRH/H7byXqjeNtjeDsO5Kq9hrNGgReh5Zyd/S4w8i1Tct7yx14f
Mm/QDGx0J444u/PwyyZkNW3LozZHn9RJBgGsCEobbGhQdHZT+d7qPlReBflb4Ov8uqUW9UuT43zF
wZb/uMy/SW9G914WsJgnrl1KQB4xTMw4CkIt1mQqz02PJipkZHcx1ViTWtsasQzHRHvbzAS3Lyiw
FbWZcilfiRho3Ha8xZ6HFnYWM6L1SG09OJWjj9q1VVqNK8rrKvEm5SlAzhgqPM7hbfx+OaZKodwo
CBCQRBTBcMBkl8YLB/FOnkHgGhOMdvEfbKO1eHS5cpdmD7kuOMlPd71Rw/UvFO2Tj5Jl0kYvTPc8
B8BDi4HgkGHCl81V/MOmSNTdAsXD1Ab2/UTNRLas4LM2YTUIsQoQI9z8UVTGUGj8uYrguAA/hOJY
WXCRsGHp1H5uT8QIOfeiyGYJ3ONx1yo82f05vWlnwHa8W/Mm66aahZVeAoTFBJoWSoahrioW5k/l
CHA8VMUPOmzMK558c3fxUvJhHa5mA9RW7GHn3Db0oCtUpI6/Gb7YuT5wMhoV6nOEqFYCRzlA8HZt
T4x41SzgEsF3PDQyB36dW1jK5zoq6AGbpKnSTX+wz0LRiErd+WEdZ11wq4q3NtOCgonXLkkklCt8
w6XN60gkX6to1LfpxmuMRUdFuSLONX8m1Oo0hS41JTw81yZ5AoXUrzLhYflLfx3dD76k7tgGVfFu
8YNiKWr8OLZtxFMgPRHaxo3IHIclEacELLsmdX2uuaVwDdsymNkN2RTY8SZzDMpjloJUBEkdA1yz
NWS2pXiViAwl+72KESzA2kmIhSa84YaMdMrxXS2vS2sNRpU3XfWOIrQjZqjdngshC5nBvSB+jYMt
wRaZlThDZ1OFrt2vKLGXI6aAFoUcowlqnDV2/X/zVckU88aVJh/hFJjb//OAEBuJ2QwMva3DKKF0
epB9xlFW0V7fBAP6Mo9w6A6CY3057vxwToOl1BoJFRibbeKLQGdZsPk3QRAO+PmTjI5DQ77tW1jd
2+DobmYJErubNwOM1AAr3LiNPT752nnH1022GxOsB/s+pAIuhaSXiyzRGUPaJwdh/MmL04IlGnQB
xcR3EkHWa+Vt0KzhzxvB7YGEklKetBTf6TK0Du+0nQkVvuHZQ0OrhtHaqIg+vV4HqUslrrLy8Sdd
71UYDTtqL3cAgwoZRgWCmffqd1RpHxd7PbjtIPIqXKm4t6EGtTQiFkRIB4c8gwvgtgQC1F2SDBwv
obOfFzOVXWkVsrrTOpUBB0UMUgzR4w+kNASZ7vC+nt+N8B65fjzw4zD55d/afjHMWwlwyWy5yRoQ
zhBeoKzs1c489P6EaAuLvxhK0C7aXX2NpdiJHfOdJ8g7NDfWotFE0zoNX4y2ujDF22I0l8UA6EHX
ofQq9mK+hIYsugENaNC2st8qfDP4/51htwCk+tZjwOD/zveA+BJSaNb9gGqPy7txihjPrJnsrszq
gycBPVqdUrUQin5cA+c1q/2YAwCTtMTsKa64uKvgbg5j2oW/ow2xYMfiUHqRuS7J8vPHsC959AuM
cBs/A9I44/J0EMx/W7339q0xfELgpGGSBlP5Go6LwS2XPHpgEU8pgtK1e2vBnbgy7/Yz2FR4bEzJ
PjfSnUeTjzBD0mDFAxmJE/2lUagvlbksgbqpif5TnQHJ0VFhcPsSk780VY1AdyG8ECYWZqamL704
QgrQ4VUjyAiXFvuDkm5dwXH9G8w9h27W6OczRm1B1cxELZRCat1iEdJQFbqP4b3O43jTiVVTQG6O
mGeUHbjXwDrINctir+Ble+2uUP7HXhBjP1FPJh0IecKRn/c2e8ShCfDFIyzmYNdS9rVLLt0SFT4p
YTLfjo5JapyWjCOybdZtOLAVUK0WJhHvBA+VKnVqqwWLRY4fhuENqauHZSrvp8Xw5zhkYJjrFUob
de2JIc+ONNdf0ccLqp+ZWyqLXOzQuw8pFWyTHnB2g89ZxDqC1rGsnqYa1e6HhVpYFph3G3VIsS8Q
xQ1ce/kfkLTSCa8OPY4976SZBCZQeVmy6aVcs1zCC3wx/QOi+JlPh0se1L5ovBvcr5TR53FFvIe3
Mz8kUaFB5kxlvtEA99yfleW0f0Pp+70WPrGIYt1Gyii8mrxoHvWxcmQ5rye5ga6VbtzVChrlUhhZ
C6p0AZa3iZVuucjQ5PGn+0vAaYIhZ4+l30BkeqwO150uVhxke4dC3/3julf2b76m0ytHP8FXR8ma
XeyCLrStdECt2W/cCblj/zV23O0gmHW56ADxPGZGofwAt2JY8Hmmc6t6hlvqaW5va31NAYW8dmue
qNWF8pzgQlzEKTbOwxgDKKXyCKV8k8CXWkQfUQ3P2sDJWuk8Mj0zbImr01zWf7N4aHooQVTRGb0b
2N4tWTWHnv2nYm2wPuPEG7EBdpHsM7u05kRLWQdaiUP5ZD04rc8D1washSq5DhT0jbxkwEzfXhoQ
E5kf/1jmU5pirFn+9P4qwsl/CCtIG9TiU0dUD+uJiSf1LZ6AgyTsiPmiXOx7rZtYOi8/CZ+1cqu1
DDvb7g6kITRhA2AJxxp1FtFmAN4MffPoY0R/c+bS0phRKo4xM0sSBIPatcn6ZNUGpA8xe8uSCoz7
6YSKyjEhNxsrc5wpp0/r61ENG0x9PerZL4FypX8KxHnkgbzFzSJEJNNo2pP7b+30yx2SR47e0vYD
ZapwzszDGiaQzjHFCcPFUVfsYQgN3pSLQ3AQ2+KLxsKAIwJs69oJ5ZVTASyq3Ex3ur263hZ9gEyF
hzFkB9KxhS17jO0vBOrdlcdbMDMBbqTdW74LMW0AZE3rueCwmNl5FGEcI5RF7tDZMvGWPpURy/++
wECV0isGwHQA32ZPY0J8alzZHR5cFiUw0CAgJxU5fRb8Y7tOh1nGKxzymet45BZOzJXfS7MrWXYc
CoytM2wpva3TQbKSqssRJT2pPpwsUAaKia8lnAQfpz1gACn0LOCezErjCyg5T5TgQO2kDm05Sc3H
oisblujPvlNREjOrmSiWoop8RN269jAfu8RwBuw7l65HCc68Z56ZLvAOFajWXXZSLn/tNPUfoKGf
P+HQ/asBl27ZwRXecmq7NYv8aK4js4czWk1zJ74buNBm0GptuWEPsc5Gdv1ZGq6wvLoaqO5okQ/I
F36z0yeYxb+ZvmCFtouqYKMIQGkCtmxG0Jb05Xl7bSDXlUDGOQOJYBZ2x3r2Ybj07UMLWDcox5CP
HyIXsfegUBckeWY5Jh5Waz/idgK3EF3vJgs35NJCcbr8KoOjgOLUgEayj+aHGDuEjHcedBsjStVa
oYkgEVZCZvOuEkD2Vkx8BZ64zC2/k1NGko5qpjtvahxZPEh/D2lTZvp9dR/hkZo1RnS4h4xj0mDv
KnXtbT+Vkr6aYzr4QCoXQ5o/gm41md5SkqCV0fbUCB/m4rU5WxoHLisjZlmJMVs/NdxqVFMGNwwg
uXe1F4sC84VXRIG8QhiIcawdu+FRTrqK8Q5KmWHDt5GMmL1kRQorlbdYSc3AsLsZ2NJ3JgCiuQFl
slTgklmvr4WYlU+Rw0ZfYgb2nWSZZMLTWDijVQLFxW+ghOM5E80rUhkM1wID+KZSUaZn0Al9vasR
OKNpBEs4BHFZSq67ASowy26XCKHtnL9GM9CsjUSTatfPOVIaovfQLyRSlxZ0FhjCrIg2G4M1QYol
NAGL3D5s/O66lkmby/XF2iU5CmurtPPQOT5uWQeZtgituW6odeoE/R/R0D78Y0FvxprOHhKZhP3C
vOMH+sQ7mmIQW52EbF8zeIozqhoo24wHpmWbS+eSDmpglsxzm8PbLcB672FiiunZFKOYAX8TYBKX
c4A720NXbWcRk3fS5YNsNh8KnZrs76rGsi+Ayk+VNh1s2bWlulwQMEypJ7XDqzpw5NVOTEfEHclN
P5bTeM87Gul/u3HJt8zdcS7wG6TcIxx88yt3DjAU/CYtYw+oHM63Dx7OEwTYClDWGrwswwqrhCYt
hxT1VmvaL/oLYvj5ZSiBM1IXAuI+pohIhPcyIcaj4Zp+DE3L3ohroTDflY9F7GASTJfvHiHBDbdT
CyUCXTAucBPT90uDcSdw64OxORyQ4y3os7Mw2ttUZb681PPcN89N7phYnJQhnUd29I4k/0Fdh0IR
B+sNp7QUeQnJXSJmft9MDKKGvAKQQb62/1aKIxwimY8qZRzw8J740IEx55T0K8nlg5bYPjrRn8PM
Rmk3kvCdihCs4t8gqRcRxqRL/ul65vz0oliO4gpYC6EEZN8UyZ+8aFXZJudIhITj6FQQ+ly2WSz/
MTptPll+nGIwY+YcNP9y8sG0pmKuGImFsT/8svkvVNwl1BkWuzYLL/Rr4PzKkzy68pVj04MGsTWI
W1hJ8snGbRr70f6+YG8oZ7uCgh7FZq/Vao2zWcKo/5QDOcUXwpYJNeXZBnUhDm2h4+JpS6FW3SVU
RvmWMV7/YGwCw6HaaAYnZF5YoVBWdcnKbhw3ek007rbVSz/4uSsqbkw/TMApDouwWESlWH0rJDJR
bp/X0cc0O+3FqIisTl6RXg7W/xY2SklViSfwBqqqneffTe3gBEC69VRbfwm9w1RXeip9zUdbckz8
0T8PpsB4s7jW/CnaagJAHm6WVmBQOJIAYabQDB/WN+mrT8DJdVeLK61rOjXhkmuA5hlHSsFg/msY
DkXmOX2jaZAfMjXS1lpDnSmW6Bfivn3kJDVJFD7CeVpOXWnvtTVQ1sYVAcrtlKgX2qm/4vrAbHrf
CmyVxBa7EaE+0ofTvzSRwYh4vUR1q/cCaS2S80Oh24GykfJ15MZ+djOyjcoQsPM7L1ogOF5OA6cc
byyKeZIqwwIbe1wKyEgGLyKAR/0lQrcYINZQifl2QnFUnd5CZYp2UwPezf72YupcgNK9YKb6JbD6
T2PRyLCd6YN5fO0Plp1hEbE28GG2kNvdREw+7IKGG1sEl9q7St6n69KWhcMq/f6tDDKJaLuSz0Zu
rok1/MFEYJ8q52NxkMluASYs9VskXw7Ug0qOHh+Rb0Ukj5jow2CapSGO89mQdKnvOlfCtRdlHV+9
eAJX3TmNwq+80CgN1OMNmFclOOtDtCpxW630n90qcnn0hbUSExKZQppxszQAfr+v07c8b3h8bHH8
9bh7sO65g1/1WMfKpYPwcQrw2S5wOD9i5NF4ugkCAvckHtPkCWOgus0LZptlTRnFkPZ9wpCyg4gv
Da8xM/KFs4v7knb2JlefTqx3LpwbqfX6feVfe3hvKTjro603ayDuSG8MxGCcQC3iMJxaNm9G1t54
sSSp4FefOqaY12kasGnYNzTb9cPbpSAAtLittYJgRoamyZV8S0/c6ODSCruLimX7nzjyRoBJ2Rbo
iantSnhT0h9y1RfdeNzaPUlcuMk5/CK9L9MGerUGHLKkvalz51VsOvQymgIHoSl5WCoslccqSmsg
BN3xDHpO2TfX8pql7O078OIwf4KvxOZQJ98S/V1GSnX++UBfMO2h8BHpVkFS7exFt//7cXj8Eb4F
Bi9Yn577Re2oVZEDV8MLs8fzq79fvrBRRgUViWdEaMu1A4r5g6tbw/CBargXpy1iUFQExMc5423S
aHMSoZHH+mqq/YBN1kq5Osgm7aXYFIAx83pVkrdxkJlwBTsYw7jwrMDPt9B7dcmKBjnkkQD4FfOm
KLky+0dw2OTUzA4N1RKeSsUG3kIpPD/caqUAJzdzhQ70qnwaAd76GKhDIWaic6KQVWz+dzmrZ0bJ
L85WAt+4rh+dRumhOO4oTkbpVx6QNjZ8GtCGH2vFbfYJG5u79SAaGNY2PuOohClRBsP/0EU8KeaS
zxtmd/oRPyiYeq2yWOL8Muso0nuEV8Z1/1czdqtf68Tdo2kLlV5QghFBzJdUZR4Qt5IIxxyCM8ib
dgCKAELf/RIKActw4u/I5OUNDOFMLrVXTUD6QpD6FXUttYP2JpZl99ERlLEeaRyiGUCC9VYaBJBW
nmXF4LOV16jrpNR95CFmqQlxzg/ojHOhMPALyWI+vIwACTiG6kmrLFRtMOv+10seq7+cGxhd8+TC
JbaePFUumS+nUwZU/9UyxNrpdI3GBsgnqRhwzG32UxQh8ViYBmoSuXxOe1tD3PLOBfrF/y7UDnzF
dqlawnS2BG0qqdIgWYeBV9suMyC9OosSFLrHJJGEgXxgthPJvVzuvmo1Uq/HoREI++ucwQxDAU61
e/nAaFyVH0lXD/GhztdZRXJyqmiOgi3u10AvCAhtcecWqXXhXrFQZKbwJ8nvTNKMmJCPnQ10YAgR
4HhGqXL5DZE/xsqvgEbOVMZDTfOEjO+hrK9MD+ucSPe/2W63Tih0nF3IMcLW+aM30du01LsiW/ui
5jMCMFbcP2je+TlPg34vWNgt9Dlt5hLoff8H150FULXuJs6diNQVBn08FkoX48sWBJpt7/4cktR3
/y42hyAkNe5XOu54H17o7Qgn/l4yVsS7m1vFemX0+klgpO+dIVXx/9syhjOfCBWYk/kKvaxpJX49
t+tztpBS9WWJ16xcjAQcQEIBuflaUyNd/l5LNcUTT8YmQHROZ6TRsCeduQ7AMA2kCEljmks5GiZB
ZUhPi7wvGuyGLGHAjbFIbNjxo3kpsjkp/utszR7U5wWk4AJ/KsnKm1fRsTnjFwiNB8tOsFLWpthy
FpvFVVerWopGuzF7lqQHAJBJGarUC3HDxTpkeBNewxN2CVZjQengu6E4D1FsNa4doe2K259kXBC5
MXzMOPME8f8UEtEoFYMqlpphnDm+SN41tJyt/h4NlhHpjXn/p90uupi0FGIwMHlfCHTetrzBRJrx
jpWSdABcclZVNYKOr012wYx20/RnWMi+nr/VfWhTiXYg0zl1oagLj2rzv3NpwjNBAxx0uzLHgXab
iJirD+RK4229O3QaBV4qHPZBmpZ8UkH/wE2CM4Ddc+Z2KyJdw9BvWd9ewuMmQv9iQq3E9D4n8fpR
MHExU2aAGRYoI8cpi9sEbLqj5PY65UWdLfbOloZqcwLsIsPlOattmdnA/uVuvizzp3GIUNgZ4fHz
Grtpo8PluEAFb7udvyUgT258FpuALZ8QH6QOBKg5sfWz0ncTQPPBsbV0cW0fXwqmsEqiTzRTaGOm
N9zVu4EFWJQydxGMpToWnXHL79j3eaf4k4yP5voLvPTR1oFcy/waLuRxiveXSXnpSaY+hsiyP+HM
TlhLpbXRpSW/6Cda/okZSzoC4xhlUF/TFdE5NNus+YcSn0feFRpitu3RMpH9EEU5k6yiCo9gHNdR
g1AZJjz+NjFz9l5AIslzjdqAAUjMj7+nAUxXI2NUzxdC2c95HPIZxRyc+A9RPJaudfIznznE/fy+
4cyPsE/BkhAlroEejJhCpK4x4b7Ck2laGkSkAcQnKHz4vS9i9KF1rLXj4+pyy+NFSUxIvL7yoiud
9H1lxf6XCYndyJfeRGvD37HXG/J4CuvOduqT9edKk/lc/vPdYHvb3KPkCrTgWQmALwi8SSuwOeOP
KzTSJZB1UEgDl5DG6v3ro3aQcX1LGrpISYf24Oc+PBlDvON3k04sfMZVv0nUlhOXkQl6yexg+sCx
fAb7+/4sFuiBBz+70/roDRyGvxYu1MCyfe7/s6XJHCwEqa32RpR3FnMsvlJ9elBFa02nv7+nEUxA
DAAL8Bl+p7B5YR/2/IXiyMuEJ112sfCkqT+TdUymffzC8GraUARd64rQQ/KMiUWk+uFWGIQpYZSa
O+T4QTXLvmrfxMKPgwnTJg5tyvsuhty2xOwe8tk2EY27/8sL6nn9XMSqOBXAiPDS75SXGdRlcIAX
HgSTprlmkme3OnohPledkIblvbBGPRZ3imo9honjBPylyIk5dHtRk6trKpIJ/2vCVh0dlFq4KAAG
Kwe9bkG1BawRW0wza8FTwK8cF/9r/+kdQgZw4t+fZyowDu6qiSAU519AG87XeMwbp5bBDmpoZrzh
tToHDHUCaZ4vgURTzRulNIFQNLK2NFvHlwgddpCcIWO4coWYkqtn7m50mYOeKrj/fL4d+9rIPY78
H0u0o2XbLI3lnskl15zIwN1DqQvqQg4Fd2KGaA0pjoHr6ZQboltq38LaKsHT74SqIybU+cz9wcLj
yT1IcpBWf6X7279ZNq7ydPktAvfPY632zN8HzNsV6mSN3DNNd9ULzciH0K+UncTWXupq+HaiPSh8
vRc2oN/OoY6a5kcSzx03i6qk9tMVfdapNs6oFdYIHfAdQO63JkGrponXbWHLfzpHUmg3K2MTY8Xr
xQzWfhoLJDoguMcgtA/m/7jIwGPjlAXi8ciMZK7OJFKS5uGSebOctuglpkcUsaRtP+HLizDibjat
VbVTfa91tAwfkbHVle4z/S9mDUF0jgonRSfAPSYYMriPozhRVGJBNCmsWpVt0aoYLNm8/1+hDDFz
TyzTfRqOVUACdezlLHPfOYzOE5+YSQ3TqqnvW90MB8xS0+gKn2D/1kBinxB/lioPcFWPBmVSTV7w
rMop0QRKFi60moeQu4PmTFrq8wbZbJ3s+R63KJDhU4HuPaTlRMKpwNbhj5kRlRiC0bLqxrU5SpSv
+vZHDx9xQTovTeWtKHPPL42am3Yu6xGE5f6PKhGzxA/81bE28ZL3KfV1R2Yo3sloXWkTQCwLFKgT
iGOnltZXIIjwu0zWhP7AansUuTcWuvnsyApdC47LU87qXKE3eF8kPVKXqDxUrB8OWRaMPzrt7QOj
W3GfhoSLRRn4fQPsJijpcI7ek2tWtIN2zaCtbqdcO4S/LoOuWHTiiBIqE8Fyl2t1baZzaNaYk59C
3+KaydjmmcazXjI1vYU8MW5zpxoe6DGTbC/lkyjDVwp+p13I9Px/tgt+AHLvD/2KVi5KDSOe+/I/
yI5+FnL5Sv+VUXkq4R4WC/kbcjhzF7y+prujWaS7TscB40DY92PrF/gJKf5QK9R8g2tWJHvaO0gJ
4r2J81iYUuCD1F13ZhdpTy8isNb08Rsmu7LjdHzkaR0kAcE5oFCySaWVZ+MEbFT4b2Wo5lcCPx1w
rRJBB+QK3fqMEBU04tT+U2SUON7enrzdNiyI0B+sFLGrrv+U5dJ3T12/Xi8UleBCBXOnQcWPQnsK
vPi6dK8YTX2rt3QaA7MIq2v1u/OqV+/sTlwaKXkvw8moXZh7m8R19scE4KtTwtmf/pklrEiFIdk6
WXBxiYp5CcA97Jre3yaJERQdITSQP7kq8QEiRj9GeYCqzJ/H2HXq8aRPsPh7itdQ90iWuXj1BWbB
Ki59Q4fll67jv1iHPUJAI22eoLqIRfmuA0+Z0DFRfUXNL2F5imB3zG4MvIq5O8NbERMR6BEMDpzP
dcukgYTZlLXeN0l0KJan7mEWaLI9G8QCLQsbP6ZOZh28qXVZLS26sI1QINYnZgEqeSjnfk9rg/oO
7dSCcRlbA3bj5Z2wRhVXhP5JsuLM30s6pQ/OifNTU6C6CW8BCXKl9pEHeBUDxPze6IYvoLtD0F7k
iyLGmPBIKfBCr7BylROvH14CphNt+SCjqX0VAjCxZLjMKsnL7AmmyEU4aAVybn46nZjXJ/0i1gEU
37C10119h9dSpeYcEoaUyPVc1CaIrmLEEqI58+AyaHKZju8QF12nQ3e0B19Z5KP61pnngI4wi3Ol
84kJKbSRXm4meDVSaVc1RQUGnZboJEtiYkBv1VlKELgP/VEXwz/l7utNyZpdTsRI+90VNqUhEoO/
/zpvSz+ATEkLj3qD5y7oozQuaaijnjNzCRuIMVXNFXeDXt/TX37IvuD4x99OCNpGtY11vj0i0zNg
G+j9tfNqfUKYpduY4eZ4SOuDCwJwqfv9XhPicxfRgXXz/JJaVXvd9ic4yNabyUIt5lzOXk3NnIdY
NCQ6mWHSG0Dpl4O/lDwVPz88JnW9YCVJBguHKZnWRR+knGImOib3iU7QhsyLJykFiChmVl/BwZEh
zBOeRzQgHnx3g4qN6ew2aC608vBSPG0heQ2B1pxUaRzJktykoyHWKauOlWFJH+dzGUp63Xh1ANbg
ZZD8FEGRF9uhzUwNBOS7E/XoB7gH9VzBxSs56z7zwmUva+4fgbDSSk5XxmC4Afl4RexwRo8Boy8b
aoamJaXKxHqTbkFyUQ9hjcpDAh5x2RTlSuQR48rwVb3N0Iy/aAuFn+R9FvsvvzsJglqsybzPKbWj
8PoAKUXw95ctNbKzNdkjTEBSgsok1Av3A4w3yZf4bnjFiyAbvbNLewqs6FRrXknN6dpfndF4Oid3
LRk5XsNcDlfBW7A3T22m5bVZwGyDnb1w3UMJdmATJx4PoYnOcVbQUpTy0LtPvjbhac/vAfCoFNl+
SSyY0u6YY15JvX5bbAoaa9kD9HCx+4AWlx5YmQBX7tLB0xGDfFXR7Kk0u11/RBa7CrC1o1jyy7KU
1tZAh1ta/pAnk20DJMe68dCxOVmptGfzmWiTk8U1rsVvl6pS8I2KPqelZGMyIVv85uzbdlN/kU5A
ahcZNJC7mIQg02LsGOGNht+qZdeZJPUkAc5e6+fwyVlADqPlJSi+YiuK+lQ2yGN1nO0uhaIpFOS8
H/+Qk4jFq4mPdfJiyOopZru4dpMx9czE6FBlMEWqfoqOHppWYB34Sf3nQnOjuMSTZqUSUGM4nekX
nxSWaGLp8x1MVXPy/Hw5FVdNPHa11kRwdadrqdOh/uy+ECqwqSWdEbWA/8W9c4g4qJCbYbElUqrJ
+RhlNeXyEXzSmx+rXRpGJXBp877ruca/iNm094YwAPU9oCW+GyjARHB9/5ggSK6prImoVdsl5PXQ
tIX1JOZRg9bcka7CxyySNoevjILWU/0Ottpd3AebNeRyAapHUkI97e+ziN0n7wfb7EYwm8eYHnbz
yBjsGT5cbAhMpcsGuRGu2ElQMoGHQQUjDqryqHrXSRZRHvrNoOgC2tgTSKoMPKnjj4R6oo5bqBUJ
PaSOd5wyNXC5dww09K39g4RbFB+INiftELSvBTE+XOopA3NLRwhhWEi5sqBO8jPuFeUzdMikdwDP
MzWnxU5RDUATZhxxVI4aEIImlB1+JaBLM5kkphgJ3HoHhGZxgNJn3iSBKGGtrZhWYnEQOTBEGyn+
IIecKa/bHgRrWq8JGRPobkhmZ8dKwHqFYhYtokxfkViqcWiBHt1yuWOJNa+V4PnJMD95pVIJhFxZ
EAOH9dduv3DLBxTiZO/tfZUOHTKqIdeKSNL7rUB2HqB4//nqUkrcFvZM4iJi98GY6IM+f6Ql1/y4
E3nppjoU4hK+KxpKbDXex+7vT22STsvwy5FP5Ug4WwmbuOptf+oSQCbyMjFDD1gZ5lmaMy2V5LA8
vj+OZyCQUz9R5GUc4pcimFH9fkoyvy6QfHBX9OenXuxYZlt2ktSVQ8Hr6367hsH+eaPwCExvBWxU
DMPZhuZiuqtcr4/iJLIJdABfZAwyw2TSLtAaReRp78Y4HBMBi6SvrZeN82sv74sraOcXZmpRbWV8
ub0AcCGcFODG3aUaM88r1RuPdRRsrhihc8VVk72bxBXJgVmTlsZ9ZtPpkmoP4IOzKpAScjK2cKVX
mfozt4ymDFLAROAZUPsA/kpxGRfsN9E9zKxY5iy/EYajOjnUn0BZIjh2pd6MdALQxICCWRJxXZN5
lKnNuplig3hrspVsT5s9p/RH9BppxIvtRHGw8ttOP/IvU2yXAOqRPYEc04svclcTt0+TgUGy0U0S
jE9R/NGVtLxjHHPC33Ue8eT0uMfGZtsRiNu3n9N/DYFVuB9TH/ujimPyQsnzOWpitDpe9XVHGql6
9QyEARKZSGJeqqJRGB5lMiI1YXOgn5SS0oIR3sGMjw/vPSvavkRjxcmK0rkB2KC0edKkke4SFAYw
grNScWiD+zMGwxEnv/nkEVpYKJ4KAaZ8gc/2HWe4mLi1ItaYPsae4YUFRT9FevtlVagf7uFTHmu+
vatQZCujT0grboFqEtcV26bSHmBlOOjLm/b8qEwPSkfvvpXHcZWh9aB43PFBdqF6gz/jQuglNX8d
vxguEr8LXaGK5+IGMHOyg3vkJtDAvRmRrEsXC9BJhIXl9hQ+DiI14cAoYbBk0G0nuNTnxbwDrn0r
Pq51DDlXoFADoWgR25ADeHGF6mz0ewzw3BSh1G6/0XqGO5P0DckIg6CxyYOLCjqn81fy1z35IMGc
iPxwxR7iBwroaCCB6gHScQJ7GGBUNJHtvlzobDBJx8MQi5tLFrGjDSOtK1z2Gu1TDLlP9i6ChWal
7sNU0FTMZU40IttStn48q0LqMrmoTf8Xcu3c5D+vQaiUWTJvrE2/qEsWO8om1lCdcD7r7QeLCgdS
vUQBDMIptYPWT4hCj/iNXpMddlZt4lZFmy9It7sxKR+9crtYLKz50kgi28KE5WA09EEPlki0TOXB
ntgxKyAS4WDzU/VsptPqI34IYSfRTSLFAhuAF5ky7q4scuAoQ0Ui1OPDhD2PGLN6dzFgqG97MIt/
WKVFrqrdPnSXUab2cppPw11n/BGrXNSR+yIfryYCuItKwzV6bRZS8DghyS2Za2/FVnOk2F4X2qkd
+hSZAm7DH80tMTtl79UMmXI9POGmENIVY+OzRvdBHjz0DXOUdgzud3fKCSsKjlyEzE2Nwgd90bPZ
6aa1ZBY3qMpcdSffPlMTrqpcSnHBgYLXqevRR+eZ9JFruTLHXoBGX/8i3IFRpzXcCFBWjJAPof5r
vRdeGW6S/wSyUs8Pzs/31rMkMQCIoCInifcSJA1AS80D2jsgHj4etv6Q8cajP2bQEB5Q0XCZcLzA
wwMB9Z/HMLWQ4t1eDxSfUSQPqiXCcjWDmYrjyOro6+25kyUc+9ncBwh4SzjCWtvp7rKp7eNr/b1d
zwZbFL97x87QAOIiJREXAQOgnftfWH/qZmCy5Se0SBNJreh+dPA1dA/H8dL/SzowWh+WtH0iUoZu
QGqTEa+3CFRjO0Q1dXF5tX2/lYEDa8zuHMsphsTTex8nee6wxDrpM62JjAmEd6dsmGOVGvez55Vp
Ak75G4r+gOwuSG0/o88v8Vkqkcfzi/6tS6YRzu8Z8D4ObpWKdC6GukgAPYzqyyspcHHtT27zGB5B
t3PNq7AP2wp4QtEgBKS9o+X0r6RVtOIxA8Vohkb67p5H/AXUriqT5WDOjAvG5dzBopXNpWi38U68
fcI6DgixzIAa6wOfJO7vGxyu7Ap4vh9K1PChD6P9JDW0nK/DFmVFW6wWDvYJbwqcFiooOh+TK/lX
+rDh5BEok19TaaQR3EdQo5AGLmE6MOXjynN/Gk3+COpGWWpYPa2UupSNtA9XVllM9z83ST/MICJK
r1zHWqnbyN9EUyhLqGo2/FxiXCvpGxzAat6mgMZ4VDDzCoz3+wddzOFEtcXMBe9JnClxRBYBK96k
nRHM5hs1346JRB7HnFVBv2Ite+Y1oRZB7EXTJxtpbg97nzQme2v97SOLlGJAK8tsAFqcXVaTu2Cd
c+Vt4ftjxK6/3UXw7xt4JBkU8qT71Zk8cYG62EkZBVCmZUF3H842XlH925/wV2NHu0NCS+f4snQw
9ceMQsT3o9zcUqAbWChJ6e2GHyTvKO1Gj1jBDV8Gt1mhfQM0In7fROYeb75ZJTPuxDo/2xYcDjHx
cUai0ylmVd0fOwW3zbM3QqJ8q1rPpyGIVZ7zqhUMox3V4ZwVJR/pt24ZrmeIzQCrNtfDYrV4Qg/G
uO7EaGYDaOlzHUm4BhRM4FUR92DsRc5LXRIrGEhcxNemX5Z2DIZi2cyp8nkD7C8nzbRsjWtwqB8I
8YdPQAhQsyTzFXmJ2NsIjUCDVLjxsWCHEBERnVmtgNFwYXxBMgbSsJda45buaB8Z97pOifqCnmT7
Y/EmSMXSAnfZCK8wTetRCTHISk+5+Srx196CtdGN0Wef55e87Ga4f8Uqy2+/svhHMx3zfwQ82f12
rUgS+YtC+6JkGE8tMa/fbElJkATjWBruQW8O8+WLC2EzfIzAYNKfJfsqwVevP3iG/TjY+psL0e2i
4DMOHknwCNju5uQ5TjcI8bhcgemm7e5AHJNiZcJI+Ti2CuOs6qEJEGy7Hf7h7B9lNDTe1PMxbSm4
n+t/XOa4S/+Yx0x3l/cwxQE2+qM7IjsyKlm+iHV6XqD4g0VjXb8X1tZQ6BsG6sh+Tv1vr0vK4SgJ
9+EwWbiwBIKrAtWb5hg0oa3ugG+fVSgPTqtgXd01tFdUBTKzYzmo1fUJSYLQmn2mPSbb9MlhAX1i
u8Oa0SxgNoZCxyc2XWihOq4I1+JxQWClFpg48fIYdEQdT0rsAHtI0R0K9mD7/4HHpcnLlUzcYqKt
t4NwKxJFyFAwAgyk88PCYjpkgiP6V2dGoIpXvrkHy3rTNCy8Via9tiAnKiCbWjX2cAhg5EDj7X9R
qCxls0G23EvQrUi15hSvHBA5+gGpve/FbnWeJ2G9X2Rax4x0a+NFnaltAeOpu3/XcbldKiRE/O32
6fRA1Qmn8EPEdJfX9olcwwktPpNCsdyeFA2vSh5wM+j06zIIby+BiFEVFqj3IfeY8h67UlLRPcuv
YLuQgTdtwt1F5D0WtL2E8SJJOZLWN3+AigNC/FTI8/w4sMnT2/qEgYGzj39z2Ca586sTEIyaBEw/
lHmk0oZ8OevtGWdQnr7xu4yRqgwhlDZgIzQ9P+r25THt/+I9AsIneiZIy4LuSy6HM1YawDCjhwrI
RBavtrruGhJZ42u9dbyevBlJzj0wMd4puLfSM1vJJYR9zdpBv8Ke4jpfQkzOOg/F2QnOZ/gQf5dm
j5IpLMiREVllIajnTJWfFhbk0BesfvSzBSDhM0zns0zRs29BTO+TPlnz6zy0HHs6rTKRKZzK9NVe
y1t9RuMJ36r0W5OaiiDA60nUa5wNdiuqIH4+Cecuv50TftGZ/coz8gmEkpOOjGu3mtRIf+ortUDa
YHrbaY0Fms2Ep3anLdeGR5oLd4mLm4RBvUc/JrQdn70tmvgDXVyeWOFbWSlueGW/n8PcA/gljF6O
PO+Q2SZRmEl2EURPPj0FiL1MAGo9x3D7YDTFy9y2uzyu9Kho0YvRprSonlTvKB+zcAXFRjpnRzK4
ILw1OOpPl3SN0rwObATMONC2+S7S/O+oH5cdTy/tdMDTbPhFMUwYmFq7KE/9rFTISGRK8cCtZojj
N2a/Kt6KKdvLfudTW3ISeSxBWF2bDtWBXtMr7fcHmSLSJ+sFqqBQNnyp1YYUmoH6mHL2q2ILloHJ
D3QOvXmaLhlqN8ZC5tbRNv3QAwpRF4Y89p9D3vSQyM3oU8lkSaSNiPYstqr5aHjwyqwCkJMJmhi4
jL5C4iiIP+O0C8h7isonADCVidbEf6iALH0D7Mdd44nvBu+eAC2GtWa8hnMj7iuqs2a2B1jPw7st
oK/ec+vVh+vWpasAVUyGUcvWb0y03aBWdYnEWwSo5hDY1WddxerVpk8vb9JJPz9sOmVCUEOzcQLY
DFm2nSzqw84gMRw0fRiG1YRnpahKPe9kUCa1V8DscnxLZT0RYwbI4NgeCpyPkvlrztQild4LjWSB
wNUkhOABUDFfu0a/QJbLNrxjxe2vodsNLSlYGPFzUhvVR2qs5EGDoss5+qbZqQqhTsYVFKdDiazp
ikWztB/62WQ2GAUriOxNRNU9GnS8YoB3i1Gw5F934BI2AWJkvroCS5kE8Ya7218gGezqbCYGUszV
JSV9jNVeEjXVWrSXypnvLTPdrt3UWouUNlpUzqA6SD/JxLj28NwfVY2u6BDOSQnyoq3f6KIc8lCI
OfH75QTiAUYyBi8ePcs7kNIQ2QICPCwfy9G6+VCP6ex2PgIPrD7STvYEXWaCAoW5t53H3Qm2lK0k
aVsbpyDMGL5f1OrzuO5vz9XgPAuGAaOqlSmY4jA5odMJ7UDS9XckKpmRnLF7gQxMKpRB5n2q2wCx
TcgKrO5RJZUbnmYHesz4TjjiCt9FNAV1//vwcXTDTwiQQNmFHSDc9Esy4RGneZyQUKmFgzQE4TEs
PRmt0QxiUThffa24U0wanwwbJtBP9sEQ5+FvePBaUyt2T13ZFuLQUHHFFwX/RnhcnBPvh9QzfsVL
gZYejWrUdBcvzh0u7rb8BY6W7I+vae8VCcEYkxn70U/zo+Lz4vhQwnmvB/fhPfQ/DtusGL/Ts6Oi
ldUyxLm7sfwxEuUrNWg9ETvAsJN9Hmv2DJ/lx3rDFTcJxOnsdOf8TSpaaJsnD15a9ynx+3rfcH5g
kgGPkgIiCwdbXS3NdvCdFvR5RS+BiZwOKEE5KA+svIPyJ8VnTv9H4ZjqTNbwTX+1sgbFSmN78sYC
C6CcMzIm+Ca+X1pkCUvx7xQz9A94OjcLDyboNER/ZKrWjf5Eqbfs/y24YfVHOAc47AgTCKfUJ6iN
AM6eM9nlThQNxEKj+eq1JrkAADf6MrGPCeqm95lNTrc70Qpq+iKZofhbcF9SLLsTjOCle5rFdZ5V
0gzrDJFctvI8F9mnzk+14g7IOJZrSjaPc16hH1hF8O3acsY7l9rXhPlbl8rmOV38P175IJSwL8zx
4R2Ltn2jeKdY1Vssv8TrJ3O/652Z9cXoysnAnlL0CSeqD/TNCEmcLjeX4cfL/77aUN4MTtAjKbbq
AXFcsFlVRq/pZITCjprLVVAHSFalc12MWoKYa9LdSkERNOnyymelu6HFt6969EbS5xLa13mx/OvQ
mTqwjOBhKOXXQ7ADMBGK9Cr0Z6JOVl11tfgcP4fS63IdGiMx/BrnBsuyUEnvZZwCS+W0eoAY0fqQ
VX8JShFq433tOeyXd85k+MSG+YeRvnjrOky0Rc/dMbzXR4TVMcaVEvbeE0pa0KIQpIqG61jLX4oX
/ZD6MINTb1UrL/C18QJi6gAPtfnlXE2K6V6lG/Lefi/zDb+kVEjCaHeov9kRBlvUzU0JcUuIC1Rc
1sf5venHLiiB+BdkAtOE45F7vXAKUprSj+3GY7Y6yF1GdQIWhstKQ7uv7Z7e8SBKgbZsBO7vHjdU
jL0xFq1klXKSYg5EcJaWGacuNDi8IqRbzgatWAoE/Iw3asP/2BpZkM1ex3K2sqEbpXCUknOxvIsC
tTAjD/crJpeLDMYdpFtE94cmU1BHOslnrwhm50rUHxfsz1wLCJHb5WuxY3CaNTUxD8LybZRKcCAz
fZi6bxEKybGHZaY2lzPbKlz+yMfGqGYgRxK2tIfHUunWc8EJU5KkUX9MWDZvLV7W+odmWbm0Mn1G
zocTb/td+v9FWU3+N1jEalbT3Thr8NmNcx0uq/g+Ju6G7kes33OX4R20rRBYVElEy2CffOOHok7H
78W7kIm0R2Kanw9HH4XYZtWBj0VAS9CJ26PH5azuE+MVca9Nyi2UBj/9iqyFn1XgOvzhwS3bk6QL
WyoqucROuWoguIYIN0mwOv7HZK/VcA63GoL+R0xjis2GqUXf9MXY+EAryL0mpBrcfvO8g5RzW3uz
0EU5gF1oieVfSx3pMIGRNR+9W+lQ47/SsBeAEkr16pAmK7z4Tj0s2o3SP5tdXI6GoUIfIlOYf3KC
qwgLRRpwQkbFlisyT5Nz93REQ8643ipMiu8I6Ux4BA4S7uQRC9m17J3gQfc10EChLSaojwsV9oB1
xTY8s9kS+sEU3g2xWmHWHJeoPXE2zIJnVsVMYHnHTHrEL4vEv1SYWlxZ2BzWgJ2ShFeyUOdl4hnv
VvjmuDay7df1DG71xlZvo05dGA0L+4XE2LJSzv5Bh6CMkrXXl90lRFkgXhtVuDZmTaEOq8jdG9PN
qtVcZoq7x7ZUwc96iS2DbvtdQspJVvfKNanDpWYL1Cw0tbZOcuHFWR+mZ4ysbBSD3z4/7CTeC1N6
+cGAxZCJQAa53KaInkZd4t7+1EnA0mcgef5rkyNui7gQA09BEaut0Xb1uaM0n0p2mw59WJhANK2U
73RqVJCPvSZiyKycV5yW3tngeZUGt4Zi2ulhR9ox7euMouNxsY5Cg9z9u746ugiBJimjPdeIKt2d
U+AV4kEwf6cOqZ9D5bDR03H8CExXpZpTE6b2cFKDepZ4nxGDAxyffilGzLX2Cub+X3JLYFlfkgwS
3AmVhzxnwEe+bhQkxGzTwytodcURML60uUV2NTcs8brWJSmy2LMX3lk5R/2MA4e9UH9S1Gl0jCL2
sfK+2daGYsK5NXQLh15Q/9HiAyvZXPSyOIzY9bpoI5rvaZiyjrjpY0jlQOEc4ptRCOHbT+YeYBSH
zeD/h72iwWyxbJuWgcFL2KLYqkV5pAlkkOJOhRc6yQPQfni4PWmrLhzVxi3LQURw6YrtA17Ig1cw
mL5WxHftXUaV44ivG2kOdTmNRcmxoO4gTecyJE6rFVFNptShFtnrL9vMHShq5a9gpxeSt8BH2tee
kGMI9xZgERwV8PNo3+glWbrsRVUWIoCTGWWEbqALayiIJv6mJeYlV64njeiAeEdAfBnzxagiPmxA
9MHWFx4hG8DdqTttzo19GWznKygUoc0XdUaNDuhgE1SfxnUI+XtLvctnZmZ9JsP2miqp1jdDmeGG
XUiz3+v44BN9gNGhzXo2hJH6wI5M12E/kimaPKtP8XitBqsui75W7jsK513gu4nFVddT+PVeOP9n
jDw2+G2o8yfp4avIDVAFzbph6CPrrYV2uFJoeJIJmM/Q3JnZnoL0qnOd1waJrjGctWNS0B76lwlX
Qb3XFATl6HiOJx9S2QTV+JSSPw7H6+ERTLECnTWfFsmOppxHohNcsxcMZQ66SnbKsqy53gYXTtmU
mafgPKY1WhWs3MgphO1Zr3rMIulBkDuOuNJbvwtQ5frbW69jrFVa5vF14rT2XiYs2TC8ERt+C03O
+sTLRAvswFyY+70IzDi3xkqiwc8a3EN5wSaL9EV3kI/6i+tZCho2v7lDTRt61pOwYfnX5NpNj/FQ
1+F++9Gb9YEhrSIrXkn3BilsROv+sB7iMwpEIcjlmfiAsTHDX5yVQNSUeMyYogwo7apaohG4Y0qt
aCQ5O2hfznYcY3qxeQFz7IDDFh+0FX73dTtXgGkRXQvVWSi35wNQWpZfta46QHr2bULsG0Ji5DgQ
5MkSPVcEsdqfLVoxtwLll+7A/07QZOvGLqEMTnYFXOVivilb6v8p1At6Ja647H4Lp67wBzY9vlCE
Wkl89fgdn9QFQ41fiDlwcGBPbIEn1RiH9LkTSLkS827gtBwEBy60sxcWNHB+58u8RIyeMoMx1NFo
P+ORNNXFJhNdcIVrsHMUFbdILQ6M2AyTRKtkoOxYNbsimT3MnmqhepAoX+0n+8YZVS0HPrRY264S
jVEnnidhDTaxqNZ6jwCaO4MKW0ez3PSU1wL+NmQML+R5Y8v9LOnaqnf7HXWAlLSiJPJ3Ykk7T5hu
3ArFnF3Cu1ncyg64bKct8olhT1o1Dg1bNK+GJQoRol8jo/2D+ACSwBWZtOgnxNZqRQ3Pa/ruubrE
hOSheg9tAnwQ93cOO89G5QZgUwFbUbASIQ4gfT445LQkIFPVyWcSNfKgE7DM7oEpyap5lufRH8EX
7IcuR99fiX3OMdS580ihydz+v3Gl/1lKGeRBlmxhZCn74OUioT7b3gi9edn8ELHEirjnvBXIN6N8
BsxTZ0zLGLMJw52kXPUhdB+Tx9H7aJrNyCTPatbU/ZUpQNe4RgPAkaG6/yUaWfpIotUVggeYVPcs
GoI6fTxMTiI+KS3sj+QYzwqI7XNVhSlbDLUyyMEaahHny11aKKl5u1pQS6ZSUGmuZj/veN2tSfya
ktaNPwH3FyALvik8gsZLmdkbPlkQlYt8kNlf/tN6PrJpOxVBDVhvfsMMCA/wFM8VrpBPvx/KMBKV
VG9UXXytGxVIfK+KbsQnz0iuhmIz6SLj2f2CFIdxVyimOrqwHlt3T/4lnUwRf+xzKrd+Uo+Xr8qw
1SVesRC+cz+Sk7a7Dx1vfgU2b1ZTisvoZP5qQE6xHguZ1YllgYAhIH+eOkTVoE4sNDDpQaREBcL6
8B65Bg04qrz58XdSX1zMn3vpk1KkR3rvKUAhGXs9xpINWQftyKIULU2t9l/6sFWSUG1ir1CSoahE
g5L1ihbFbH9EvxQbWEtRVlLlT3O+SyL5p22RmibNUTiZi5Zv7K5Qo0+XqDidFG6RbDJr2zb0AnWS
VXY0FGGGX4pkhQD3/Xk7/rrI5U/nqGvTCPDjXfqcMKOOWKiWm2oSkvEiLB+GdNO55ZbEWac7foKa
GStyukMJ/WxFlbqIqenvNGx7XI3leNz2ESiJMsDG16zkeJpdrNbfEX9khmVDvh2tNDjly/evsW1M
QWybhLdbExLH6+0tu7lrecMWdqcBSPSp4s4BhBwB2jigwDcw0lrHJFFdD4HlQfPirG6moEHx7rO0
ZHUbi2RPrnzoxttO8sfMoi6G1svoLoHwsb4Rh0rD3GePmQwy6HQSKQunCTy8b29gWnvDPkH1gPol
xup9BG2bHNimcLUqJqXeid5OcnjFWWC89/0aIYkdHElHGVgUD4o7qSfh4n6zgaerQAs7c57/vybk
q/anpLhMJrBVcDdUocmCZnt4466OUY9ASHv6WqzWqSyuDCEYBxMPWruFR9Zer0O3CF4mthdE96s1
ackJVGD4DATuIx8LGeLGBwD2LH3nCtMFjubAL7imy361K4ZBDgBj9839aqhgnTnje3nBzIwPNAdY
UHblZqJJ1mRYKgWyqPZL6QtZqxVfFGrsRAJG+RRoV9NqsvDTvDNO2xDQkvQ3NOsuEwiPoa49Bb7U
36TcGNAk8PiErHhXUgdjypfIsO83B50Qnb4HwSFCRwN7CcSZwegaoHIo+gefmOV5lj83WYjXPaZT
s7sQsD2bH87eMBAQBg1hc3IPVyDI4siBwt7zHkhyoqoFt22n6HSvpd5/bCRnf7EK4eMK2i9OwCuk
XpJ3hDbGB6/o6mVXL4MqGzpaFDq7nbQfSKd1lehtUjASojAYcE4h/iGggfooDkpUgrRTzm5y3jg1
Tw9u3T1bOS6VlgskCt6kF4a8Xky0LdDIt5uR/NkY1BV/b+08Ejg7VVS3CLJtyQEBBXAPMMCytceB
hbaK+p92xFmr8IDqVsXEhDMK7Mn4r7uLnAnKFC7G79qDNr8RGkJzwEdsdM8Kwh842OD4utQpsk9y
Z9b2KC66zSGu4cmgEDXwJv7BTd0oK+hjTaNbzD/5yIpXqmEvOOeIASHVmUACHxtLN543RiE0w8z4
/VNKWdi8/tpxWgbRh5SvXFaYm3UCOt69uBaOFKVo0/JdtzbREhmWtHxjBZdB89Tm70NyovasfI0Q
N//FP5qDSSI9GbYdzgN7/US0qYjbRiat50Tqj/AFDI9PtlrXUgL5KfYdsxOW/o5BMwQ4UTQK1QaZ
NDP1he1l99tS+LZK63Vrn/Gbnp+VhKaQ6SKY/lIDPjB/86cr9m3gyCGp5kjLns9Cu2bemkZPwwd0
4vqYsQ4tOH5951CaPYPp6wpbgAHUFakqyOFKaeoQuELAZBA+FHYb2AcZ72A69GY85FBXz6weJ56k
UD3xkK+LsPMwE8Rvv75McZiZd1XeL9fwWFM9H2Q4eqwOZdJtVVZ5DnrtP1RlwJizxYCXi+U6V/Us
rAy+duf76q9htqlsnd1KZ11bbNDYU6d4x9hn0nqtmKYw5a43SU5YMRHqy5IFL9EAtSjVfRxAEZqv
Vy2qRgMR8iZV09ZGqEEGiUAehwhP+B5vgnK1FP5jvSTkBzPA3+jtVkWfuEaqD4ot9XmUl5EbpCkb
fUKcLtqklPxaO+HOJlycRXKlN6dAu6J6kHfzcyPyuY6cE1kp/1UPfNLilQ4VIF63cIoDv/0QhlKa
Yss24WBdBhBesdx8QYX87z9MBz/4mSjdheUk+QuFVl96hY9CVnAPXiji9CzJbS21bUOf4MyBcOoC
mTDDDSfZSuwp/LrQ6LKlf+ZRE28PJol0YmO8JvZk7DOE2S0lDk0+DKwpdeW8lwgnCUlQGF9xA8Ql
6Voajd5+zNfO03lj0AmE6aII/zy/6WjfLloDq5Y6k5u4oNdwZMbi19t1kq9ey/i5xG9Rve0Qu0Jt
6ozNnzdZ4p04i7lqNayS0LSRnkWU4murA8xm31SZlR44ASa4OXPUfZh5xgZvOu6nPHLwX8lRAJWu
yHqN5Pq3mBP3hDiLXLHER31oxKyrsdGLz7tME2vM+mo9003zrjVoHFmTHTPT1J3btEsZE/F5nb2x
zBE5eZJmwbDUfeYYxatsH+Irol62dcEyGEKd+cD423pEtXsvjVtw98AUIk8AzdJO1U1UDy87RS1s
EWHM/XNhM1BVw8zxZ9ZbZac6IBZO218+SjcD3g3Zor013ldwpvuMmC6mcspYd0qYVb0uVFTgz6hy
0aZ8TuWE2L8Ns48zOObOkVElHWGE86TVghb4dc1YQWlx/kRZd+sbC5qpZESHMjGogpo6b9B1Sd93
9CrPPNaUos/1CnXFyK+A8mU4xZD49cC1npZK6ekLdhrnrUe8kc5o4re3jpJRQU8RndeBx6m5ws5j
JhA/xgMRRNMy0BVSd3K8NDPr0g9/ZR2YxEDcr71yXVLfVQ/nm+5DGVwWJ505jGXra+3N/54hE1Hz
47vfMyPlH8IwiTDVskJyyVO/fAFwUuEOUQW41F1bZjibKaXdq+vLeRgLDG66WMKUQs0HXDEYMnov
ilRnYAW/iZnwA9h9+QBo163rxOd3SIT/82q9dBmX1EEgx5fUi80cVyZWV201n0T6qOmSzmNGAr6I
EHr4QO4llxFBEmqZtMDXPoEuI7f4TxEy+nY69mAtNXTLZgcXjjSMDIEHxBF1U4Zqht46zZ0+hx6I
GONH3NqRpdEvr6Kay4VBCioOi1UyUu3boV2Z+9gqPm6A9ZCv8TmzqmqLG83ICAfzxleDJb5sDic3
mCImZjVZy9D+EE8dLwMyqnOhSKqFrCMSPnXBhY/8yh8/wQg3YqiF5FLmwvhhTEvrPmpNoAUD5Hi7
/3wRBd45NMRcIItYPBtMs7gV91deQSUhnCQ0gzNspIhHHp5u6FATqDHrj0D21i3CN9Qv4QC02VF+
1LszTK7Y+MBh3VV4mfVMCnBEBCkNTqzcVFfnHSovbleCYgFs8SNFW5bdAcOQOnW60QShIPMpcQGr
KEFQSvQpnfLQHvcUkZ5l/bH/FoCHG2/Z+U8fmHGO/NwHTqLYgeqYQ2MKYpe3TQ407LX1TzN6yVDU
EOoxBhViqidlJDbSo5W1Fz8ObYTsLtALaPrit7Pue/IkmuqAYYLjVHeNMqt33jyqop1ikC4TeGib
fvHnbq2He/vF+jPlhId5Q395221aPiwftR8Jzz6x559WzWOk1r0n3Y1jF+6TbdnfHFznQdyftcaC
RKEtGxJZybNlRD5L4YElJse1KN2+gsXs/0Q3t6RjgOjeinB76PKwRDwzEvSwAIdlQjHWdCtHx4v3
utHni3Fi8zc7jMEsldNHe6x4gspfX3Wbl1ifrbhYb8Qxqsk5j9lhBG/l03Emlxr/Fy55PKqNWuRG
u5UZs3sR5zHngrwGOyQqgQaT3PyaOCPbqVZ2b4b5ogbY4hYasnHLCe3OrdlO55bOLsOyURVEIMe8
bQHGF0/82f1yaVPsjzUlQA++h7adjjlMB4ogoZumjXEmsVw9jMv6KC4Nj4OtYfHFLaJ6BgvPDSp/
HbZ2q8w3HLJ74nme9eOdIK4ExKGHBB7eJU98gzck+ARegwwQHgcaAWCdBoZX7fY7fKuAN9/qWHCn
t0rgBZ61RbxAOSDY9qYmqxnUKwBRoiQQvk+8kYLLGUEBCT9imHmj5B1oR9RIuLLSBCw49Pr5pp5w
kGcXGuRoxT3cWqwk95+GCYfWwKrGhFDjFDL4405ZyvTfSD2g2IEYcuGT28DdQZTsit4lV2OIdu8E
f0f40EiUZPAZlywrsWodbUzMNE74ZhKNjT0joP1el1sDFWaxUpGYmsrVYsRlnxqG1ADgupeQFbnr
OfJg9B+qCJGvNjMtfzc/P9gyO4Co3zx60g4n+CtqfTw2K1yV4py4wLKod3q2Kw1Ofq7EcGkNw7ha
WSjiqQcRuHDfNhbpuh2ApLADOhryLSXo5GpdSK5rFwKWlwrywKbXdWsuIUNftTkeaYsCnokR+wKC
DUxqBe/6Oa19TCYvCzuHsyegx2gJBRW2Cwz4LFGxhJijIyU4rPCCljCaDfX+FdoBFRb6xeZm0RyF
RU9DaPuketVR2hD/D6FKtQZh8iSPrje8wkIx9+U4xRgW6HO+zlcZnPZKxnGirhec4BsCg1cqgAgL
pWNbCJcsVoEVu6dj/5PYkSAIuCKUMFI1CiNAxvCUx+WeRs/ZJu9RvJwkZl4596IOW7rD9wRzy9cw
sZVXPa1nLLSw3lmYWUQ1ZTc9WIDtfKQ6NYU5MfP1jTAYTpmLq1bi5d4G8OsYydtv63A9Y2XSKflF
wUTuAMwD3+aYVNrKne9aE/wtHi6Yt4B6pdRiQ1fQpv2Fiq1N1ejjz412DZ313HqITn0euFvnPsr6
p699yeyAc1cgachsrESNl9SD/EltnPiYDCRWF2Rj9+Ek4rDkPi4nISbkX8hzJ3eft+vDf7GCl2pe
reLpAoxI3ON/goIsfckROrPNunHFgiWTnFPcUoTuADfkkGMtbODMN15xqC69K/Q73AR2VC+BNJms
WFlghT4tb/aVYpAlvnZIYSoK0RA5sX0YucjUYpkTP0quethd78aA9EFLsoPHCCUOsZ4CrRHrKP3o
CCa/P3KF9x8xxbvxp4/C4Mp/MlQGxmT14+VTsctE3CNWYFRquU5MxwwmB7H1qBYzVvoP1rTuDxCU
ll6ljD1pfXSFIljgPUEu+rV70ySGpWHsGcQmGpdv2ibjLA1+P2vqDZ8iuPtLlGrvrNH9CAk4zdH4
7YNRnY7PINgPxKuq5Qxz3RxUNemUDnP6ItuCG0a411vRvHpbtls+ig5mPD/LUbwX2w3lw7N5Ij5C
TwF1vlHPIghqMSeTIsJyiWwo2wcbWms4ajoCnuC0U3oGkfvHkXpGtdrtfVIa8paazhDczx3FNxU7
rkLZeXhrPb4OPuKUJ1u9/vhfpy/3m1BQS7x6hKGJLxbv70G97TAONL2B9Epk85Fy4o8xzLl4NGFw
FuQg5tCw75Z0lIOHMnzh/9OOdlmfhYiPq1kXmb6qZGkFZZTLIkUZIFkFtb3iqAQo5s0+PHhMJU+x
8IQQhO0ksc3d2KvA3hIPQqg6DHjcuBRHOy9TVFY5gim7XI/A5ShmwSOMCAI9lmvOsWbRreKHaxuI
JPUKDyGTmpdOuCZVQ3Cf3uBtumhsdek1/6WS3b8qUb1QKKM7Tlrg8BytaF98hyKYAKhu8lko6uB8
pZesBCT9FvcuDXfEgckEQZW0QhIfbUmfTlphLi2Sne3uFtDvfunx/ilApXAwDt40M5INfbZ6FLdl
WbG7VD6GJHleSzeL9zA31nrfmunAi4xX8lX6SptWNT9aIbgYKdXMEuzUqxrdCCch/unsY8UjIL3z
0VJDh7REuRlVPGuUEIQOdNScQPybYP5nRqesc5IP8hBtMdSoF393ffs8J+B0UV3Pjujip3n5ZS/Y
XuPrkOmOR93+pIokuziCi+m4Y2eAsPIlqNZbwJnWt18zFmaStp+wDtFEwpVLtwCHzuWyUHuND/k7
INJBqNvb1Y4+Naz2HfiK1GDgej9lUE22ZB3fu1xadQp4I1JKbPIcwpQXuS85y27U9VoPKiCHbfpa
eVQeC6xWj5t5FR3v1LdCzsCJDnwjiJInEZbPQT43hF1TofnU88y1prgCEA6tUFcB8i2k09Zt7yB4
g/o7/wHn9zyoCt6zfhHDE3pP0gpeLY9TCM5WOo7Glty6qVs2cgTuT+9FkTK0lrxsn6zNGyzugRk7
jl1+6GhBx5S3SyB5oLSGUykQtmLQK6rcT35G3xDclIIgWYu1YUYf3TnuDYgROOkgdE7rFBL6PDGv
VI+p8MVQjfd1cfXxBSZPBATCidcUt2kr3DDY33U3Ps7MpDfCAWaQuG2DDP+urg/0SsE4Xh+oHShq
hxVrLp4NrpNlgC8VkkPoBUUN3N919ZCxF21KGfAAy4PI+udejDYRh29BQLrhZ7XKTjjaPCyJ42Wo
cRsZkS4//wP+rO88ea+ZRrevQG+Jn1z0kh6hZmm0KgcjsvozpsEQ1oP4lxylpUAz8Tt6bFSH1NNn
dQwmQXHoHS4C+/ryQowXVoD0iRV+JmsnxJeEpe+os94jqaorWBcBwlDPeVvwOmXOVMGvSyQ9MnfX
Evi8ZA7r3FzKJj2PvbypSXQ7n4nF+Fdt6MoZLGX9KZfGMSXOO6AgIJLcRUrttBFXuDy3IYmkPSJJ
jFYVVyub/LVwefUH1FWoaEBJUNt/w3n9MuDzfgSfPm0nEE+/dhQtMiZvmhRlLcFDtwcoMc+yI4Rr
NFNk/YDge36U89rsK9bon0AuS1FnI8cRQX85/3WT4AfbTvTb218IN+3xJukiwa5saEY7+pGy6hSF
njJn6x6tCHasCCf2LEaMNkYsvsHQexYAhfllVAsYKm12cAhXYNFzCQ97qFaPLxN5E6zaOIdslGJL
aMoeX6GHILSoA+r5nOUMmmLKa/tk1rYl2NZRQUKNXB+xFIY741iIsTmQVKhPOEDUv33MuaIbtQ2F
c6tG7coWMqXSUrTUsJZfhEV/mTGnUe2mfN5tXcfF3N1QjU8vHkYanfa09gR/CAoke3y40AXQEpYt
inzCyDY1yF7gaHO1nBD7FCl26GRrxuQs7G/fTc6AiliWYjR5Aenk4N5ekr7FgzuVi7JQ5/An1Kpp
ArOKgL6QADwT/qq8tU3R3UCJYHaOl5hRR16SlrCShNibQW8eJ8PEIbgTcGPmDosavjjE1XB4JsPK
4aNv/pg958IKZC2+sQoV71QVRt0pryVbIZ78aRcxmUmG6HQsOYZ7rZvCaznBGVrafB0ogpXy+GC+
4E78BzDNdzq/RCpA6e+5ka9cx5Uu6Pz9Hr6IP1SSVyvVwNq8lGCApaZKUTaStwUJKmLDiQ8uYLsu
amREnjtSL4KHTXFIzV8jr12Wy6XDxMn9jTmGYk8/GxmTld9zGrW7DxbPQARdm9vT3glcLmrhw54q
PmJEYUf7Ed1nBtJFdcihSfEl633mk+kCJm8ZRKg7hegFsvyTnHLq3iQqb4Q6WK4eQOpgm7/om6rH
LgiUZqNI3o6n0Un2WXYy43+yonbKJYrcoS0uNCE5L42idTjyR3JNNroY/IiO0IUffr4nMjv0HIhg
tyUfhC3V4kOX9G7ImMDulRdm3+TZO6yycq8UAMFPm6sivMNpy67BQg53cN86tZxP431VL20s6eqS
soT7ot9EihEUeHVn78W8zV4pCmqvxgd8lsaCfgkSW/jhdrr49Wi9yLwTMaa3ubpgkZRdCYFTrV4x
mV5/HJv/M9NsoIr+9yQ9PAeGv5w/1mISe2XrDZ9k8T3JyUmX0lYuvwoSTZIaDkrKAZ5tc7QfGhqD
4qqqxBCB7TyMDUTjaBBaJDuIvLJNQDxO4QQe8/pHoz6VNJ/rw1HufYQGUFuZqOuprbdMCVOQ6fpP
MPQIsNplLxs2kGvbmHZBhZ6KXmLfTMBj1C9KMat9xK5oiZHoDrUAAfFTNnljNY6pbsRKkuEK++Mu
UqtkkI2tmG1E3MLbwwd6ZqO+HT6NqAA9jvLUtU289+OPqglEicls9k9K9ONAE6X2YJVnfwWgN5c2
L0UYN+IxUybzWdalBDH6j1cSRUtKIwueR6bvsdpAzNLIesfpiYfby03YvleZy3YHAF7JZvc080Wl
EVNj2CS7Lw9XfgZCRYPgX4oGg/x34wMArC4UIr+sd09BXLYSQozsc/0YOymNQB/oKsQMAIQzz2b5
oC+tbtFOCfuoISy9sXQ2HiRx7j8zHKBy7KCKAwEjRT5Es/S71lQG2YABEMQHKJM8t4Z9rKZySxH7
c7p6qqcGDhXcZ8tVYPCWCDC6BFCVjJMHL0+SgHvxaciYzBlQGFHvdCDx1fA4vgCnIXNy2KtlrOyL
8oKVDFZEvH0LLG0om5afd/Mxu3SxM7RC27+7CcizqcR0pOU7frU87bl5xGrv4H5OQYe19G8dNfle
kWPCt0xQ4rIf2eqQUFBIOZkSbUe6+xwgLwvIVxuRGL1hx1b1ILd+PneVPif9K2MZ+UzV2Yp6SBd/
hGn57F53M0plY2JBJa9PW4rPb7MUgwtFDIO6ZiYqIZ4u6om8QHCBhb0OFboKAvLJPiGk+MKM3c+n
+JdNaw+7vG8KSKOG9pqbFlUCmKxXlMzYnCFbMZStpWbBeiJS/O/l/GDuIDu2QkoEq1Qov46ZwNXP
S3Q5Tl+utHVEwd6QYhHNKG+2ypFDEPJEVQUbSfDrOkoi3d1m1O9wZKcsXCdqyJiyKw5ZtC6LOplw
N7YlRYIiG5RlFIZ/fAlwL9knM4WZrRJD23e6U2CZKQWsY8PdXWFxdAYr6v3t4TXmwGmeLU8IgVpW
C54KAsWf8uObyg6lC54TIFb/YPULt4nc44qLKRHc27uN97/vQZiTprqN6y6KyhMPJYALRmzEkITq
e4xK5t7CPjFhEMuWqoKLOCznwg1aww1Ch138vGIcJZSE1FCx9GLrZoNGpPVBsUFty2GtqyfjLHuX
fD5/AECzMR9DK5lw1ZzZ084xuUTqeKrX/sFkAp2CAishYNi0Ee+cBFPisrrNPun7NRh9R7xjEJBA
ROdRL/pbwwOsXsuKB+FWF3vQMlsXQ022yXAib31eAwJgqLVZ2d93RNCEKBSgamau053F3BX8Ttcn
s9HkQr71IrD+NW4AKCK61Vdi2O2TJIFX3MHzdvGaxxk2K94ededNbXilM0UeQ7V5ople1b8yvwd8
zFCW8fL1qmgBoZAlcSd6cGP/JHhRkMtQevqPK3Tb4VSWA6ecfs0ryEd0IlT4iXCnxHcC7fN9c2Ox
ggVFn0p42yIoTsF9s/n6RV4lMGLPTbgxFBpkjV8aCxWKC43BvuNxbkZGhfq5RlJduTmfirDqa9JC
S5kOWmUMXM4MP6LFuUhpguS+ZMHBEru62VC4o+C1MDIl1OWaAkH/JJy8/jHYFRyTcSnHIMbh4GC+
6x+erVLPZRyp/r9mzc+hvqf8yF33iAr7jCtRBf2PE2TSi5qWO8qmLQlzLeBIYPIwpFna5crs8BId
U21t3PW0iCHvbk7pSEDOxOggwdNJLlBCTXS4/ubpvAS8pMKaYVJSQdrkH4rLQ6npeTDyn88cvJLT
El/2YqOGCSO+xMSG+UrEHSzxL8VNUs7Zrdx4Y9BU+C3WxMSfgy+Y74jXBivKYjc5NlBtrV3U2IDH
zs7XbV60Yns/F0BqKxhtJA6/tr54ibLjqN43wx6toAodTAi00NOyAML/rJTHlIbe+1Z1FIMmF0LV
aNJVyKwQYsH+Lu7i13q1iCtpfmFmszE9K+xjo25ZPchIc/WNPV+g9JfA6TuFdfH6C6r2SxH8eu8E
NLp7Q8PMh4tLTozpfJfeuwAw59aDr1tI8nqiSFiXBqX+M7+SoNRQZ2vmWwBGriAc4mW3tDQbhmRa
qmpGAVsvcTdY0ClYeBTuutbp5kpj902y9f7pZ0ZhgR6ucbsdfudz/dZ4xZXNolpdQn+5ZFQToX5U
tQBGuMD4XRPiuHJNCCZ+o+mC6SEDJMYUSAkEJ6y6OYFOp95iOGMdnrpds3k6cofumKDdlcjJqtwA
2E1eGMJtfFbZdwujg9CUpDG2p/NKc3YAYpfHyPNxG888ibXwWeIhaJU0n40vs2CHJzIdZbLfpEIR
gP0k6OF9qW0ElIb1MKJMwqrJaKfDLWn/Tbu/sCVfaoXqqIKHjml7u0H9fe7xxhdQ3fkgFEwYiFOq
gEVgFejx70T7W8I1id5CPhLDn11N+dkHznqelK4BQJ5+17m8dGPVtK2RGQZiGrsQ71sv9XsG8Vfe
1Svhmhg/IYvjAJNn0VB957Kiy6PX9IprDQLE0Z+O8GgeHTQg43UzwFdWZ4flbHP2fKDrKPXRSV7R
Z/RTRT6ubBeWnMt+9OXV67vN6YDDgclh+hYc78LOL14xY1gR7Zb5tkdwqtvjnWpfTKgGmJgnQb4m
YcX8Rae1Gy2DSmOmodl92QOipMxD/z1SuOJru1Su8QgEHTVKmmj6rst496ljLd0krgGyh3WIzxRZ
nwhsetABnPnLHwjoroL/lLipJy8qrAjobj11hfADPSj1heK1j6oj0uhyyWSPeum5oQ+5vvn+thj1
8ofcsLHqXrBgbRBTzsBVrtxOS4P+0mKc4ZcVJLmXv1N1NINsWPrhfw+Nz9MpQ7QI441LJvPKL0gq
6sak3NTX5rreTwsLTLqMVpDdMQRtr6SZetD2w/8O3KZUry/koCN/MOH13VWdENnycU1MGgyPrygs
hzuRDlfEyeoIdWHIq5zuyCrHAhHfYxotyy5AylmGlc3Qhv6UsK15ENwhgLI84VNU+9i/8NUis6Rp
zkPGHITLV1pjfPyibFYWjZC0CHyLxq8WemvPJGdr3hZCYuox9PZlAmuZv9Mcfk7z9ZlZlXMsWXzS
3bOlfTIWSrjYPN0MpCXhgnewhqUl8KfXzzw411tlwCz6WOg1kpHFBLPCD3jTKga0N67GuL4Bi/yR
RzpdkRqR/ww0K7onKM4VKW/M9My3VjCNJ2ng3x16BR+bsU5iQ8xtbQoZyMhvrIQ02zrrv0M05M5j
goI0SzwavUDuzs+cHsGLRo7U+oBOgup/WL20lmMqAzt1rEV9ZJnnXbxfCizCois/cCVZuUfYpHaT
VgqexWT1xX1S+7w8n4BdmDIpDzDdVxT0cZJDxQGDVjHZkKgG0nBDqjwQY0rTxGJDbZocT06VuXXZ
+kpoVevXGrkCCnIIB6uc+D5wEMLEqWgUKb76QcXf+GUz3PYi3FLQRqeyKUt/7dPLhT8Jj/PEt1tQ
+q6lm7kVbVgYwJvV7O4joAkwRpOaZBrqWgbHsTrgnb/5pjhOoK2VhUIpAzsEca85NeQGBu7GqDdE
JPjJ+2FQ+DcGDx7AooL610hWbOZ3i3DyNma2B4Tsi8bLzd7QhAiXZHNT23asg07r/XSmd5N0C2h0
i19+5Sk+8gP4Q+yIeE3GcaNzwCDJAdMCIeiWO8yrwhUIPqV8fwV8RtDLYX/43Qasy/IxczkhR2DZ
/BjwtHqJwzTyUQZam/MrTQEkPaVB1+9WCEiykWaA4+/eE9YFlU/CUrGUIqVhL0Tk//IIOmV+2Hri
J/M44XNEN1WG8QAkNJojeo2Rc7aKB8gjoFxn5XeGnyioLaSlqrX86kZsAHtaVSGLJenyuZyzZTdI
hgVzITuNnfOlqhxNbV8e+mYJRKXbdqxUTcEcdO5PCL3LhgmEl0Lnjp0XdVcSc/xYrmYX/PKJvSNm
00BwdPugxe+Qer3sG/Rbc1sRPJdtz7pT+rfXZzxUxA9IMLq+pd15g36XK50YHHbNIbSqhup+z2el
eLGkyTg51wQyyOOv6L5je70rfV6dyNWVvwavJKSFXZtOQSrIaYPX/EGn45V4UImCVLfvhHdyyVPJ
hOgbyedrKwSodfEyuKDTKU3FxuJ9oNTY8ck+XmZUIJHUueAs2CCCinMNrzlCC3zPn/YxBxZ9oOZ3
EovBfsF7GeMEO5Dg5kvfF77sAbYMge1f0ptiH1JqXzsWCAiSOt5lB+FKx9nlkhvFU05YTVID1cBm
WFx1jOU439BOCcHi+/nr4h4pqICnw420n4laCFnuUv/TEXUFrNWqgAdwzCXYXoy8zBsy+yA+/uY/
WYaY6xwHG7fzvdSBdTjFq5AS/foXKmInj0Jh1ANIjVFZDlGUATcXAFUwiSOOFyrlydbifBxyyNkp
mx7rez1aqka164oiNCqHo1dnnU8TQCPLPC9DiTZTp0J07nE4Do4TeMNzHec7u8zzDJpIa1FGVgYK
CpHnsAt8cmMLXqQrpnX7lUAfR7tlS4GCYVCDzDCxw+nY/bRbX8U0qHhQSVwuBg0m9hrlmw3pssC3
nsy0QW5Dq7EahgDLrsrBhJjSMljuqyE1DjFbu+/3GqTaogUejsVSfPpnE9acFypzi1Uad54H5K3z
efETdQ//pC37bGwjdST1L4hDqbOCO+6FY4+UNRZTlzpLSQ4csU3SVKYEw4mN+qTLYpbCD9SYerq4
1hQ3iqICNcUlazqO0YzLlTvVqLOcLsiHCXMagfaH8xjNUjd9Qan6lZs+ml5iVkPwGSo6br6DGjkF
syDbqMNqUu3lyhpAjgfvUINdwHCgpnSZ78F0acFMgSCq+ZPTjBL/E36KIfjiRp76P46KxIyxiT1f
qgT0HQbQhdqL9cjNMTfFrFrQzdQ7m1ncspm1sKOwabWjFlPxjRZipqmWZZG09qVW1KjmTrFzngC+
BupgV3LUiKWH5W698v5EEfzfMtHoeid+hLIjf50EHHyaB/qD9fOZ8GYiFBOBR943rEKizLgGDhNP
YDVJWFXRQ2JaTW8BiYa1X1vs5j7E47ZR7KGHGTyWAE7H5Uynmp/v+Qc2ri7RFImGYbOkhKn9R8+L
HmoH3Bq3LfepBeNHgWXx+Bf1ZUrpa3Oy7GeEWeUXFpzEGli7JqdPuP9h6yUHKvhbopDRhNLw/vp+
D1hbi9r+oD4zg12J0tus8BFrT5ytw2XGkGG6Y/jrZudQ30uWDYm4QRoWm2QJkqt7TYzatdncZ9Fs
GAAIIo2e0NJdw5yfI5FRgDcetLH+E637Huht2j6b0baSZnL/G3HDZyrRtkiepmAw92axMgzr5vgv
E1FmwsSFrz6dsAHRqLbxlVf31cjcySErxh0MahWFFuOgJeNBJNwaDsGzNAvmXyEAESm2KZZ9rBf+
s42BGUbwWyRBH6oHY2BMOWcGEFqz6RbLaEDtBs1KGE9eRwk3ZasJglroERj2b6qccRWn0eT7F7nB
bZV5vIooSgC3Hm5KHkFInjdquI/QlwZw0QGY+zxlZd3mKfyi6x0l9S+s8AfSm0BsHhaKfJQq1FO8
osBjEoucIGX1HkUvCUwyUVDeohj/84CixvdYmvD5iZBU1ZrLqFlY9drkuEtTN2PT6VjZl0bXEDn4
bQqRiG0W2OZ+EBdqUmwYn36Z7JXQuWwZLcUDaXLqVRlZrErR3+xhl9sm9QKArr749/3FdWoHslJ9
SqPSmTsLWlGZ+C7nn4W7/JgZBTC/+XjKtGg9wovC8sR2413XQWUfaGEH7eFwK3ciWehO5577QPWX
yRWIcZ285/ExnPEH/dwOZ2jgnsjZsS7gwrW38nhHK6MMNWLs6EC93xWficZiwIYFenz85pmk6M51
wUnpFwwmJd/ZUC7xakK8pv6bI02/7rJicYyP8CuCwY1QAqyuK0jBjEsDkxS5V5BO2Nxl4HzQk3nL
n2L+fPQzBMl4Z4+A9Qeba8ODA81aFpsiV9D68V4wLvbTJCTc1ed7EUrtYQhlC5DYjERWeLPprQlo
VClfl46KwqvmajLbHCEVRdMQej/n7wDLnmPSO4wOa+1RnGezyoF8gookwD/LVI4LJtxKEVZ4hdqr
JNzp9uTRmvwSzJD7FFSV6rUhhPbf0jdaimfmBs2qA5+v1bZw4QwnhoFvT0k/le8S+PE8RuLPfZ+K
2BJs3xovbiKJ3loAFFdiL8NPFzYjCnYpUqlzgslSEOScMQeQIJx17LtM7UkdDkRmmiv4UAEMMQbN
r7Fi2bVfz9570OSillDnkKU91u36vC8dCITMmwbEGpUyQU+ijhFPvE0x4p8pfXZ11fCaf18sO76s
QS42AQswCnR+2lZkOXZAx9V6MbBjPL0Z+bkqS2NXBcy3IDb8q25ZpMH0gLK8HnKwyYT1dzgyNVPh
ZQj7U0Quz1/pErMvydwRQN0ikNP1ITc1HTOA1q5T1Tx27Cu0+dEzSGDTpEJePCjt/8KirLQm4on6
6B2WbhTzR/Q5ZL2J+xKuD2O4MZ7Qrebvfu2d05Qm/u3naJci70x4Qt3/Re+ItA2xjmSmq5rBiaK7
QdHrwjSsbzC1pI3fKK0fBDCRiusiY+C7lCIoUdMIEHmblHCQJAo9yQ3nQrkZsTIto/Diw9OWOUpI
QWfzXfekvwl3PnVA+MriUd1y4xBWrAO8llPs0mgBpwHm+kerdr0Uny/kByUoe9+Ecr+Hb3Oijv96
+HaNNCei3s6KB/iv3lff9xRhcoJmSXXQBBlkvBwI3Ed+VguAxbINL8lOIGtHGDYPqMI2LTgGJ1gH
M3PIQdEPlTkqp72ExkXL9TDLsLwC/sE8SSxk5eLbXQVeKz55UT3l72axJiuaTudL4vQAUmacVT9s
ekWkat7q581BcmQ2a/lEkHFqa53EKf+LrHin31jJSci5741P6xbSi3hjn6UdXooDGKocRRWo5pFY
U8MX/aJU2anRoKU3jVH1GKE9lBN00QVES2aawQWUZzYMt9HeaZeXLG2g9aUqC6KYLZQ6ECzEKKDq
vK/Y6gE2uPbmn+6OgVfPLMeHkWA1iYmKi6+NDOLtHC3JrAcesa+2RswToAB8idggBtrFxuG1KPmD
a4EOzPQ/JD+P0DyWlyv8/AKtOYTLcxLmJKBmqLSnHKu2jo+1CfqUZg/eG2/r4jqlE4eSqCIGuLJ2
10aUaDt3TEyFWBrdkn2VIfw6OTUXN0vRU61YShuYtcA1TOmC0GEQeY24I/MqWXqnZsFNPxVrHmWe
PWkmV80Zhi+uXJb1pAfp+KVKvyyTSI5YRTs2bL5fX6Ao20BSm+zCexEEMAFIvKMkq6VwTG40cZWY
RI61BbU1NYQWyNitEoDst+01+GCtkXfCauv3wxrD96Vz1CtHoAOGIeFLlTxsGzLP5RW6gtpu7gX0
vDzS6oIHA/XaNF6y89rlcrFbQkpDQUz21DAchNylDFeFalEsYHC4XjODSdw6R1PmFGnUkIWXiNic
psdwiveZGdFEdmueLDYYgFfD8dhhYDYZr+y4Y2uFGSiypVTNrIccVK3b6UG5D/zAnyNcixJSZfQG
QiVCUH0BNplC/U4JzEPitSpFAaqObdgbI5DN6eZn3YYXcqQj3dOnoE/LDrwGcosw4xv/HYQ7uyME
bQMhkH3rV7k2VVLVdRFEchohZW49ce1ONf99cC4DU/b2MMIOe6AyadtK5aqVPSjRIsS+DDSjums+
FN7gw42QnxXSACzUdsr24iKmiaBcJIRJA0uUQsScgGwsDRTOpej3b5HdLBIRys/pvtluEgsojAhe
Ym1oQcFGosDstavzleAXy0jzlEeKYev2dPeDoJOeBrliqFsgwvijXpcj1glWYjHQPMJ3ZNkmFkG8
LVMLM16gRlBieoKIRSngg83tMAUD+YD6PZQ123xlH5JhqF+mqrLzzQj5iSvNJbmJu8okQCB1gtWw
IvK2Wql+74pAV1O6huDU0T8DBtqlouASRrdXN7vdCulhOpOF6QNRBUXNaBM4O6IfuvEpeza34dR3
/VevJKoefxAJuszHKcBOIjTZ1js5oADDM4TD68e73ukZ2sj7o57Sj9Rv5tj2UQGyU/7gFjwh2BBJ
23F/A+Rjpx5Z5IWF1vL9kbwDgKl8YAnLe2Ivx5Tm6sfUVpprFEt5jjV3E1w55WmC59IvWjLeIPnE
mD52rpOsWZC6CzBJb+DyK5uPS0RJOS+vgyYaqbc2dUZo+cKvKHXt0rz65gHBqBcNQ4X2nWuyWZEj
r1kiXgC6tWrJPzgP6h8ZnM6O4JxDy6PKxX9aCBEVLxT3dFF0atJt2Sx9R2l/cYIRLOSqnkjqjIhY
hwNC66p1vk/5ekaY3/wT34MbM10S0kLY7h4dX0EFcPkrHWcyC1WGRgHY9lnCSZG8v62x/onFHrMe
kVQqEWsJfwgLKclRxxlL4tHGEBjZlyqFrtCK2wtIw5OeCHMX/lGXd9aJIS32KBHYIV7eycc7iP1G
VLkeu/+UhTNh8Z3PYTNQlu/mwUDxp4ErdRymTEqT1M3apOHaFsdcMIUsSXgx50nZiwV4hR2IIZOH
cnkdwDAK3dPMlOT+bnZqrUWiq5la7/OQup2mKautFkuF04qmyT4z2F6POl6guLgg285OnWsmUW5y
bHW3QeM3dejlJe4gHLLeBGgLc4n/fS6/10HIICDBSSt4nLDqltwrq8yQ/8b8FfPMm+mI7sUqGkY4
eOZIUdPu6ckwMrwWVw7AJipwHmJA0y+5D8vfMG0BjyugGdASUEklxGko4OOEVmfg5ENqRe1p3B1/
vCEHgvOEHq+oFt1z1MIBiNIhiG6csFGj3Y0h415isqGh3r5FwU0jgmKn4fxCO8LlUNzqTrvsQjQr
FF/TojCqrf8/CojuUIU3gH8FTbrsEC4UnxQlZrIDc+2IyJp4OIyREA7pfTznZddgMtGf6HlgXygs
k5/1jMo2gNBuxE3pH5Am97Uz4lODf854O23kC8Zw4RIfkLm4KLJ+dtnipUjtG1UOgkj1KUpE9fxC
WlA+t1c1as5Hyz9dcPK7rp+dEXnlKupWsJxhWq0gJf+QcSSl2WX4Mt2XdGA3Ry4XQ120LdAIZyZq
NM094bc7eIO2arV2uamAimWfuf4aEYG8qpl70sYESY+tnBHE7w68oJrWj/H4Bpm9CttKS1PLRwen
JBvzymNiN5Z/8irxFIa0wwwmq3v2Rz5sDwW27c5NRRTNqExlBPVLi0FsOEZtHjoKp4dUgEOhas8K
KR1VD0cuUt71Zxn0yN56yjMSQ4li5EBsxJNiTPcSr1uKB9GnPmmatmKKNH2oX+zhrdIlC4m16Do8
ViuvAcExW18mgoe4AYhQubBNKu/6cOQtLlbP/e1UZnp53LPRkvUvXTViPQfBL2EK2WOUAc1Eohvt
AvrTv+1FLXJWzA2bVu5fTXmUjRaLF8mBz6Bm6282rS8GbjTVtdVQJcJDHd9w/4UoB38f4yn231vh
If7kZ/K1stxcSGj4ktuu1x+o5yf38LMQUcUmn6o2pSuMuM/xmI44oB9ZTD4NCfk3W1JpT0cic0fA
TGwu6tzlgLeXr7qzAjf/tUh2AXs9G7dD5nLhtCR6bQwzdAEkM9ctpXiLP0ztBj04dBV+vdrzfbvh
5izJxljDhruAqCqXZ9cOnZvWfxC0m1LNYyGcouRiLJ6JQOnXsLLIfbIsnoG0OpSMcHc3cZA8mDFA
+QxjtWIuqqFRPl2Hd/QDvBJ9VW0/w4zVjdq+ROKq1fxX1KDbBcPkIVs+rcVIJV68EPL4L1MoFNh1
P9lzvcp0LydFuIzG4vtsVRjzqIdNNlTMygOQmKIIufC0ZD2dWVpcRZHIYG2lL3lfjD3FouaW5XaM
+iXFgnVSaU0D9ic/ir2kltk3FvX+y1TxjvsTc7mtULpdPj4oPxmE+c37YAecFSMKNn0mLcmx0gvf
TYu7uELifxQdnHQl2dCVsd4WovYyKMHXLOi2EJhdMjNdJeDYjd3VvKbxXgE+hDftmwnnwaPe0H7T
SEeTX6dGVkhJwoYuhj2r/AV0ytTMXrYRUFuUVqh3Lwo2Km1aKOyFjlXmqGJiwKVF2yYC3+LCrAod
C8qiLtMD4MGqXWYVeX7Qqni92zm4YZPBIoa7dFQ4idT6HyMnyfmmCC6vEwzZn+wW9iT1y1qzB7Xb
eGYIZWSTeX0B9jm1ApWCt2js+ERaY8oSPL9gWLSEcuTWe7lcM1cuKykgwi3W9YS4TEWP/6evfE18
PG5C6bH3T1aINi1hKau5jSZRAK4p39euqvMHwgRguTKJKBv4DkZ06Mcu4BtAHRJEg3IG/TElodrN
rJcsyPC2HezF73fa6D1GKFEhtkDyA4S8jHt0BSd9/CZVA9v25Kzoll25L2F6Uot9mdxTNETQY1pF
c7CeosRLV4f7SEwUPE3o0KNCx7yktbTSiYws2Afyeh6XBf+9wNsui/jla73kXJ13wHeYHoG+DFs+
tbHw9RXRe2K1USNSeFw6j0t1diWG670v0KP4hrRAG/IvQv47VH7M62GhQvOBF9WwAhBflVJpV+4p
TcX3ZlCHlAFEhHhLp76vnJpkPv813BQzSPNnDGpO1ZAkwuVEF494si7o0t8/z3TLxChCFCdlZUAt
b638etQcnwYAaOfYEaNe5Onwh3m6y012AgA7VNcL1bgr1m/r894mKIddTAxlHpROoll2LWdmedOB
tF1OFSXdhg+zOi1QujuqkKsyLYKY5GsnXRFVu8HcoVGPe3wlMhRU7gZlnp252xANKVAdYINuHuep
MAR/7QatTmWPSDU3+zeCcbLKvf+lnpj8j68r0NKYNLUuTfsQm46cJehxz/xXbkd4wieLFs/TZc/Y
2Re/AofDdwJ7o4rsf4D2cGEGEwZ+QAXgwhrqPkivhPw7Db8H+udvv2drnlgr2CEIbYqLBxf3+08j
6Z0qD3+fhqkHLJYx1cwFz/JDE+pWDrLWoShimhq/mVwkOgK4isJ1xNc9uX9Z2ATH4wB+MBrZFkmQ
scTYfuK9FxyOtkMR/0I5YK8PmuZept3uKEGUhVFRa9Dhlxurhg7R4JLirsT1qe5F9ToM5V3dKmfo
X4kJFgyC1rZ2nSABpW6HhtxABTe+FBQZzni2DdPTZ8xKzRH0DJkL7nSJQeQNF20FuR6fVfnoKy40
XjwhmycHDA+1E2/30PMRHknb689E9HQAXBW834D0Cb9Ueo+pmv6BNY5yxGZHfOXeMvkj7qWmpDaJ
ttIp8kI6KJBpnSLaAPFxovp/4L7oBCCg1ZTBjVUPC5JaZFXENDww+qzlYUGVLju8/PVmZbkn479m
cF3CVxk1c7hLUCVJzEQOe2Wh2PdyhW9zPa+8zszk9aw6+Tcl94Z89JUjtyDWeeN55r5NhEwLNNHp
ztHYhWcaUoJJaXQFp6lU1pfbfvoVFC4kqzcsgzNDCmjzisjdrC4Ij2bCZfiRiDSah/xiHjW/+XlG
qFOXqc3tMgdXGRz/rvLtM6GKa5UYeZYPLSD8G2/dFzRj0NW9tx31LS63DTxMhad6Lv3eHybwxD9j
JduNpuOSoFyjCoh/XFmuIhILX5kuPuU++1NIsa+QDHNPG7RRmFt8ZgisvBpX48icivvRpE4UsvV7
1XbcKpuOIlSTaF2BhL84Bos5jO0KHuk5yBGMWx3jY9qz0COXNpEb59kU6UnaJ5YZWdHWQcSe6Cya
s8QIhDLjkWGRuB8Gyk1fqGNl3Y9zl1pibmY5up8n5375uBpVEY69qltgTma5cM3W7tZ6sjedngM0
uIoYVhpfDlNJ1F2x6q80TdFVjJd/OaIBpX7y+3rQZ8J3xJoxZZuGIUNdkyAY9e+QDIOL8S5sc45h
419Ijvlks735C1GKuns0Eb5mc64AS2b0K6v2i+ZQFftn9VBznMFrnboYucSNIuFQ7SoD4wDvl+2Q
c5ZQA4zs+jb0AgFeI9jBlHz1Xx89uKcKiW9C+bv0zVFhoJoKdpG5e6w+DMvvkP4kDra6mGXoPSo1
KOTBnUSZdC155/UaCK6TQKI0ZA/1/cuMyWuJ/rJKtswM8N8uZI9dP0puk5LDGgelPRRdAzTlQ8gb
SMnaLC+ZYSWee5ZMhEWzv2TFBZ1zGPBJvtIlYT1CzhBnXSPxSV/ei+zjHHoNDV79A8kYCATOuDYA
N0d7xMbnM9duRZZsQdrR3MU+tnQ+muctGYp/EFC2qLg+1vDS/2JiHsQXvPPW1CbYdh7GG7VZLyrK
KOrTQ6q+Gc4++vrdiA6PwXvifmkALdKhXmDqIQJZsIpm/T79rdOlLUB6NfTyQEoOS2mV9EDbS6CU
xCABpzM0YtP9GzW4fd6TqOf5AVagJznbv527Ped0OjhJh/DxmeFae7Ui0FRl8lWK/adjZCgYF2jU
0gVHhryoPWopWQmq6kGjmcb6DK8DLwWBiKh9h82B952/A3mhKOVE7bLjZ2jPxzVIklk14M2yl9HL
YhJU5Cdw/NmhWqLc5tVy5IFHE0WwZmtOHZWJkhn+o2afuVPwXE/+ryjsFcA0Qqfwpcb6cILUsjbi
IvhXnsu4g3Vb8hqF9y+MM3VwadDJHOdI5gWqHDZov+IYvKuDdNNCdpAw0rjy2WlUyG37Y7+h6YOV
EVpFZfKCrB6N5YbYLvtiosSXvIMMoE0lFFnse73DIKU8inyOsm6yD9L1RysN75SyYyVqM9eQS/YH
R45y+PnZQGS3xHV2ThsBM4w1w1JrFr0T45meGouSxll6lPIS5n9NjtaRYVFbslo5+4Z+iiy2uXIj
5oLq/YUPzPZDrXOs5P3e0KfvPbj7hTo1KfybsLCXiYmL8usMFctAft6JiuJLF40SuQu9IaVjjPLg
dD+7KhVVpXgNNDBMyqKsxzug38gATS0OvW/4q8QBmHqOljIUHZc3nmUMakWD+UrCEOBNOywIf+Ys
/4vubFtsocRRWSPqdu+10A+QniDEAuBCWDixDnO7YEkyMtmdaRKhrQaD65fHDsRrODCqoriCutzx
+DN3YmKlD+8YWTJ56U74c5iwNW6VaFcE/959vTKHzKqVsrmFvNqDwUUH4lGKDhpP4BDdgshTa2km
2XHJ5vXTdixgHDcrINqmnFKhjmqrJEqMVyevytF9MLeL/GxOZfz6hWnxUAA50qTOnRxAeQTx/TW0
OFjBC3xzE+WJofEQMYZtxtPQ64nPzzWuIyb+VsuWoG+hNri+qmJSsGXudz2XIIlO0jrkf/MTbjmr
JOscrjFUUjMYRYJtS9j3Hek22xm5CmhwKr3p0dcTa2TMeRJmJyl/YMrf3ff+VW0PvssFWmzddnLs
p2cy1RQMVU4HAc1/TgWiaIAkaczUlTuTod4z5FuuBO+fvgbVixYCxnxMASIKEIXzYXeZAhkUw35F
VBGTURKadWXjh67BOOc5JY4d6oNJy2QjcisdgZ/SdR0HBtF/qCjQ/DkcHm2qxUwl18Tm+s53+qTs
Toyr68aR0lz6U+dr9VO0SNuGMFRqWDcmQrGIATaofczYtU+Yw68AISV0h6OHerrTs6dfNwr2dJUY
0aiFBib+CCUXyabqlQ1lYfZo/+1+tU1ZWjAU1WSGXqxBY9U5DQZlOA+PYbiJEi5snhsLF/7hJnax
EjWCgzB++xR2k41lJ7rGKzB95gB/Y7FUscR0ncED1fuAWQhzXSZEWbtDcH1W1JFhberDGICEyDlw
qp/S5ojYh74ut00wuPP2mD/QMHZyLtIKvZhe1q677RCxBYiSZ7O0x1/tc9LexV4Ne0Dlj71j01K2
2Lz6ETFKRv/fNVK870Adr6HlfSO5bvYiNrgqADYpnJdYBNfrmiDOCtmoi/iT5fNaBJhWHNE1ZotC
3cPX53sktcWRNwh9uhHLw3Pa0Et93UkCCnu2mauNclHBNAsSZaLgHGVtgvJ7higoKD+OitjMR+IY
MI+lXkPfAOFsoienYEKMIsB6kEDjRhf2T2HVK01XjMJgFqkvckVey+kljuAUJkyritOfq3Kn3UiE
Azwuh39bjqJMke2g8r9qOM92OuICsxNWvFTwVcxisRRe4DnSCqVw5RQJJFhO+9WConMqKN0UzX0D
yxIDkwNLzW00gKkTUtIKycStOyzSdTqW07wlNLzM2w6sqCTUPGm+H1yk+F9l7Q/NCUb0X3w5dZT4
7hPzhMIjDEQTJtRy5OYCPIAwCwt2sF7EL4BoOEc+/0W5TXtHjB/EQR1/G5yA+0Gwk+YAPu6W9S2m
eQ4fimJVqiYIltnwPqoWTadojjN375L3ZqcmwiLggnYTPkU7cEbZ3d4U6GE7owwBZuPa196l3fO+
WbtihqaGdiHv2HIAs1gY3FsDSCa0UiZnAAGOUKBB8oj6lzG2IX2D6Wq9n1PVPkUKXNTxOQOGpaSz
kH1jiAEFzSCzQ2yQzG50o4ZH4orA8GQXslPyK77Um3L0oLXy3Ch1Rb46N+B9B6LUy0NF3ujOo5es
iaQ36nHz49gHjdJCOBV14OXRvSvakYYKK8kvDN6AmBHNbvg2/o+4Oh3m8JMaBLwFF1MHBnqVza/H
mUGpqwgxfE1zbLov4HAq9f2WuYst7vYd/xn6omljNzVu1vHImpoYUHtvkm65S7BX6yUaRsKmcxKP
3Xz6CFkAfE7btx2Q0z0W5N5F8pjePXekNkOFXOfQyWLhkqzybiSdg7TlUUNurNrdZlOmKuxiGq/1
9M3jbq+mX7diT2sKuf8z9l8VgZ7IV9EfhNHfY+jMVNO7a3G4EcUHE7fyP/xdAQ5wvKo7kHn3C5Ow
ZbpjEA36Vc22Zp6tGI0w2P0qIzxFmLBj9k8C3Qu85VHtB0gEwEqMz7wH6+mN9R4BYCZil9eK+Q9r
UnfFBzgG98Bv5Iwwh2Krnx39Igz4tgveCKZEc47on16ztn5L02TAvjIUDgladeZRvM9mZV+kWr41
XZeAVAUgbFtw3F9+s19xQBDdtplBphaS2t9aQvwsDaqUrAfpo32D9+71GjvMl4ZlnjWGWYUIa4gS
wRmE8kxtlPXK00u0VD66faZvXYOGA7F41R+MIMuXwYNa78l3lYlgWOjSIYsFILwfK5iTQ+INi43r
fDWkzp4GD65Qz5P5nXR//0H6bpvZvD+hWtXzfWks0iB+5nRR3RJQJ/+kLNcvcnJwvb4n+IUMXRyM
h8ALABK8+B20bzso6JqkxhVsQZAGoGEn7ufQ5QwnPDA1o4+jRYCQqh17R+jd8B5f9dlm2EGNToAP
GB3m64rQoQbI9it/5TC53LjOf9LapADuEFvtGzfD2CBiNUxGD07FkGwEbcFYr0xwvCJzocu+3LNY
V1fJbPH5x4qpH3c35BXjIHf+HCEaCG3CzENOSKU2LaPKf4YFRXAIM3MXtBthtah5MjVji7iukOcR
yHAtUZPkaGfRWLQnQ1qQuyTB3c8SMYJ6911a/77wQAZZBCpH5Ts09C9oj7X0XYEJXlJIZm5sd6O0
e028OGzqS3rCxOySHGR/vMhw5ON33hwOvxgDPz73ybvj8AROQoiSDWlNGhmPR+v9Qqmz7vaJzZJ/
GHACP1IA3Ht+m6tN4U3UycOPu2Sd0dlabstTvDJG4DYybhYR01J5C6P8eaovub3lIY4QO+IYdi/b
jthg+yjCHc6c33xbtsd2XXza1lE6fk64xb5Ayjio+tRmeK9EOVm28XZKa/jHeysMFWEP3w95R9o+
bNEuXAfeEb1vLztjDSDosyNR
`protect end_protected
