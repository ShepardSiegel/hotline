`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jwlxV/vkCTFGZG8dKLBNMu5G1FUPnQLS1zaSJk7wvWu7+nCWZwt1UFMJhcDJxklXlbkT5c5jqN88
xTnBy5kJuA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EDqU3nOUWK4I49qYMiw+BQ3Xw6+d30y/7EWRWXO84WJClvjjVnfJGKLePrlsi7wFDrMdaNtgZkrT
X7FJHM7K+L+r87zHzR6IqkODI6+I/mP/d9gx1xhwgtQ8rykAdYWkdZoDB9VTjilMgIEUH9a7Liyn
YGQXj9yCLztnc3kGasc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Aw8BBea9gPI6Gh8WZ0GiGVI/OzA9BeJHTGTso3N3uvMt0w764EIiDYzWa7RPqww5R0+WVTq+UIhT
nzQBr3upIxSswFx/es+hsHUDuEqLHbFq76fFtvphLDZvWMjbCYELVF6fZXoi4auOUluZZrG3yz3C
jy5m7GrWGcNLIomy8yF53OXfqVtWy07lRyz8RTGeWnQrC/0BSQkUDecZ7gdzFW/FukXvFMB9LStM
M06NpPTE/cixi4RJAYAaVZYNcmJhJk+kUKHNVuwUSHZ+TUBJ5RChm61+Pf3a+X1glrXqxX7TPlKm
qdrgz2vqPpyQY3HciC446yzr2hGhrBBlNMEDTw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PY/CnUxO9QvbGaOzmqzQs+kLxye8Rs5DUwWCfSTA3+5vG+r3K89TENj86w8UgIN9tA7srFGSD/l2
vaenjaisHVBHiKhukE+ehtHluXvpOiVyfZXahGBQJBVnyyw+wsPPrVS2zl5xfZ9Z9d5ZfIofOuLE
1sgwwF9X4gOampxBU1s=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZjMCin4BY5adx6qAtkTk+OfLU1gltpDByQjADLAl7XwnDfK9pca5dhZikTow/WfrIsH71pd9jN33
jipA77ulIh/NCd03HqcWp6gVVySicicAkbu/4bV6f050V8f5uIi8X4gakznPJEt+TFt2BN2JY+k+
IBhit6OLLeygnNOvGm9nLnWBJ73sHZM9F2koCfu3z0mwoBkiBOBYPggrWyx2Mv7sN/Cujv193I6W
J5btkUmG71BKnPq9DIhhUWDheuGifFOF7Pwd7kexRpeYd75QYTIDagI253uQV+BwW/puGemg32RP
fRe9crRZe9ckqN/h+3NDEQNjY7FH38LIfTPhZg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7264)
`protect data_block
1ChTziMjcCREJGxZ0gBSKWdkzLA3zGL68HW4CGse2OKCg09Md+JRyM6dkk5FeMFK1LPhxkpPnvCp
+AhdNrcbUjErZru/kgifPLeKfr6KJkDimBk3NHPg2YDp80O82i0u0omav5f0HcaUeI1ii/eTzAkT
60U2KnWBS3KfKEFAQPuE2jdqEED7FMt+ngNPjsDj06Pwylqei7sAYhUe86mkm0AD9INzmFObsmiI
plysHpAER5//z+vOibpEIfQlOZHfAna9uhmMVhLnhaiMT0FqWFuIT4jT48xzFujUrMloFqzUhfO0
Wy5h3D1s0Cd08HkLyakVSRbZS5cjT/oqzfWV+Yvbduw/3SbIJfFBi2SYJ5ZyW/WAJATlwJie0hiI
tOY0r5VAECh4oo3BIDYmqUGOmwl8c7W++mBPLfYQRMpR17kxiF/IXBzU98lhtZ8/9vAz3EQYhick
4wMdpcZGY3ydsfm5J8uLZr+Tn//Xwcw6kne5VF6AVVM1u/Qd+KOWu4mSeaEkGnyznbfImnFwn2DS
0NjCPPmFfaUBJ6QtRtJDQLVwmWKT3fQvyA+k0PLEjhN/yUjlMXpoRh38cltpTzl25iTZcFiVeGHd
WjK29s2x3poKoPEWTbXwOFvZ7Gj0dlGClTI03p4ZnfJn7ZDScCIpExj+bDZPfjZr2W00kp/wUNvG
yGxmxdB4MvMyTN8JxK59kTmxAiZyUxVH1I3kPfoRVcV0+mfxMXTlvgw6t2AZUoXbq54RMP1NZePk
5zl8e617aZy7p9QtrJf5Mo1DA4JSWTfjQhBIqOs9fBCm8AG9NOkuksloAOg6fkKjW7MGNzUUNtdP
hSvcOmRV3AK/bvpLG/DVrTiKzdd9R0Kqps3Jh3ekDin0g6tbnaw5zZ5mpNN57/pwIkoh5BfwuiV7
S5I6G+u8G1KbFqB4zy5UrchTrfxwqHUZfafST1PQFHENfVqcXcUOYgpLaQXQUcJulu3fsFAg3bMl
RGZE/CttsVWoK85GGEOMOEPxQ+A/RDMo7S7jeNKV2x/DALQ1HxXrMhOQte6DLBZ+STDaNEDbTd//
+kTETkzRZ0zzUhiFouNpxXpRn3EF/YBdNU/LGUZHnRA9NlzfRVQRJq+PRngQ++yuzUpjJTJ1z9EL
KoS5rb5XCDEWFHTMaNSMeT3QeGnuynFa4YSMgWhUxOkx2HE9zaHvImJFDRLZV2crA1bh8rAYPhI2
luXm3Cz4mQKiQJFN1DmQehtVupjdKMPTOlgeq/ufkMg5OZV41xDokj3FodT2M5lApV+/Q7+//3S5
EE4s8VW0FRVDTEWUrFNJlAi6lsgZqY4aEeFNkYcPXSR55UFDH0QH9neMqH1sGPpcF3itldEFjUCQ
aDg/OM7d1LsRnSPN+ICS55c6pRMEpLGv3ZpfluIzgvx+TLkcdD0knW1MZn62a73LY2ttxHjZT+aV
tf8K6dhjVLQofuolMYGLUXNSVDuavxrDOubsd/B7Hcp7QEiHLFlg/HM/9LuUwNLZdN2bY9QkLjzO
tr2g8kQTF1SUVRRwHJr2mTxdsKEtuX7nSsquaFi7VORhTqOOhZw56jUhxKbC95L1OjOvxIIsq7+C
7wxf9Ju1GLXCzWtrnteVyoG1mgu7v724GPG9CP16y6j+M+D8v+fstEFvpWprpABayeQ+Z/pYp4GJ
Q/wl8vSWyDIoI+crJxP3BolTMD/O+Y6tsKwZ2HAC9MEnCcDfydqooQWzqfy1/OuL5z/ojUq6pSYb
RJx5NJdI+UEOgIS9ECKoUByzJ97W4iU5cIeTSKNp500z4TLu7/6zBdkWZrABVhzV7gJM+wulP5Ql
6lBAoNHNWOPq5s418rl6kccCHUboG40yzhVeZDjC3nd3X++kVBRtIZk57Cep1yvnehC6xZhqBEAd
OVqgtl3aAf0cV4tXgc605+6ZOo0HKZkZyIz5APfWgH9e7abJL5hvdQyo6Xyh1TKAkVVW56So27hv
v4y8C9MKM1x/v8fMezJom2qQOJiac1IH/uarwN1yJ56q1MizZZO+TDM0XvFa1U4Mn+C3nY/xDG2G
n7ThopdBvR1MiO5xrTYCFdAuRZSDs42yoVsqgCYDyqA1JEJ3yYsaRgT0Zu4TCR6171zj+fcKYd8V
+sfDJJiLmEIAy52SrTDx5IZ9EXaxW+AEscnB3LTSMkcJkPO0d7PYaQg6LlXRftzqIvZfDEj9CzOV
zLfVhStOf9/pTRsJYHxI2V1YWi8tzqk1kRj1y4dN/FNdH8fMaz9+FS8mGyIrSkINHYc8uxumfs0j
o+rthWrtSeFLzgwND2P9B7dABHZ5E5ZrYTnEwmueotAUANRhlYaxvm4zTJDwMab8awnm1Sgt5PqI
esEDQEh2+bUwHNGOPTVE3isDYqPzV5OGDPlxpwXbQtcqpmAXJ688Rz+149fzt+dhk0yty7Oz7rPa
zy1uICsipFhVDmyGggPgz1tQxsk8ENXRYsgEhBxMbImhsx0Tl3PeHyPnYVYgEEIwbH1ZnYTsy0ci
XdlHHNunt1Wf0t2Cudr5vi3YC1g3PrxF86LA7F+WDrZNFY+PADMPr0MHIYJ+Xo83RDNVOBzFU+Bk
YToejMN9g3zo9LkHLqVgKmfHoP6GRJoCIdomSLIHsFCMuuVwb2VYV0XhTpD5e+aSRzDLgRU4CKLa
ddNp6sOlrh2axCeIYzzj1Pa1AnixVVDmg8vMN53QhkubtfDo7fjhGnz6AY1310pmNC+19p2zP4LX
vLcC1Vmu/kzLMeoK01RfbYezpOOrcsn4NuDrgx8etsXUa2v0rioys34u0g7LBSQzWDfs2xY9NE2G
KHAZ2nNCia2+q9FCbse7p1zFYjB3z3SFH78yepuKusMWLRrdPgOkntPXYnqn/qUuZsXWvmCz7d4K
MMRcw7G1wzVmwY0XRMh/VgcrMX3vbdzBcmYEfkpfbgJuV7m1dFnbO5goC3YFwc5yz3N51W9kJv/S
ENcrxr8dhoez4dGonwz4fJTU9eybD6jXKz7zCQXsDp6qDZbM7kvfk+GjpqpK0zdiDjOC1kvwzcbN
JObE9h5pcE4svBEKZfnPmgoujIJj2A3ygGe5p8BbSQQ73ozC6sZM1INRaWOZeZEC5ZjBIw37WNb+
iUDOW+KPD3AWJrx16KgHRoT+dtebyJpucmMrNTehXohk2JgZj0lLml+grGz+YRB2VTILavC29EMq
Fi0e61Jp3yVQF6GWO71z6GSX8LvVm55Z4Q/ybT/i7I15a847T/F2YSgqcneoh1preAydkVUSUN8S
YQOQnTr2IctClMaAHPXCfeVoRdzjwKRvmktmy7wZwelAcPjU61h6iyjLyjmBJispyHda+1j0bwN0
tYB+9NUltgViygL195R1QhftsDmLaLfLxDfjwtShc2mo+n2dgnLj9vBHD5X4raBbQ380MNy1Rzf+
jw1F+3Xi00hQ0vII+p4RdIIIm/bwVuut3x5C2tHhLkT2X9gznmC5hHE0KEoxtSWwys3jv9fT+KHW
cTIYBZxXxkm92SOq9z80N2POCWsh9/1nEsfeDvzbtmvb7OR88DmSiQz9iv13Q/kBm5OEFNJRBXJU
dVbV0sreXhrKPiF6cp3sP4/cWhuw4LwqJU8pI2GmcZDjx2kZ3dEE/F/QXS+72luJH+tWdGg2FCah
mmx+1clvifPzhKC94ATahdosDVA1pbBuV+Z1k02o8/wkWF70/v7MGTGkUWiF/gsIgv+/XuTVEQqD
9kO4Z56tMKZsIj7OfVt7UJYHxdBCtEe3E4sOsYEHB1z6gzQs3ZE6MVbshXsHVRHGLqbEltDDTxZU
nflGgaNBE11XLS6XPNoi0QDVqel0E+os1e1teqCo8ckN+QENKwTPF6GnNL922eqspVKkQjV/ob14
4gvNT7yliugTWaLt+UZWIrydfztW+rvZfTXdwhmAQPuHlYDfsEX3QSZyi+ewm+U1fMwI6uiY7SEx
dX+vbVONgYm1qYd3TMCrwLrpjuCZomxXsFNPbZpIu8+WzHjRLNKGdDg0RONSSOmIWnHlMIc3mAb5
zi9TAAdC0RqF2yN00rQCPHrdAYD4zZ+Kr6feWWyp30X/vmc5KTSSa/ZQdYyXUhPYI22FZq1s+snd
awP7CB4sfxp763UJ88Mn80XbR3hYPx65W4SRtsEtZwNzZy9LpMZVwOMMoyX89P80ImDsK4dYRFLo
9KvrGuqxGKWflgVsiOvW5feaaOxu1LNWhlTkskjX9d7uzElTR82LBrCn8rg+naLhJidOnZt33P0U
S6axGsSgRiNFJWtS6SJWVT9rf8y117dp51szP+jqiD/snWnVwRaO/tpvtQTwWRK9gFuwzreQ9azW
n8VZKN94LRd/xE61y9goovmG2loOTlGBsiKyu/nrC8D1NlmWYHvZllQlnWLC0Mydude2unKy2eLA
NV2zRRV2E6ospG5ADwZm1ngxfEuxIZMoCNXF7gmMZi/K/RcD9xpwa6CkDalsC9cJ0+JlL0lL9znv
5ruPnkWeZZizVK0uahAEU/zY3W8D5IP66vPKWWupoEuGnjd5j/f9YN2CTVPA9FdKZqMTjSJ6ZGsg
yB8hkSNTKctfpRIxvV1alyfQHislbxMdKKnjQ739/uGtSg/x5mXx3YJHhC4I6liYYmO6Hge2rEu8
1AjiR4u0/kcIgi8BhHoligChCSsCVF0mj8opFDFNgRLa6HuzlZurlFPEzEHTMwepzJShWZMsE6J8
NMyVG2oHFpPN2Himwlv76WdVhz/kAWFQFpxbBInHsEQJVnmHQ2vvB+nLeZiYZ2sA7WfGRogCd6xN
Ww3YBrCnoxkt1eFrKbL1qt/RTIZ8QxRPEStGsTCujcecBF+v0kZLAIs/oks3JwbSXs5b5Yn+/CIT
e6EMsSRPKiqTju1H0rl/NsvJLqYOq5MnqDrTl51n4MEBSrMxzsaD7TeDog6ElxTQNN0KaPJXJXr2
+wcJqVtyMQVTtJSMvtzBzyMAzXUvLy5gvB/Cgq079o9Nic/0XjhwAMpJiy4ET7MT/QcBMzYtxEzJ
09WXugNOtxE1i3O5b5R50zqhnd80P9M6vIBdRYzsuM5URq7JK0CL/qEAzTzZ14Qt/j5pEltJRFfG
C8siQWsJnPD2MEB5hLyfY+WNjBcHdNh4eGDTgfBPvT65U16vYpAO+PiP8yKWtDD6XhJD6xfUpYMC
7OBLbrl3h78tmq7ckrhgT+R9OVXcOaMX91ZMzdMYpDhv2hB6cA6hmxuHasEesSU4jzrnFLexDOAi
E9J7A2f9eioQy6nV2AwOCPL/TYzkxSlEpD/Ua0PR1BQOXcF+NOo2C1Wu1xhQaha1nqRaztfW4zVs
xsw8NDOG6a/IpcP1PrykwrAqLEk5ByAfNNnxqSNLNh7JodjsB5bQDuibMTZuso+2rN1dQGGAFcGr
Wgd7vc1o3Z1HWh9JIHOwUu1yRuDe7Ogpg/zR2pTJsHEUnjXM/s92sZt4i+yWbiGNsIpxY+Iw4S2S
DxoLKnk6UVUe3MhG24pE6D/bsjCL92M4lxpXXvMdiJARWTQ1nJFEcBkqT66qrIEf8EIrV2j/iYrK
i33scSkb3zQ596HbcfaV647svhmBnMCWtW+RCsUzSu1inJuCHaa2AOEh2ed3xo9ENjyzZHAltWUd
fbRgeVaYKHBETjH8i3kFv3vFxUvZXMAShWXVBrKCTaRlIWp0ZPWcb605TivkkP4GFpLyypq0BY6t
3oDmDTGVikiVmzhOC3C17sP/3MoB0KMTiaBekEvorEvsKZGhP9SsV+SGpfakSF8FlZAJgc36OV77
NU7Lz4cI905NLWImrG59qYZhuogmlumVnRPLp1IHNUEV9USY1ThuNUJvHqAHPD8wWgWdiKiaSR7m
oBlF2ypMCVuwVIdWqr5FYaGyU+4YZGZgr+ihLIM1q5xfuzyhxJUOd9giCUqJMdqEM9fFZMcnRNUz
JBImoDKxeO7pBeaFewmb/kdMO5zgCb+I+JX8S2H5TkmG36cBpUeaLetqlPaWVMr+FQubfdCJnSgm
9LYrHZouvb+vAqic5REgtY/Gaswmotp8YvNQ/YAxOe6oCGCPOs2jsBBzIpyFta83V9NJk3A3Z6Fe
nBsB3QvSWCYhLDijq8M3ww5R7j+x0Cxba7ThFiPbYUAevBz8UMnDgpCVSb5ihTC5nn207Hxpg3n/
R9STpnRC5kWKD0LfUvRH/tfsXJvc+Zu7fyHJStXH89J6+TkAm6v4jiWSsEDQqwpedtNJLj16NK1N
KwBHm20V5Hx4focP/W0jC93FrOMKJ8MjbPz9gOSnzIxHlJVNU2OYQzC8gyx9KUeqj4RiK+V1MTuU
JyEj/OlC9w2K8+BFLx3uAV+HYFPxpo5LPDOSS90ZAtnfBtLHD+WFY5kaurEkV0juqSxYr6rlDKFW
5Kc1idLkElvO4UdcT5WhpqW4t482WnGIXYseWaNYFOIWsHDcAYmrgbO37GYcjzfHO+BfyQUOVxk7
Ce9smwGcKndVihPWZIPUGI/U4JV4hRZ5O/n0eJHQz9/tZPYxnC9uMOull8UILoBmfFw+/OqLIfNg
xUCUGnqeZzckERft7SA+9liAqt16zcqw6p1B/kvdsv5RzXvqshqHRYjiU+Zr0a6R+MFOQ9fHk/eu
BrjE2qvqOCy0InQ7kQpM4f3bzC5iaHmSHxJQO4V9uN2oEZeipBsRkgP+GyBfvTatQ2+H3nTOLCkc
niZL84EHwnRjJ4KopK6kF7tC6+pkP5/vIGaQN+f/0rT5tz+dhV1dmQOShr0Gfm+mGL7YoKa6x/e1
HX0pvNshzE2kKCt99ORVaXKfM+cBhBJs544j28Q+CRGYQNUg0sOGqGp0cnukKRPkW+v2cjSBLxjM
rqSuOUYV4Oxfa4MOLHsXKP1uAkoShWsWLVpJCPQxVGviLs9LEP41YJC2BJnkRMgdVesOYZP2XX+V
1iYSgWeoO62JpXc1tbmzE6pq1aJSbe8NsqQVDFThzJzxDBwYwTwkVMNoLxVmSkwwvknGOxNuV58f
U7daXfd1+4USHQzqtisJRZGjALPl/WYblCpMjpEaFoyJuU5GTbgrg2pCewiSGuOY4KfxRlW8OquA
sgreptL6Y+3NlLcDb0z52J1DeDW7XMlMSQEWCfu91uWtvyL5U+Ct0IF+PrdTaDBATmmudpulLQXk
SPpShuQhsDY6SNQzrrK9pXad/TnX1fO7nhw7Qbsjxuz0KoS4ijxDXfk56q98cQuEIYyEvSfx4K8/
razHCbegHxwGXFWBz8aA7PfDW8OjNS5SyDhbXc5gxAnISi3uX5SaFoJ596rsSQBxN3lXFRKabK0g
rUfbmkFvtz1oK9AA2j/GDl7B8PZjNK8YLnP6NsBrVmTYGEM3v6nMViw3n+dPI77wgjP0nn36k5x9
qOhuhzI/MPfg3hAw7P869w+twzZQ2fUhAxhoM+ohCl13iHhQ4/YcpU7s4WP0Lej8Glk600C5J4up
fyx7XX6wsXFfZHv5JPXd160CcQCqgwaa2MfpnxMymYq1H7M2pxzx0UMyUML5jdm6AxRfMNQok+tp
0rF09Hyh+ppiKPTRGf0Jfr7GYkBWatDRoaVyt/B9zLWhuz+qtFjKzCmeRUoWgnuwFzd/A/VOLaNI
2Gea1h/LUcGc0dyalgURS1+CWjh+gFyuRnom9SY97SBFR2ILfjGRtT6H01XG4etXSIG9HbrBprmP
WVPKFaMUXR8qXbe3aD6v9IGzp3HXOUJIhmlA7bnZouw1dHrq9HHrUf7DtxgLfAAzQtpZZUVPtXYV
ERmEx/v5ob2hn3/6hQ8NFRczR7fiobCP5Cbrjnj2IRaBrdAdjr9h2GbnrTPVGYLvJ6JR5e3RupBF
jmM/oGuOVjt30ZQVk/mjF99AUJxxrS+NQVWwbVI3rNOaLC92oRx/V7P+TSU+yytP2FiU/gmjrpM5
mWFnDtljMe0Dbkswr7ekJNm5LFZ2tqtD5J3vJf2DrvHnSGo03NZVavMaqiVUjivnrxqk4J8QmlvT
Db+GQvyswnJ4Gq0Z5mvm/IfKl2b+dCMErhpT1OoJjW5aNitEODb5Bv8qYBNwfnJMUZYZWS/ZIDyf
EyIXYBhHoE8aq9cwjI1wdyfp6tLSVjT0nuvb0onv6sujh+dy0bpJ1Jb9HE88+noNp6vJamG3S6Q0
TsxG+M4dY3YUxC5fUTDO/wAACiaFDKlQ1hLcEA8EAf1LR6D4MXRVFxZLBa0fumI7H65gZlNXBVuA
1u6Par4DmgOENUlE29lKcZ6X4+FzbkQL48ME1JPiGoOiib1v07R420isYALMw7zc6/5unXfTTEAQ
MV+H/pY8HAAnatiNSEsJq6kT17zb6ZGi6x++PlVaU7jpQef+/ygkBasXlxUCcDNbzqB7kVxfATEB
ckodGo00lm6cANJerYXlYpRQeqQz02gMsgP+paHhQUiuxB/gXsVYnMA3g7VJL4pM2abCG+f9I/RK
FCxj4sb4MrJl58gAdfLZF+dH7glh+Sr0EWkufF4Qfitv4pYCOfh3zZ6GrBXmBap6MjTOUlTNGadh
dDivUzIkAQ8iDV3fPWMhJkIEY8SDMMxYYGPA5YBv5fUZeBRxYwmH5N989zkv9GBvpU9wMIb2kFql
PBtEo8MhFdry9DC2khYGU6gD5OKVyLj61EgkYa4k6e15y0hGNH8/HxrO9H1/vH04B7UQ0sdhvSUN
QxaE2q3wGg9OXTAnI/P6sFv3eVT3LzE4ZSPcGVYZCP4A0SxnuYxvvESCO0ZxEWFSH5kzLrEqU0gB
8UKjQ74XU9zR7M0dnCbhw8lceuAeE2T25agv1CfObbho7AIW3Lm2KpYv8rqrzj/QbpSlbCz5lsxY
rRdjjoxZZJ1SpDVOse69ShH8uGAEqck5JvAb43v6/FQmzZgBnLcLLo84J3TWG3DmjmxG08OGBr0t
KhKJfWFcPT8an6SPwaGJz2r4PnuRreSXs6omlYFCAjF9ODUffckdQGpcdWTC7tOB7wKKtTScDFwB
9xy+zoX5C/1tGdY9fgkAI62TwA4+4AfAjmdT+s1TUByUbNuoI0oAHZvnMgd3RqKs2sC8PMFwbf3E
awGOX/p1GDzMWXn7lstB81vtyBpAxFXw1hq7KCewsJdQQgWfSxq9sp0gWCgFM+ztN1goUJIM07je
c+5Cc+HWDnRbDPAQ3uCDKyXMEaFnzoYtTrUzm4Ta3CfnJGitV7WFzpLW6cxZxuY8MiQF0WpUk1Y6
LA4lx5Z2su/NHTUV87WTTNVNhjdFP2Lp7GV8ncZgBZRXxdEh0AxbuDav+vgzgU54HMZr+h8W0z5z
eP57qxYysggMUZNfOLD0N51np3uNf/tdOrV4omQskrrokwLpjxaNyfugAgSKqCPezI5GsJQD0zdZ
Pg8M+HOYahIPuNae4Z/evlQlWwF+IGyYdwdzduy67Xttg66x3EvmxYwBCwSzv71cXwlPY7pXLaQS
yFu+kJitInRP2K12BAZxFLaenXMC+OFfxjqGYevF7eWDoHmzNbRM4UgqtiD1kQN6Js5uuSCl47Qc
rhj7+Wd6NH3BhansoEZcJv2meydM7aQDvLXgLZvq9QI0wV4UqZGmfGSWIkXbOIIItCF6++aqnWlv
ukhFTH012gtr5D4tKMNVjkEvlJG77sK2EV+xt/fk58jcoCAI5EIVw5nuyd31dKjeIqRnlpEGq2n4
CPMC4Y0S3vYdd5M6PMV++X2nqok+m5Enng==
`protect end_protected
