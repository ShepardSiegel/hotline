`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
l/8kmju7qk/MO3B4fc4fotFQW2pwxQxkmZRO/caP8sTUV+NA7/h8/6qoVuS61etF7fT9rWN6X/Tl
GLZLSIW57g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
arcFEzw+bUi1enX3KUulNQct4QUGD8gjgiYiHF7ZBW5MUU9QzArMDQ0hkrZEUzJ+hMP7b+FF15h/
c/x3NGDqpJcxMJMeCmozYb27Dg29IzozdRdzG/L9q+xW9NHOkTqEv3RhVjksZNWb4nNFZUBFcFgK
vGyH+KpQqVFFnkADMuw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dcV8qXGvjRHOFWGPBs2hMLajhBH36sZVOju79gorZoHeB2pLt4/wcPwkLxT7C51qx5KR/QX7wQ8p
XJNQhLgQY7p+B3XLKMUV1gqYNxB0IXTxcoVPsFDaAWemxPjujp8YwMVyfB7mn6qb6rEKtPHDW8Ab
rOLRKLukgqnmPFT07CNUEBqEkRCUvtk23jO28JCSL64aKhaLJer6EdSotK3bmiDmvos7JpgRDEmA
3cSPEqsiRM8LKDGkk7BEfMpeyd4oYfYp7PfYmHEFtPvQ+Ssv9mpyOHIjeP/3j6Rd9SF6d5tmxUEb
vPXL9Ea+1EpOs2hZlUop5BOFJJqFnLRyiqZYiQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
I202mPV5zh9XPeJ7qQP82XfAaAr9pxpIMgecsBebRK/T9vMCmmKybMGs97naLgok4L1hi0l8K01t
N7UF5ZJTDh5i89mUcDgVxjbz9XdfhYYHS4iN+vQeaZmNcCQz+LO+ZGobpaWBpQEXN6gxlMTQzBoh
zHDiNvAHpfO3TLxJKg4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GKpR2NZEz7m7JWKX5FRFYEzTRYy/tFUaPl3IYndDvyS6f5Rgt9FpuF8l608voPx1EDNLuYCbPe9D
EqY6W/HeKHVPAdycHBFgyabcW/UL64ONeNtfBxbhaUDSkqlKv8TMoHn9UKz77kqMu5Ay/mXy7zDJ
Xegsb37yTHYWASrix7KTdgWhXl2PwFJtjZQpLFFIcbdFvKSfGYx0zU3Q269QQdu/sN595MkDMYIu
72AJ8s59GqS72zQOM2wB4iOfLfjxfFjo11PgRsTqgp1r7D69bX7GRJ2cnBJ/yUpVveRKYMzrbyhG
nHQ7IcqUu8gaGJzDx9sytd9qTMIt8o8Xvshk1Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18240)
`protect data_block
K35Fbc+jjIGTNGIHG8cYglizfkCg00YLG2qmOfe504WWimlFEs5Zx3XoowFIo6LrZ77Ka+v5u7kl
XD10dR4QGpSvygC8tLeRhU6N37kHSuT1W2lS/AX5mjXSyql0SgBbIPniCTwsOoFNKAgEG6Iy+jh8
taNVwUbnIbWQ3ATkLrQ6vY+B/rnArRzQeP9Ps3wbiA94YBC9F3htj5uHTJRuUi5qbTRfR7ozF5vN
OTgwKotCaDU4rInCLuPgX5VZHcFycR67otmccfYp066ljsXZ3wE/3PEmcCcWcGEVMyq2w0qoH6Yo
NiFIIi49XOfk4+8YTEqL+KRPbR+GlTpxphO6JgcHTLz2NG7vGnjHpxf9mhLbMw6K8C4693u4HUlA
94VvWWcYGq5337i4UmyTN5ijEe5eBSbWvsLatLC4FN3Tpfhc6bivBzxk5H10zqF8DvZPensd5Tz4
n+CklFEglsMInEGYlrkGSs7xFcSdV5azRdxWhgsN2FqlyJC9O5jiyqKCGDe2D90JBpNIp9RkgvLb
9qwFLosvLwrwzHrUOlz3I1qdgmlp+mzoWbuTLpKoOGihwwqjPqS2bU0Fx5lYUBh8wUimSMaDsAgQ
cC65zBqV9pQ/cNjlEC+VQDTuXJWHDlqr1wDd1ruQ4bSGZeYutAQQCGlsDS5T7r6LCr9f9J1cIy6d
New2xq4kXe8gAv/dflgkvntDWlyuGVVfs+p/l/85oHsR6QQOVDul0FOJNiy1g1Ahk0hEgypvXjVh
TpYRJqBSxxtAqd2jvtApiezu2RrLbrD8jwvDna4OqR2XmiOtkEGZiD0dRORlWTJAG8Fct1ZE35Gm
H5osbz5zfkwF2ShH8DGDRnw7uncVh9X7ZkLy0Tu7LqZPreoYjbDtatphg9s9NtrxIQmW7gD9epes
z+Xe6+l/y+K9RFGW/W7dk7z/5KKEXAoLH5f/LPpnV8WeUtROlztvGiKi70cc7+sB9gmfHjFQeH4Z
DSiI8Zv7SDyX+sISGDhkfhfwvEBxg1TdT87s+kAaKCXrf0H3kHLkw0YW0TMJBuWvhQeG8H66cXfH
zOlNUsnzUvQF7elq1yMKhsnUv2SB+uhks9kXu2U2DZnda4gtmxih0RnFkYehrjL5pVvcpzGgalZ/
4SvjRShwgYbTy43zQDy+bDbD5E2Bs+0Hsj/+Ng06TliZpt3WXSgdXaQRtfkJEUucNRljL8Cfv9mE
ldfTwFbab/yT0kQ8thtz+3h1pQjb6Ap5pK26Hqizlou0FH1PPVMx3WIPvDQrEncWJrIvlCeL90WC
SFewST+U0rPHN//GJ6Sj4wcKmRHmhAxh+KlnhB1mE4L6kwDQvi5WMUoJErdrg7JwUSg2KakPqK9T
+6QL3dBBQan4ppxqBYnBAjXGqgyG7aJkPK1Ry7rlav/tOK2SWmLFfEJbOl96vja3IeVVVPZbU2eG
2deXvut4irsb1i/arMYAXNQ6ku1gc3pDbVZfpQlz11SmDb42NmKD+Y8SoRBw1tH4DQXVarDn+y94
TyZXeAt0VD6LYYD1P6pSeGBTQH1fVYfYet3XEHak1ffflUo446Qom386UODizJpNKIIE6BOC+yWw
VpU8nYu48SGV56f0pLS8vBj3MzVQnlZSTrMGNCgYeNDQn6wIXSTL2mY3MXEuURU5rXzpNjO2VlC1
AZ3lxRqmq6LnVConfA31ct+g0mzMSOlwvrJIpTVBxOw4vw32NO4XCwe6CfFsHuBw0ybbVlUQQeeU
3NlDkUrigN+4kW9dWv5oE9cNfAyBjlinVvxRxFjEoy3tj0K5ZH2r/QCq+r+P9vxSUBi++PiFaXv2
qpWdL+O7W6qYVz7wo52P6ksdNPidAvzjm4Eo5IbVpoYFVnwivNDaHRc75fLJtf7omcCGQvjqhn6H
uyhDNyfvBIc7rCinWURr8WotIXwSSeRFX0SUl0eR72ZEDNvm5a6uEoGJZ0iteB2CyDHFxKJOvEbZ
U0Jg0pBnSzZoiqyYfDmbIVWYZFKm2ICQqjNvFP1ASxarmVpOLaIq9M9NnzBLmx+TcSi0KLJzbnrg
Qb7QRvsp82nw+673lcBkRfQMYXfjqUBOSqAVUUdfi0vWl0DCfTamWoLR6wRFFLu0xjatTHLrYM9/
8clgyZcsiuhXkCt99bE3ASNX+xr1epQE6LFA22HKKKP9o/mZ3ZfPB4WaV/UjU8HrsHcSoybv9d3D
mSyaAE2XShpDFc7xGWGi3aw0ls6Sdwhupa8QHm7YQlIRvP94vAdpwVj/dwohCfK4S7nKdFDEF6Aq
ju7QwWd4QjZ4oozALgV9KqD3OYVzfrDneUswfnhHa3ml/hPkQvoHGchGTzaJb79u1C49Qosziff7
vymFcUDTWrfToKBClPGLEmgM26fii+1uxGbuBHzVlK4Ts3h6D4FErZnKA+fCoP6ne1m8pJ5E1uqX
1ZxdzLOadrgAiAOLALpoonflQQdvtR7tX6akHlNDvYD5uQfDiFKvka692i1acF8Z3wOXrj1/zUuG
/FMyyWfC5wIEbFZRgrJkzbsDTcgAGnlmc1YThkvjSIQlr8hoQ32LC4wR4u+U0+trtujiODqGnvdW
xdw51Da9LK0W2UHloesjutB3Dy7UXzMvJaA8o3zvAl3oH4xVJEU4s+yoQlHZKQVNak4+YDIvJtom
1WdHb8di65D7aE7kNDqbq02jQO5wCuyWVl9dR/W5WceDQykpTSsPFkGJp+75lo3WpRe3dAa1+TzC
JNn7uZOFcPBlgeESf88pF8fnrk20kls5IL9VhhIMC6vCd/qfHaA5/PqaaQQ4wfT0PMgXo7vHZq5r
+Z9N/LciM/zBEypP7GvmNlqRp6CZ7NO1eoVxvS0lrVbER6Tmxh8vFYivDf9jMq3NcZBcQx80GnMT
Q040Ksqjtn0km1wQ7wcc+rbmU9HzFX3Df0Vb8CBg0e7+AOC3oqPOEJpd+p8c1S756THLHqDYBTxe
EuCuTViuwhgIuwZ77ruJYPlavJ2uIibf6rlZ9j0HTDRyLvObOJCrZ5OYo/6/9XF73r2+TLbkWXEa
sLcGuwFPM6qfiEIn4qgnduJyLkXF3Z1AH/OIA4xpxw8Vi/HLi1YVjwyon+g94aVu5DCdPOIUqGHR
F9f299fZJ8P0ExxtUbmw5L/14c2n6aL63U4VT0rGVY3nAxkAtPSG4vdXa7WNQPUecCBcIXD3SH1a
JyfLztOmZFyijUo4tuLUeYzE21PFCIUpAr4ycGVx2ZOKascNB8mkGEgqwTybCE4g4HzItyTCy3A8
t2JYUFroLOa8kRgVC9KjN3juMEsvBtpoSxeBT/fI42YWxnTJhKtjQ8VaYItmGNHJ6UpvAlKKSXoo
GQJcgpvIUHc1+fk5DPhPg+0sKdoPVuUWR+QzYjNYJsXEEcALc7c/6isjf/ez7gbO8+d1yFMhWFHR
K17vU78CBji0rYYYK5i/nw4hWX14QRz5/Fq90/H5PlyMtYSdcHfhagzWhXdjC98k9NdBZFZaKQUm
vT/KTlaEuXWryTNhBo0Ndli5gGK34oCiakbUhEluJB77XyaSFS8e7GqPBpUjFXXDpwzaAPCsLPzZ
7sT3LGK2QiGewUQsw+bEeTo1ys+nJTQtZs/WMNUbK3aviONmNXGYj5QimyI3E6UGkU1EGSx80vM0
umfWVUgR6d1JtNMzOuffDJC75SyzikU7UmtA5vZyg83mQr426w8uwJIdfgYn4bXPmG9kbEk7rjfA
WIHTlkXCox/hcZB+OE0Ns9f68BUrMP/vAFMAicU/+xXKJir9vRqkJSB4aad++9yfZ/yt+3L5v9yd
f97GcYvljnGa9whkp95b6qn6HnWKsUnXhVr59NLSHkU3ww4Ry4iWo5eqM8iiboldbwv1lJcLusib
H7W/yQF5By5vZ8WRYCsxc12pfKDOcBWiOdnU8RInJjqTzUcqVfPZAlkWtFoOyKATVfOebclMeqYN
RhEWcEmBVHsSnrhYKc65V56OiR0IkqwwcFsZ64mooig6k6TIlD1IfH/xTZPpDt0G0CnaCYNSDdsq
1s0RRzmZlEYVyO74olTc8ByqRHaRgwbdyLd5v3kwRKTsv0jroM1On/6xxInd+tK/rB/TcvScR56y
OLeq7NtSNvvDbZM+33oeFIY9kT3wdUp2spy1TuAsjEUozb4Osq8j767CXeZMO4BrU7+pzuLQLX2i
sSuDb3XtcY+VmoOFqQYxEYn6Hq7Ub9dEoUy6Hj8TgVabjL54tZpKECLRzRf55ZefJ2fWqXdjSDei
ZbSJsKDyPBuxg6uPO/p2GAEy6gnCrUtQsuJtLFwrFPacUB912WVCc+tDmH576xKQj1SqLPk1QPYU
LQ0YaoKy2xR+2OemLajjR6MuVx7KOxkzYRIsHM7qRrxPVYEA+I907lt3KHNhrgfDfG24J4cl8DcM
oB9Py9CIy1HJK5QIfYIXa0vXQr4pzTdxZ1lB/tSI43bL3lQVGdls3hU3uv+QJgeGF/LvuAbgMxG9
jAfaYZ3UpxfWH40h4qE+FjgUVevCfL0Yz1MlCRb/IVEybB4Uiadw2IHXnIXQoS1HVDUdHzW+upB8
Yz7OuW3vnPHOzabGJX7PMbWFIkW/nb0r4+JiKNK5T9Co3KCZU9Lm85tXsFoFyotHl8CrbZ6J7kNH
GDBswMEz+wwMIlZbpRjmLBFwVWFNMRD4xiL2JOpF/0KfcAaP/koJkkyoLcN9okAS112ZrUQn19PW
lsOyJydNbqgnT8uGnguJy2UJN1TK7yhLvSR0QNJUV8pbUXtbRFMJwWcN1ZyiWMQa8KuL5HnGtBjz
swm0rNuOBk+sRYPSyftRduQnalDhC+HxOnBvDNQQHz142VbXJ0mAmsXcEH2mw0aXJW7x1OjprJZw
pa0wXB3bWB9IDZw0pj90dZWjqIPVSLjxxc5vh0GGnC8A+KN6XBmxB8H7b0o13EqDbA5wQZhW/nzi
49+eLbSPSFKx4Sauk5m88aftRB3QBTtnA70CpbsPxXVH5yOnmSibXJ0pOJ6FTxuRARdpyhQ2uXsr
3983RnioaGru4MOSGQT2W2FwadnN+CgRpS1irZSXGgwRNYpDafNAjO2DoTmIWvxUkMzrcfC9VU7K
WwYQyEDp5bXUkjUaUdlkRj47f9V9vCBDwknsKYkM5caok+G6IHvWL8RMgC3zGNBlk1ROGU+ndwra
3oe2IJZ1biiO99/qDu2cWMcf0v0AcDMMX80oEq3LE1GuGiWpau3WWGb4S9r1OfTOJ+2owPbtfJgo
1/phAyJDHImNvzSArx6rl2DmkgadnVeCoFO38yBQN3yFSUw2dTYNOTiT1n1gnLiSBbGyMOHK9UT5
UKrumLVTzPcrt3Zn+RSPjdW++Lxjh5ngJrolVzlfNe8lNB2KCoX1OZLEjgKdmgg6N5K+reuoIIBM
n5SxIIxgYwaLLDkZBI47h96SL8Dsh1GWQtRaC8S7UISHXEe1UxnxNW4juMbfzvlIuJGo9IxGkj57
LpcWv13wnMDIcsil6y3MRiUxXarnyWl46BDzGpyxvmxliT0LSV9QCtVoXmZd5m2hT7k853DZocB+
Bi40dxqSJY4BizDOdirbAkm1jua33eIvQhkRdxbdLs+5GJ6b32oBNcn0tEZe4Gc1laGmNR3h9IeV
Au/jnbw11kY7C7793j6CKMAh2EVjGf3LxK8bjJTe1eVVUqL0k40gdg7P1eJJ0G6iWLo5i+hIc/eM
62WeI/muriMjJhNYXxjGpYc3JisvO9jmYH6/ybuZQ0QYMep5AJqAMuKeXAATi0ynJZq1xjs8z9IK
MZ5vK4c6z//gPWWKPWuB6q+8D/cm3Q8E8roERjWKVoMfGYyzhr9UGjKyN6ohH+K5m31oG38XucGb
kYAWQV5X6iKU7SMbIjGCANa3HtVDvflxqrH6eWf4WOtvoRgy3MqeQVpnHjktSUCtV0NQjLjBjpYA
HcwRosXkf4XeXdWfcAgeo8/HGjSM0i9DUJNaihL4+05NxQHTNAyhnvbx+n2JB/WaLWgtX13MDcUr
2lrfzpK5RLyLMyPRLvCpcspx24KyXff/+o1fgZOoyDI98N3H/t1gts7s2VWNajHfZixbmunFWXrY
VN7RdjuZCIG0LpzWdz6RGetaCCZeHDaTRgl8OdzJcOTdh5in7MXW1mx+VS4bA8B2yMwE2M/XV7Vq
eeys+dD5hEXD2z+bUCdujcI6lG6TnieTYikj+13L2cuWnJsuksWgIVza9eQbfbuDzNoAlniNFdCu
iKx/90fFLg72m198TI2bRuyBbliMGjTou04UVFu2TCtlExbvgani0PD4c1oTDxL9x0+x6SiEnEdt
ocmk2RmbO4KkB9msjLJd2bKjqV4LRUfggWeZ5IP3NLBO5xxdRYUzxk7EJdG6fx6AdYObhnzd4XfM
Kfi8J5rb258kHMx/AermGcAe57NvqjwtkeMWg7y8inoUdXTppqM/wEXFuAqvKhs/RH8BcTKwFojY
X6/CWiLse9wXAlsmO/omQYbkS0vF9LoEiujEhqT8K6zAE3aZquHJRZ80x6O0btPvsGwtYfiPxE8e
fW1FcLFqf3V+xP1jE0QqT2orvyhk30BpYPtlvihpxNmR+2nA8YJAE5/GwwuYyKkUX5Nrjk9WZwKG
immUTZJM5BwsFXryMC+K1PUic4JV+KQkX78uSnoKUy4gPxgOac23Uaiw+RqZ0w536xHcDB1n4l0Z
+Z1qkCetKhff4GvQhRul1EeRRfVXGPX7yUnJ4IzACh2cif2Ik7xEbbQio+K83jqd78W0UyOvDnK/
Tmb39eXj/oQ1AEN9L8KIRCIihL4/dwAqZQsODINGh6XyzdyNZJ8AjBwxD4E8N0ir9b9u2l1xDorC
MB2+kiQ83pKDawWQ0JmKCQoK0W5VpU2ZMtUIJZZWy4WsR65gufezpnIMZS6X5YNgdPX5MNHuaVAk
4ipNmsq3M9aey9vLOCnAuh1H8caA5RE9ID/gMJSDlxsyYUqcfQ6wnH+sK8eC9ZsUuYsRfnePyP7F
SEaUKusCzO55LFHC3u/IUw7E1IFSbsMh/DQ4aSq/UoiuVdm6x4Byrqp3xarAHgnHKpbiV8FT5aTl
OgWMh4y3IXRHxESI0iuRgjhZcw8FlWkPIt0JBQhCch+9kPJmUz/6WuJCnjSbJ7NaqliWpc8qJYIi
SphHe2iwp1Q1OTfi9yX7sZ4RKbVBGnkEkDJ2GqDnlMfr0I4Tdxw6DdR4taMngoSyhcXz8fQV8uZM
8XcyBuWDztzC6HiK9isxGVBsVql7JGwxcOnmkzEwJxf6ZdmDDgmi3/HREC8XpL67Rzj3+H9x+oiq
xr8vHM9vXMkfptoThBv2SQ9NqNo7l1QmIpAgrcM2VINU/CWwMfTt6Pdn6uCBuJzf1K3hFxgVBYHC
IbfJ2IJA1aVVrXXEVAwAZuHiEcMd1Q6Wmz9xNXeHWviZ1R2yRX4uEADKxVaoqgCyLAQ/GKad6OyM
FLbxePO3FUFTi+QYedcHIqyCIW+mmFORKd/6fwJHhxilQQlVxRm65U86EuERpEXgadJU+jMufNG2
43sozI4nHsd/Imm4XTzUHj5RqqQGeo5SbrXwtvaDqV73ZGh0Nt3PwVLTcoi1GASGuh5sZszdTsWo
T67/0Wb7RoXpfZV76CqaaVOMkSxHZGwmWuFxxemxWMyrrlVBAuF9mvSFG4R7ac3GiB5WEbO/W7mG
F++OBBttrJpBTBUTSm65bRnZWEls6jscKp9nCu12bLW9FVswa2PRF5owASWXh2MIkE/bMZ7qcGU+
vGznyTMhw7yBQjA+rbUqHiHiQcI21jAMazDHNvcDhtzAVSEf7qj6QpKhy8slIYkmeixUsYBseCxj
KpcIetDhPj6MWmR+ALflFzmjJRKcvYzKi1d3NbxSNV7hpyv0BgTRLCrU7ORbhT+0MqW9422k5Mff
33goZe9EJqMksc+pv+9R+aIIuvzfI0KVwkadmgyVGYnnTpEIedOn2gwEpmUcbivGePS2xn6xNM6z
kGyQxHB/VXchCsWG8X91lpSdvfNbztb/+LW+2++9ShZN38QQ60cwYSn9lAMraQw0rhiSlnMn3k5j
qtr6vWo0ykva3whALYujdP0l8nguKnI1N7PiJvjcMfL6KVK+LtE3aM/z/2Hm5vRaQiJ2Q39ETJoU
9p+UvMWYozgiRuGpZSJhQWep1WtGqiGXbN38w3itl/ZBmsmJzy4fDFN9QrDEg7Z8SZmfZ81PG8DL
62Cv/9EmjMyR2RVa5zWNFBqFEQbQjW3Tm7DwLiOMXeFDTMEdNGZU6bIq1C1FHA92tWNgM4GGpiXl
zqedu1lxhzYRE8jaWPuW52rXqLIPnPjHniGPvYNFI5FkmKBH6wExgugHYED4PPjTVHOsD4nAYK+R
qBk9cDiCYqUXDSv90Cvk7QV4ExHAWvCF4yaGniWvEMDInEpsqDO9OjoShlSgBY3QBQ7zthOzyxur
jujhAWRfS04V5UEm6hAC2qaab/Ei3IBfQEYvqehICUUXmVV6c+y5P9mIxOt6fw+/Oi3jE330y65x
B6AWQzI4tw9wL4Ussr+1Xh6qlUH0O+ne5laOOh+injuaH8jEkwHPoqZ+LJedf8mQkxsfKeuXIFYS
osJqcB5M1xc8pamcVbix5n0NJzHs5YzIQQdWIetP7BehU4N4xuvCo+LDxlu2mJ094PD1cEfJnivP
Zv7OMU0b3//S38kxYjZUk0O1ufSWx9H3BbgEKvYb3ZQo6cuKxJfULN2XHOX44ZBKY1QQSIaJ0dDY
zMes6REDuZg4NP0dtIM+z3mP1M2FoytGTb4LdwrycV0EJbTiMUzwDVwwbCn/np6/HXa91QOUk+8j
l9+upHCubDSy4bA9TyiWAjfnRz2CjIYc5hOuK16B8opfL1BRf4hmettFQQ+j6IgzQTmq2VtTsqiP
/tfdGtY5mlMBDZnCaJ1XkUHwHbsLoZu8Xu73xsCQQzv4aBeMkDSPgP+pePydN6e49hiofF8asd6n
8FXWQInqEYdbeY3aACC6y1vNGQVFqeIzIvcJ8zd1FBo5AD8j06WxHtDYACWv1hRmQgRfBvnL0mfk
iMThLXAGRRTLxD2fQPvEyon2th1xbCKwxhQZqH85i2kfwTNkdZEVtBDKJddMfQwa2ar/WB56fHD8
FjYWGkBtKZipeddbKXVq0uqXVKeTfYRYqWOdGMFFAI8rK6CEFzEO9PX+rBLvPCmvraChTKK6NUnq
gmA5s2EwLGGAjvjQ/84wmYGQ0Fy9Z9jNl7XsU3i5sIwG1f3ICpdSrCsItNM4VXyPungFoyRWorub
/MC4u70ricoE/xN1x5gfhPA7rt1XGMAHr/aRiBDSgolluZ6/2qkSjLjFDjqU233c9q8FOe6WwKR2
bx0eKyBruUjjJnBoB2NJ9qLd3Pk2YME47Ry+FzaZ/acL+OUHk3M9ioMCxULJOYGbWpPTXv0r1RrK
nef4Vs769F18vDoyVspyWS5Ts7OmH49CvLp6VhhNFvb212mHxYma++4k9jQPbaW9paTQqiOJd0db
qqZX9LQRCFznN1IYUJkrill4eZbq5ZQOPbYWob+X7kBYKaR4vyFDazvRJo6psx4eJ78TlFwfR/aa
kRkUvEXio3Ql5XledBDZABvmDfNVYwopwv4a5clD6jiK2RK3MfvLz2BpjTCSAwgzg9goLXrBH+IS
MwuZpniVJwJp6qY3gM5AjbnGTXgR1G462leoCOho07PZs8gZnVX/uJ+pJtni+EJXfvY7DEvgaMzZ
/2RyhWden/RG89qg7htNh56ZL9YV4fhUhU/BvmirD3uzM254jnfEen/7+2SNKJ+NQLuJm/H4rg3u
3oPTTg1rnz8ZFFbchI2rNuVuz+xZDwdzM0wJYIeaXJLVqfe9oJUoT+51EkRinYUqG3BBLcIEZ+CY
WaqRCfvtrLiCepYds42AcZnyDuyKgl+BGpCMl4xf3GE9JEB+j1/h+2U3sjW5Y2ZVZPk++c4nWIAl
Fsot9Vj9iRG49L+1Gj7xrJB9YSTFH/yXHP9ZEQC0vl7s2vd+7sCX85eeIa0lsAM6mOhm/i+Vf+Pu
KuMh/gybu/AXavQn/+UtTB762yjwfwfgjLZ5mEFW8/phufWit+iLjhiPhJUO9xCwMqdIImrO+m90
Ga4WQryWSV5CQ00ZRJ2j2zYyMK0qMN86LtKqSeoZKX1McpyheU511kc90XfNlDOV75wvwapYcoOx
j0A8Jg8RPLW8boRNjHSiyzOJhdwLXImQfsgJp+fLvUjNiuZ7xYRNRkzlKHcIYbtEpTOw26yIYzNV
QKrMEwz64WMx6XxjwBvJhWcmktc7wD30rwm0XxdrCjLESxnrD4T/kcOx6KU4X/g5jhyndr5fmH4J
97ybiepJkZ2P1w+ZqKxip9XJCFhUYlDKdJcAWtM9W3q1em5dWppSRHWPjNxYmzh9123kN1pzA5vN
XqWOR6HqD8iDL17BZhlXj5b3vVN1CXjSbVH7ikVvrn+Ftp/U6yjQAsFUzwEfB6U8D8hm3xA+NeMZ
0uz0qiw59vJV9Hld4g60iU9nppLwMdfXMfJROv/a+0GsIJbrIDjV5DeY672BRCtcsTAp11iLHVwL
HuRndG9/cn9xy4hqQLScaXtbJEqeJS2RgBdAH3723xKuB58/aXSu5S9jFhculY1GjVUNhUlEvFHo
fuWXS+UXQQ8Yx8Gozm9FEEZQP8XUaDD39ZKSJLqsR+r61oKq9Mz9v/35a/CCfQEhWUUXqNoK/xg6
po/17mYwyEWEo7Jpdt17v7jOpwjJ/Qtw2Y3htSvyTXwf7a+Ho8CJrQzmqA7uj+Nj017sn5c3mBp1
2e+afmrTnZ8F8eIwC4dP4qv/s/89wRm9Afh5NX9eq2udMcoVCPs2dTJKH5jSbTnb7MLN1mJchrGt
JBxekGkVhAPcQCZE8aCWv2z9gkQlNKdIC6uu7rNWr+mgliZMJAnwAxoX3eQFZi6xB1Akt/A2vSB5
7Rtn5KeBmDM09biw7sLs9ligynIwBx1QJgQE+0O9+KduOG3J3sm5sOdL6pAxEKMfjjlsVysrHMVf
DpO/gaEhuQKIbfLw+J28IDB5mnb7wqDlADAojrSLSacWEjxUdR6oPytrRNcgpAEHiPZvywMBugga
mhoS0DOqV6ZKEkPm10AtCCp8xl+CcjspRC5igpJcMLcbnaUnmWwE+a3z4HC+5wDMTSSiWnPDZc3n
Hs89lC45NkITRkk74s20deT/RoFezNe3KN4u5kJzv20YDyCANgtwy62AtUNOL1/EkGRuPi4ZuH/U
+GnE+BAaLNn6TNP2i0exhR2Ehth2eEF+XrCxnJx+mBwTfLDgIWgorSAQEHHQMeh++09dtTaS0cHd
ku3ttQTu56z+PYQyJw2ryAQIfS0CSeYkAyo0BGZ2hhfGaN/ONlhEw20/X1V2KS359PFP3OUijQzy
SdmDyRdmnz4C4BJ96Ufg5XC+lt5OvZ+k3K2Q7opv2k5mvrmAbzeWqowqUCeopmm1LNJKwldaeI90
d1W2kGzTWgu9XyYzSAmWljo2NHiV2s6+UQ16Jiu32PoZUXlpTjkX8JgE3CgFSZExHwVm6BszwSzU
ewPLMPGjAbQFQeIweY0yZyw2Qkz7Hu1WmuXvWSfBmlIwkXkpvq3ixq53cdEJrYyZHwzXdv1C3I6X
ndrh8CE5xxBEarJFUTeL2IkBUF1RShAOTZPfS9AUYwMMnUYVyjNKJvwOEbcd0nvhpVmdDxXZfW6+
bYPUZMLHOqUJqLeRL8HomXdE3rM6awpgWlTpeRygfqmOza3imd/9S+tV63hBbnyz5Qqs4cSQA3PA
S7osIQZlZz09y2w6T29+xAlf9wrcSXDlxK7j+WFhNVn7QG8iXVi1NkQLubdLoFeuHiSpgYcwEMsd
Q8/aJGS7lx23lHJe/CB+mnY5m4jtDi8flqUDqnorlaNEVsIQSnT3YcpOpqoe25yi5zmA/g4BUmvG
aRiYjQ40bb2+gTGtt52FS3FnJ5aLzpyVCPCHv6jCd0ohISbMbVJdFz/sJFYeaLFFwelm3Q3rj4Cj
eUYdhfPe9M8zOyPgLXoORYPIkj/qFBOjKWVU80YN6vj44bf3AMyCOeV+HPtR+DAn+a+kjRIYoD0G
9MzNC/VZ59BEFD8sxxbyk1HYhAif74qN307Zzl3kVEwUMJqiEGJl2kjc4XdDsJdQ+wNVfAJ+JGau
5p7K21uKGEMwRJwbJyyLJyBzRTe6zAuxz4SAHJ4PBDIvOZCDDamGmLhhbWdu9X1UOnNNr9CTOSqi
88VDbrl+KXsUBrxP63g3QgyWFdHbL9H52ZB/7QrawWlrqVI3Ncu7sIinqIUhCcQ+/x0CBQxsrHyt
vVk6F4uiNh1QCnfMuek3vHs80h3koegmNO4/zf0nitrtN7HtVSC1Y5wHoGkWwem7bDUf9YIsr/Bi
gmov7+QfyBRkGRQBJwKU1pHijvkC3WpJeDA7MiByCA2QKFXqC5O3cE2GrMnAc8EExEpsUEKgm5wL
REI0OaL504znRcpD98DiKQbuEoUfNsWDUBv1LDtLR78EclzkLv6HzSG+cIleWzAWUdkLE0cZ6D79
e5UB+qzA/653BAlDegZeeylbXxDUenAAtd+ooeyr+xaV8HJoS6aEzPLfN03kTPucURdF/HCYusGd
TSh67JDm3hzClAkYmtrhGvsq39G0J69lWyO/xPLs/IEuycBWVmIMY+vnv5VXHf6OdrLgVcIqRnd4
r68D4eTdJAo+PMlejZh8vee8C8LpP4AdaboP+y7xpVs/U7W+h8JEsSGMQ6wXsGSZFPLMlWLTEKnz
rKFDKBXTFmAUQjxYz667jBQG/VG7sk4YAoW3yo0KSThhIt/1ZXhLwXHikwUN6Vhc5DaTPaPTMIko
iBEdLGqeNYjwYjOwcswV6uypihDcIYIwCONfpV9IMcrH4RyR0Pi11YfL3rp3pXcVdEuomCt6AweL
5QUZbG3depT+TRZ200S3+PPA/VqZVtuShsEebmGBZ4Nmh60FLQlhYlj2QPX/DmWjAEkeLfVwD7S1
s/RxZ/rs3jK5fk+mvC/OF6npHzYivJDzCEQOHe7ZN2nD8zyJrztgACFrQOCNd7ntNiYDUyPJBfIB
+5p53jR4vtdvm03wRyzRmcL+q3DPaQZBrRwHrKeZU/VXP7f0ePsWF9kvzlvLwPMJamsarHuzvqxa
zFc8QXM7EM97qSlv4Yv90PA5AZ67v38zjzeT/rJIyO6tGHIOLVz/7oH0hEqcYpVGMrqYKFYYrrwX
QQtKZfp2oJBQa/qk1GZdpzL96jxylplfwrqc+cROgBkkxCyuT8VDZQ/Iz75XuCNW8GN4dSS7Jzlq
xLcNu3lYwfgakVcM+VX7y0otBE1fzJYnWGTEbDkxyVlOg7aZGq6+hh7esqSzD8c5nROgMyk8yMAf
ARbJwi33fNhN61aR1j/3vRu8B32l2Xk30do/sVZzXV8rBDj/fEKvIZVlvOYSwVVtP3htjAgC2DGE
XofFIZmhlfi+/YEkgiwm640xUh6yFiaApT48nrIC6xwUP1oyU9lKYj5YuLSgY8aP8YujMauxIQls
mXvLmd+pusW8hmOplIwAEIWHb2ctKyvElSlPrm+DL+eX2Xq3YIeXbR5rFY/FpmxAzLLIQ/Dnbrgw
qsOUY5KdKw1dStPa8xiQzwalQvejYZJzxSYqeOo8KUdN1bv1F6bjI5ritBlTMPsEGap7gKQeeSHi
qO5sqlNm6QdS71a98UvG0irOTYRNDFPY48/+2NRpXuImNDwDITkhEG2mNPkryjuj97wq1KgEMPt0
e50XkW/Ii160GXb1Vq1d0n5jW5nqdJKb1IzHYD1nS2VzWRZGfpeIYipskztuk+xt8hrTPMrzA0Jy
6NrXBZJBkR+iq2Itcb1QmXfLbzEAWKTmIfrCFazZjcMim7M7OfMfho3xvWaoIGxpG7+bqQGFxwEm
zeANoUtDQ8WKXZTWQVTV8O5z750E6Rr6cilRMY2bKIiv1vxJCSvuSLuq6NZl4LMBC3wGo4wKCjqa
AOfIPe878jvflBVO2ZeeCJxaqrucBH78ipCXom2JjLfFQ97eDLopfY6wNynbXeRO8zeZ4OgA5pZp
O0jF9WIwsAcI+lnFZbgAgZ7Dpf6B14ctgDjzXdwqC9CLKuMPLHPBtFvYODNkCEo6p0i7gQUEdU2X
RCqLZ+v7bPHavkwEcZJiGabpRv8sM6pHKKQkFqnY5SGF6LakMLjlNDTLEb3+Q2sqM+ElOOBMICnP
CCsXYY3QIEbbaqeKwPDBAGszou/0brbJR7OWoJB7NRnv48XwgVGHfZy6AvF7fhvaGjk7pMRNgqum
VSaWja3dStMMNxoKskSyHcG+7LuhEiaYGBdCADUuarGR5n5oz2vwp03InQNAsOU8dRURVcI287Gi
Q7v8+cRBM5lluKgg3vFd2wT3C65rb0IDfZzCcmtVcd9qkg7cH/JHnurV55OzByPMmOEWEz4Lhyxp
anT6c7ndKSRyQTbzb8Hn3L6O4zMUUv/K41b46IUnFDq0OaV1DIzdGOEuYHW4h/i1tqvbbRafKaUo
JISzeQxa1YS5ILK08sezY72wnIwmVVlmezsj3UqzFrpLhw9u+50hiFo59E2kutJOmjywCzErWfxv
M7WiycpzkH3GgMzc7e4F4+YE7e2eVI/sJBUaSnMoQDDMp67RwAzteEWszlediW92yFm20LMSOsms
yyWDGWLN4O1FbDbB26NFNn1H9wTVZDRb9ke4E+JtxvDX+/MyuHk8mArZmkWYzPb5t1hzJOLuB3Im
KWrkGIgJIHnAzVqF70SlHIMTId+kuXjEf52uYhfhUop4hi2YHObckx5uFjJRKGDYg3+/m/ktwhhk
6Z1jXqSMK8s25Hp3bDB4Mwra+T8QKE7qeujhddeO418hUyzhd1i3hE4tRlhv0bHkwDiQesbEWgak
QQxyfn162xlNOC022AxcgZJ+4RTdx/0KzJhP5dXhBDs4JsctNZ5Cn1vEJ3cgyHgi9OGkzqKrOg1n
E5ihDSWL8gWf0+fUSkm2hN3ksE2oPtd620oBBx216LpdIgNH008CyjGRbFF0U7EKcW+PxhaEetvA
T+0v/YkYHr5wfVVSq0XCLA1+KtJVRqtwNLTz3cjP0MP5AKeB0gwA45fL5mg26HUiyJx5YdPmAwSI
umgndsCGAj12tpxmldv3qnQlG/WHB5ZoHxCq6oOWgnkoOz1j7RLHlRF217V+OARLzLKXfW7+B2K0
gE83WV3yTrbmyYtZgA5Ey1qpI4XUeTFqNl8xXVcSaLPyjsI2H1BP1KRKiUA1jtFOKz5a/5moT57z
Ek7/eNn5GNIAnMHajfc7TYNLB1L9MR1LQh3XpbCeOdHjZ6yRt36lTAC3jmjGXUom5fzhVK9nP7lf
81lB3Kl8UDAN28+WmZWHuIEOvFYQsA3g5VrTF3L+icq6p/Zc3ne7/ZnrAXLgw/hwlINvCoYL/t/0
F702EEcQShmf3wMa+J7SwSiA/q+2fcauauDAbPGgxGD5c1QwPWOj/LlL93JD3TRQGE4d3uFXSc6K
FcP5b7xdRnZNdlViVD8Js/q5py0bVYFZOROuK7+LzIQwdahbxsJrcOKh3YSSHvkYxue8YXHNbnwR
71iZcbiq9Qg4PT+ytDDVScAce5NiTxQu+IUMFneRC+Efcbcr9PekZ9kg5n9A3WC2rMYZsZyDrbpF
QYrzjwAwjv5ajkfh5Ucm6T6NtB+rKpN2O9eMzytjM2KLeixM1kEzt2fjrgNxgHxzo8hsigogoSsQ
GXe6nOPimiitGK7xSxxdHdMCvx03DtJldY4BlQ7Xj3clHCAJK2SA3PWJmnLQ98r4msW8+lxcUYKJ
Qfwczvgkb2QG37PP/5Rqm/noOBQpjiDnx0Lz0jgg0KEEJ9zahkTOEe7XypED4VVfRgmkwRKtito7
Ju91tw8/HyYA0J34lboztadOYhoByMvCOG8xB4zSGBMnUBUV22yZR7A/4oA5PSKBADl6kWVC673x
1nb2chOshhx5yWk+y8BKAjQLX6PXqWtxisImQv0U60EOUihlIB0V4NuJTN+1x/NDiAX5ZhiHvb5T
5HTBtw23NPyf/9MC0sspQtp5MfZZpOlGNQylf4a0ayDHd9uac/PLFd0VOJ+CkHCt4YJXz7fnwRlM
uWIvf8xz9oCRa4J2kSQJxUWcHI0KjUTal6w6k88mwAmEA/17i17A7RQLH7hSWcLi4yf1Cb6PrwjT
Ki4S0I6L1BQDhDXsdb3QFQJL2jMy1GMYAUULPoHnNTnmuS4cUeq+WdLZZAyyEBTccg9SD00p1lzR
VqVkzdXonsZWAFovrxHQSMK3c5fONuvMpc6obdFodP/tziCQPB3YrAhEdF8ut0nC/1GC8F3Htibz
4bjm5D7IEDO6hMus+S8MHkOUQjw2CSW46HFSV4Fd2lXKI2KAgnQ8cWbhPlTOJ8LrP7M/mvazUtp6
T2SD4wI8shDCQVUgrdNizf9V7exaNivBFkSi5IRO1+yVE/K10rASFZKl7EvNAeHK0Rb9iwPR0k0k
sFeRxykgBJVDnHpMh6VotZetfAgi1tWadK1858G8b8cNhF9OXTbFq+9S0z65Ifviain848fxrb4N
9dVW22dO2ZEadyWZEWnG3ae5BWiyZ5pgJRtZfYoSkdasdpztKN2llpjcwVw8AjR3JgXujtqaCUXS
xrzBPXjhpPoHrUqzfcawwKb7F9HK1mnvhuI4ZyCtTc85dSY+EG4ZGgPHlo4l/kZ+pBhXm0vkc/f5
r2tkaff+kgqSofq/sa5vk05ek2/xmkqQehdQa2drYFHRhYut+WKAdKqRYw/1hz+D7XxfW4BZ4o8J
Rjt0QV9+/hibfNb55idd4CfSm8qrkk16dHW47PiLSzY3kEbSce+NlrKNdIqBmT8pYW7Ee+3wYihA
PXu3VZ6mq7SN8TsENhX56stuz4YWponwDiNAETE61glBpclaPHXAYQ50ZJaFn1gOaqN6AYVDiafA
hpfEvdmaaTEg2IFWCGMGwm/ftybKQ4k578JB9XopdXR4DcVkqMzomAYmnpz/8ji8nY7dL/d1bvqp
L234GUPf/5KJ6xpq/teVZpy7QD3v08uddtNsOpLa+E0ilaZ6oQPsuN//VFMbPn1uoKt/c3VpQ1L+
P6GF727r64mXVlYo0AYvykxi5VJi1Zly49yX7D9jwMinX8zMUWSB4nKW1iUa38pQbePwTO84a7CQ
O8LTDaazavEuOvPgdaajbm80+iwNHlhQljfk0Ov4DLkIV9FFEkWC/KLu+gjrTk0ux9xfhuoOJ5Q3
hraOuQyzxiinaJPjin0LWx6ktoouo6EuPRN8j439ABi6B3Sn2woR22LawceEcMlrkUmEbIcrqjZe
JGs3Uh74VSz6UarV+Dz2tDxyTSQHQUYpLInZmHz4tlAWrQVGPo0gaBHJJevvqtyYikXQth9hejqN
YSHo5KGzLJVyY/jk1R/T15iz0oMA8Uhz4puwjSyuRFgRIiRqAVsvKpLV54x3kRV3ew3etCSUpazP
/HohvdnZ4dBhfYTSzsTS1G9GrRUbGjbSKUpPuq8dN/ITM0H7iwSSYdEV7itY8MvIspSGqziPNnXg
8RG4cdNSz2UQey4iA5PhJ+1HxOG4pDkfT5bixB7y7C4hsBBFMpRSKVgJyYpeFLV0mzDHlPpEWh7m
LHJrRZTOcnZPr1DH+V54URB5HM1GYDWg8IHie/NzbiHZitz81iUAyV2eLern9Fw9FmRzeT++9suV
KkruM719bLwICwX+jWoOEp4mvoo7wNy9QM9+26fXTP2L+dnGWwIBfiR/9v+Xyp0jTnVDIztLP/hx
8YKHt+4Kug6nqDfHA5WOK6k9jX/4vcczSng5jA7BCZEom/F7NtlZ5XHiBfeY5pfcX00k73p1Y8/n
MjpTovgSCISjnn1caE6YDMrc2F4RQ0IHeqUKBXZZ9/GL74MawQhfgrVvA3YRp8PLlkfPOoD6pyVG
lgeRK03TLcgX+2lYLKSfD/ydjC3QDCubgJdhAmPB5ilkIvNTekRw+ALB9f+DhbQKrDySwOane6Xy
VclH97sQzrOwWFeOO2dCIiPJsI8ZCKW1S7n/wY1oP/ipau6Ev7slff0JWcS+A4fLfuFgpFECMzGt
qKjrZAt7/QRA2xB8LZSNQZoeSKLn7EpBvRs98vzuqOTFroaik6SIrZrCY34dsW0hXX61M+7pmE5W
dowwiDCHCHwaclTXSFHeZIO1X6wiRsbZ213Fpg+pYBaM8z/fDyxXiWfI44yWoFwayxfMWE9YfHSd
GL79VWssnJZGuSJ0GFHj93h1E9dhFvyzcaCoXb+bIiHsZqgByi7DAuGO3KQLR+BggmeJC9SYp6Sc
wHesGBDaA967XCpV32Hnr9P61Ptqfmen1j7y02ebX5yeCm/wZAaZpVxx7nAshDVC56iopGfpeePb
M+SZWMSAhiKyJuNqUKp5DllEB88OD1zJsSrY+1DnXkeXbiyEInhaa55ZgMK2WgYnUYLXh0vdQQ5v
lZWZT2VlKDObHfqSna3yfphJQryx9zXDPfbCQB+Z2Q1zzld9D89ErvKwMenxRwbLD39VKDMRxTiK
/DFp6dnj8hAF8WITU3XBHu76vXcWeO/ycXWwEzYRuNGfYK5nv7u1UEdS5JHSHbP+uTb4wlv3crSo
6eKEl74VXAP73JvobYTxpAoDQcbJAT92OwFfwIBCtFxVXGziCMntB88MwjGg1p6M1h7Vf8WfkXo3
WvSqm/C1317zD41BSEp3bnB1SCFkXh00x2rFx9pK1Xhl/hOAnphpQoDjRkbzkyN01iruE03ky6kL
dC7SscMymfmGt/DwrJBTYfhll6ZO234uGq7PWmA0tg2mN6MtxFT14A5CahiISkpXFlH3OxBw6OCd
dIjrAHnLyQMYrTD7nWCU1ucssfT2NL83x3F6gdudn/kgq2xWD7Dj9aTGRkoprA8C6gTlCwQZTTbB
t6Sq1DhB+BrnNvNIjlwuJKGFxj6K237qdR1HgLcgq9TC8HBGPPinyLb83wDzdrIOTAWF8PmoNZ2H
bQwkWOBHPBNyPrBc4FbZuBmnNgibSkLw1+uAEm2HeAuY6EVZbiqVExaBlO4aJ9UDIoqhinA0+Shw
hcBcxFdu7z3l/uZe54rw++j+xrApzcp6LQxFJXPzCVyprz2rKpE5vDEFhXrn+tDHpJwarmyICOK1
0lK/r/TN/7KJzrVTDcrte9vT5sftpTPcG77ZzreMzEjzeiiPjPuxhXmuSm0I7AGO8T0iGDSWgL8l
FnnLtWjzA1JXGIiAwra7thczwlCNHqfZD2B8kT18oC59bFvqF3pdBdmyIl24WZoUsjAVN5M0vSca
RKNooqwytzEJFFaZcC8uDpOWitbPwLQohUjp34U4Ld06nign+3xxRr+N2EnUSIJaUiup/WK4xDC+
sGyNMIJJckN6N5qWKzEPiov7mI1TKKF3GTlUpglBkuInqvgRffmjHfpwzQob6F4mPrbLGhB0nyEC
YrfmkF+w7IhUiFYON9H2OJk+3T9VG4cNLnfiAJYmdjD7cp+N6m/VAXZdSdcmGSgawSFnw/TlT4Vg
dykT4Dzinf+8QPSHL4mnH1yIXD2GUGH6lZoaJf4sStRjPNylOSWl8cYWwjreQdB+NmuG+rQbVx+m
7xW9qKsw3haz864EKYo/dClr5Z2N0e9JbWe6UYu2sO3awSZDmW7ZriuCjtivMO/ZVX1XRV9mNTEh
o9+G5aSQuh66BB9dZyZgYEkWSq0zJ0M3I9H3BWCPfE943MJt0/TI01YkpI4KZa+Pm3nBR3T52flQ
Z5TrCyxn7IbSPPL0bjn6shRuoaxkCRZgUSWO1jrkThDxYiZyMAcaZb7RBSO5wzQYwQC8GliymQCY
SOlVRi0ot+v2zWSzqCrHZoVE4/si6ACWYNqcbuOjMbHMe3Kmmp56r9+sakiUvU27WmuuXlPW3bD1
MwZXBXNa9g53VizxVidDRlzXcSg5+8OopRz3kjD7UnC4muH0JV+qKbtDfKl5dudGT4s8q6fIjfnY
LdbMc2lSf9ULoak56QRTWOYlV0rivHqGcvRpSJfqhk+HAy18/A9r2gu0viZ6K2/Rt/nSguDfBJBk
pU7JA2D+n5jwg21Qy0TFBrcmF412UdyAIwjId1S3GEkpkvaJHRBZZ1dvQ/5Tnvu6stYcMlBAF5kR
iX3Sa13jNulG6OqO6n4vQlsy3KP+mdh1Y0SD9/POG5ijAjNNotyuf92qKEpKIJs1vxEHwBvUf85S
DUN17YN2KR5v8+R+I7uTXZySUM3FMCun+vrbYKr7C9uF6LdTnfQBRGwDMluAUrzJOwF1NHsal6Dp
MqGmxTw8HH2ckjJ1dYS+86U6hTIEYUD3AbzuBM4V4m7zYWq2U6H9ISt2bLBhO2bScBRtnCp6umf8
XBKm8gpPsiv4UU4bO9SrSbKAwLn4Z9slXC84ym+d5Mq6CyRyQaHycKFklr1iwnIkBD0ctYxQsYZO
fD69pKPvnCN0D0Wh5SfCwm2cfn2EJy74oreJgfUVVedPyy6JQtgAHIGazOf4xyYEUS7uO/z6gZuU
YKgMiQOmbebFD9DKQRq3mpkaizsjwlOCCXTMq7kuGeJ6CrRLKL1qo3DYg1ujQQFl8+jygxSWpnaE
x1LD7Hbf+ebK7D6iQ808/pjC099G4FoQSk7FjD8C2xmoWuDW0F2jD8mSPVMwh1vgcBjadEAUzdRC
V/oh4NpA2gKGQVdCyhfFNSj6L9DTf29wdw5TBYg+NP7SnIWbC8CkLh14B8dC+XiufKMDmngsKWrp
CKOXRU4ORYndTWAIgW4J/Xo8P2DDIuJChftJYr4uJSMhHtbvqj/LSOnERYFkagS7Pqy2Iwt/gTlZ
IVOLsuXLP1+h8zqU+z9tT+1mUs2rl0OWj+OiHcPYbHR/LPhvcdjnBsWK/6qKY1FVs/sQSG9Gc+2j
4GTbMJh5b1vXDSB83WLGsnZAJ2PyGY+gCIxYk/og3wGsDUkMj6R6Ab0urnbQ/KPzeCmZRbpEMQlW
ktGnHvzrzo/dp3UELbDIcYrVsPP3CZGDdCn/lNC8yMD5fKMSjMc0754iy2GagvowWQFlxqJPw3sS
/N/wK0E8YaSmWYJf4o429jcvEybMp5dAPQG3JbJsKkL1/vKTKGCmGzbCOBzfSCiR65HmVEqt5ajN
eTkt60GK9eQhmXAtJX/GwKIwDn43umXYFuOnD65+IwD7rKO/w3W5w8GMPnhls0dKuFarqphEOfXj
6xmQRIc5fS0bMsvKs+RD5virh2kfTEfRbeBL3JV4Jy06vvQFCyN6SQPPSkJhksrIyXMJGVi1Ngj5
gI5FYRaKxHtrpyRGT5drNXtUIFbX+clJ0yl58eKJQ/9W8jS/D45mq3ZJc1IqB4ieNoIx3r+2LgBg
CjoJSJhxxgnZABbbj+pZZzd8B/eKDudZbNaRWSdo495TYpYd/nHtC94pjyYQMM5FsUWWOtIUpVgZ
isYl/JLBVP6IRnHV9p7qd8aa/yeyI/Qnzr2usZOF4YP1gWSHWfUklxHUhi5QhU0x4HygMl9KT26h
M5p/wwNnQEbYpkdma6KP0ueB6Lq57dAZkSRZnCeudpw8o7kR8LQKdgDn0EGj839XxRQNsRDBB79N
u2MNoGrz52EneOVZVd3CXBBXcTSms7FcikittQ/MfinPQTCZTZP5pvNbmIvWt6XuvEToRktnXMKk
7MHAC8zwkfa7S1Vl0y7px/wptl5ua4vJ5yjaM2EFf5c2nCTZVauf78c1K2rpjx7981/dJKY14Qpv
JhjDqypTDajOEymuWYsOUYT0vM4yV5+2cA7dEmuV5N/EYJ4ytP5YIMbkFjt7Ir1+cSEUOLyXOffT
T8e008oeo/rG2esLsrkuMsxcpsiIQAS0x9yyXJ+S3QK3+Vb0DrFD2KR+rpGzGBnUOY14x6bX//Jx
gaMZCtN8snXO+nfJs4D1LtdaSrjNr/FJVhcOPZG+Fv6xHu6CWqlQu+fwlOOYFldxygs6Wl0m5wtp
771+xtNHF6gq4pz/s/AvRL2JXMKOwcAFuk0AfMJB2WxXYte2Jco68/iaH4WLlKgSV2VovsF5nFNB
DHuckEaVUozMEXWA6d4r4q37CE0fZ5bwaegkeK77HAvyi5gr5o4DaGZzCKHS/2uY2HNKO5Dh7S/i
S8s9AYKkckT1gv4Arpq7xLXJoKgD2nJSk+ExkLPj/Wo1Zy/BaKJZN95dZZd/DiiMec6kZ28u9vRp
SvAYYC80JHbJps2MTgGYmUlj37r+BlWDwrEYWpeka7qr9AG7bYBPFbYtquEYxHWz6q/oX01jfy6s
rg/8V7jhzhTT01pqI6Sau1HrqmqfNG5T33fEEaorx2sxOiB3s00X5K/1zppPRLJDMDDGlP7ZyChT
uUj3AczCIuKvB6DZOOFQR+lcp5JXQAKwKCqhKJzCbzMU6clZQjXAgNfMPgHJ/9lx1KGdO3ziN8YE
cw5W8++w1hrTtEVnlIq/UYpBA4CH2yRp71LO0SIyIdQ0MznJ14y4kJrdCBbKW+g7+qsgj+3raq7N
IrM5AM63v/iabnE2UEKTZMDXHHo6Q+TPBq6QZdYWtc5yFenLXFBxKSVkPEIPJiang9d9jhWxXyEW
TR3W2Z9d1OSoEjoXF31113vaXuKMwGgy+SsW1NQs2BbL6jGBR5avRM12AsqyV5c08UndZr0fskp4
aAg4YA/GFZsGpI8S6LKX80n6tNDDrOC9g3lsPX9UvCfsWSNi6TGNeMJWXARE8g92qDHr3gcRv4MA
DIJhA8v+dYEHuYEpswmTjKem2ofeQAAre7CB4dPZYGDVJCVr5OwxLh8H4C2A/Q2R5rI6KZi79aRq
R0HrFm4FR5smx46S4DgKJ5TBGSVsVYUWCpH0nwNRkN2d1m7BuEZIeNs5RVqb2zB8pBmsFJ0fvTna
z+DY7f5KaTlhTLIBJoAuJzcvXleyCRoibNL0Naog440+Ab7sAA9i3RA+ULIxsj87ge+cETUR68/N
bnZw8eJCpHzNwaEJIPJKjstN9Xr5FJD4yxDFzj47E3174oTgyFvVwp8ZsobXKmqJm3FgzEtCzRHt
cQHxtQj6m9mdOczVgeSvPY6TQtgKDKKvGUB2WhItpOfKGABpqfizSHV8YQY+RgJi7G1W++ekwaVF
+CCNlFzqD0VUMs2hYekCsDVbtfvksBtxNZdBNJ5EdHb1vXyrTzQLIiQrSEgNJGf7cQc9tsGgx/p8
WqCY06GqI0o6g8YOcwfrBfw/9muj3Hjup7DXiYob41DF+hvVFqobqhur4ZntwRZ4Gc/plS3TTR3w
re2bvjoyHhthsLH4ZdLzqth+6vq4N1glWF0Al0AaqkoaxKCcn7G/Ia+ZDMdBKj85KJH80yWEijba
4rDAS7Qbm3hUXLa3x6KT8XnljHZZ3eTlbivOKnXT+Mcc9c65MLPVtqPg7t8IQ6Rpp4VbkLNsbDwK
IAiQbp+U0VEtDzMr/8kYM6icmQuxHhaZpk2fanArBv/ctINrEW3hBdmltpJBS4WN7q8/WEAihuF7
BiGCJjC2fKWggsZbY9Rc/8h/0I/YaFOE9A1jdsh2TwS4+Jg2tw+Wo5EDMszoYSJ3dsmGqfr1NE/W
/GJ8tvOrfyLad+cAisD8uzdE6HXuRHIsPGf/ljXcqXMsSZRjk9PWw7pwF7+4Gv8g9OmupIc2XkzB
22phyxsPHlKn/WUy44diGAl2U03nQbfpnROMN9RyGfi5GRtCtPC56YCjICJ195DUtMGCgmppJIH4
rfv0Nr8wRXxyFzAC7T5OLm3EhpN4yZhvXxQ5w24jyUyNnqpvbfCA8Vjofu3fivt5Bh42Rmj6cfD2
00LaUo2VVAKMxmpPna8TOldSmxfthMtK4jaWUeaWHVTtF8hXcB5ldBnJrLnVVYFltuv2HZcO48Xq
VMuna99U4aT5Z4eTaFkdZM5xVkHGpsyaOFIsN33OmlvPHfn3v8eqpTL89d4ND1ek2Rf3fQdoeSBh
CRY97zZ/6bqCDIqcZDHY3Y832xpPKjRf/5bXGgfcvFpDgLLCOd1kjBn4BBGg0m3ya0dCFUZwlgLe
X0xXRrKEevky5SaRxHFt32Jnmt/V8bbSJTxEuMze29huNL+orokKIfOGYK+T4rd0OtEU/n56UU2r
Aw4um3WWmLJrH2NAM2NLXCcQ8H6dmAlW0oftjm3lE2WjTYGRxs/yUklOWyJ0RJjw3O9OFz7mmb5f
7o5w91weEB4mSPbv7j212bRYnyoB6YuppteEuTBCFdibRvx8peXrmILHwBNMKDSX4c5yXwrX0sl7
DIwAeqW1zKA22SDU33B/wh1bKNUDjsctUK5u7lmBGyypu+Kshh0AhQqSiGNFXWodZZZhCOWQpFHM
`protect end_protected
