`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
m7zDuy+JJxqtw51eMQFXO4lHnioEC/qoAnrYEdWdpZowH403jxTIYuRLBs3MQpIcZPsPYrgjOM5V
Saf6+ffc3g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jCh2lS/YmzCxywR/PmEFM0uhK6l6Qw+0S+E7QzOGfgYVmoJ3I6jDSggek9Dfy+Pv1+yNFyUarK/L
Er/kBv5/oXrZ208XvimZ8DlY+96a7rLB0fuqHJv2dXyEEXkU5VD9Kg1aUf4eF3qtHJsWS5nzjsGo
TMOwMAxoOwf0UWvvdZs=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1NF5Rt7HJLp2G2EeOmkO6SlQOsUgXaHd7J4UxXdxiWX1nYlzMmvM0ETqpKSNisyGmMV6/1Cqnumi
AClq9MYiVGbDXj7A2btWRC0LXKzKKeoR5GIwDMAbJWzFhKxnSnnkb++799W9F9wQ3+9U53mYXPsR
2+svid6l4lzq0HVrgJiU0aQ1tfQJOSPSWfRxa5ZQ4UlW+b3Fniln9BFuXRJG0UPP9Wjf6VASH7ZN
BJhC7dZR/R37A6b9MUSHicaH4jtIE5LzDT+gA0/RS+a/WLfNR3+B+QfFjHCvGCLxgXBQFxrBgr4g
9F0ZCckcgq088inNO9Wm0tdWbdSJla4kKW+uQg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4MGK3Fsin+7pZVcXxjIn3rC4Tzs5FQ3pUWN3O+ee64gO948UUMfyB/qWGeGNEBJpWHqsvRcv0n1R
+vUmh3Q748I9g3RuEFOcXuU/yVzdXTFwb6dcyscKoSTNuIgKODJk7LDWOaG0TEmw06NcIRCxnj9r
ZfGjXvyeJg9Q9XwNzto=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bN1/jHX60ETLYLHIdo/cLvorMdcrbVH6sH4YYXEfkWVcFE6H2tl4RkHgjGoKIscb+a7NaBeceLEK
2DO2n4gTrn1YtFmBemKJw6pXFPi0iLkzl32FQQOsIbPa8mH4J0UuEdydQb6Fv8VovO12VOWq5cEo
9l1ol+vAzM6cS5xb+6IbbqDDz1bTW0le6K/etYOLmOQaKPya2GZYtcePT6sV9dmDtiZPkoSXwz4r
lzZfSoHpFGqF4TzVeYbeRbPNu5bT0fcdyq30KnajZRdbDWMF7CQkDklY9gmT+lk2bblExyCFzooX
PwiqUrOrK4P/J5Pqxlyy4j/isBFVBZqD7mVyJA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 36928)
`protect data_block
pkLb2QodNhILo65frbQcN5I2BsDdoryV2b23GzVbiRARl9sNZhOwzFCer9VDWajXQ65Hha/4lY1v
T124jW23THndrXLn/IasNSCCFKforA2pI5il1XC/0kjNbCwkncmLUhqIBRav8DvXDMTIKR4Xiob+
WoXtqd8PizuP3ZpRkkeNedQs6NkF+Dh4SZMT0Jr+FCGtYjO8K0BUUQrR2zPxL7eXD2UIzoXhjBHt
QUogMGkwLzkv1f1r6HRJbmDvUP2RdCIvJI8COTLAIwJZIORlfenLTbeF24B8Nh3EExZj9O/DiWFj
1NTMuXBM5DVKj+50H+UasQn6SaqEUEQ3g83+nlEknhfIse+tZvD1hbFQ0GiSZXwGl8B/oEUvKWCc
F8TS4WuG/oSlBNHhin8fa8NbY7wWwKA4nIgt5RUP/mGC6Cd+fUlhUsAUoa4sJ0bhDCkTvoI47fiM
DnZw1V3B4w3FAXORgbdDhtgsqBtRoXvscc/5GmN5DM3rR2uRN76HcLAgYOgl6c8I1J3jvC7NdWaZ
bCx61FNsuNYKAxgA06i9UHO2vhW2DcHVjA5Y7ZqjsrG3zttFnCwN80DMDbhxlJdCyGOMelv0ZB8B
BmYOFfDkjQafY0Qgm3dqGmThbcbASAbmQBm8R21PNNy9szYR2z/3yCK0VfRpHwUR1ptg0IQIdPBy
6phK69BJVmKkbjfvlM4AaiD5Z3+yaayNpfTzWPEcaQ8oNDgXEiX9xeWtGsMKGK8q+nj2IS1uDCaE
nuCipNSnuyBujh6dfOjzFqj9GKP02IHg1Sxf6XLo5VzWqsTUxtWCriXPVwMVKjlVWdjPgghUFkul
HCgK0wtyMX8ZnzgrkdP6mNrLcOeZ1/zFxSfbRR23LAcn7v0oV9yHl37aEfYmi4g/7R+niSlkBLrt
2F0i90Y38A0r9Vwv58y7a3ihLwqzWF66dnQbHhQ3I+W38RcvQSHe129ppDzOUF+pqlpOqRta7Blb
bSz+5IGaS+WFrzviIgu9R4BBIk7zkmin26I7U6UNbPb6lbwgi1DE7ouF+PgpkIHyrusQDayQjArI
qtff2fi7ZS540WsgAGGsMiEPSmILXIn0igFipQVgHNrux3ggusIHNpYaFG8iPMUb+/dLMyMHgyu3
Re3LC1ZgkZpxOcoMihMKKFEfuDiN9ult7aDW5rtiU41NseDFXAw6sqep+F1Cc4fvfYCYRPIOHL+G
tmchGrak4cx/rnuPVXPn5lDw8DB7hcOlTbQgl2P3kNLeJOWyaRfWgIaEkr3Gkpi4dtE1yaiTwR+l
pnEroSrAwmAAsxv39lokwB3fbdDRdX9zebhJ+Ga+It1nPVUsnyPIZBGvNiQ1dOiaLrjQWPXjlyG7
RkckqWuLiV+BzBZ00gZmQmv+wf5RgmgzvWaLCinE/my+Omm2KeCVGGQSxD2FhHMRh5e1HWZDFQuZ
Bo24wanpNEm9Stxw7TdTdqdAdFFE+lW9gXFCzCCyalZ8C+0Pm7Hc8f1L/nw1d+0+iJOQZK29UJVD
Bp2HO4Wemyg/YELjVtiD0mskUClqrezYb08zlJedgIOqgQj7XxU7bddnwHHJc7GObTuMLU9Ha7DJ
YyqmpZqFalNcwy1Qy4++sb9yx0Ur44FPRBmC665cQD2egn85/VDTM7SC6EX/M7bcatjVh2KScDIg
kFvec++dtQwhGWSbdlNHEAb9Aj0zvzxo4WNSdcdPkUTt4ypz3iDpY/y203IwGXcdaZD4fe5DTTeH
Q5+jaF+aAFaY/3pt6i//DjVlG7rvbT8OqKV3lvLkmYojcoS5rdttO4JIUQ+drxNdWNZFVMEkaroG
FJ4LapA1tf3idLgkmFL0VWus+G1WsXsoJb3n8fTmO1KB+JsonIviyulsRrAlK4nPGxMdw5uykyxQ
6U8MsLV0067NYK/yJ0OdSSaUCygiH9reutX+zis9Vz/byNLb7thlwzvE+3vU5ZE9TTXYBWuD4ssi
Q/jhLnPZv4XjlIlaTa9+PGGPP5E2+C9H3rrdKvNlJ8mDAKJ1mkSrWvfgZYMbnIoITRMyxkmPE7L/
J0el2Trh0H3cSCJvUbJwQJozYLz2kgVmstc9r0G0Nxa9YOcle3ZxydySqx1Z66BPCkTyZ8jrn7K+
Q+zHOvgK5Wll3Sj2ycArSkbofHGSHB2F8nTMOjxdMNA/PeWaYTxl8Uygp6CXth6z6SqspUehDPrd
1qVJyze7HhmEv8LJM7AFqCTgahekRRnD3Xmz7c3+uP97iXoLUoi8S+RwZg665Be8t7R+W7zvyqhg
62qD0oEjpSd6FoEF91K6w8e74Bpw9eHN9izxfxkWXMWSet+1DrMzOXME6X/KRLcj5uMCifDUCu3Y
xESvuxU0Hz0n1uY+4H09HnFZvNmO4tizMD6fwWJ13cY52RzS4JrFVY23tbPcQRYt3rLQJ5Pw7goT
XfbQPFN7OJfB5GyDAOv0J4LawJxc6Zl6cFLXCXeHYr1cQDdh5WMWYzAIRyHudNyGaFphnvhYvuWe
ZuTIDi3TI2ZbJwpNWcs04QEbDXyOE9qtKMlcyEz/r1yATGay0QgkgBIxyNIG2CElfaiQTbeETVYl
Nazvu3fv0XcPXJbR9MN6flkZRQfU62PihwpONRnsfVRzURqFqRVT3vrtE7HzPX1nQgveCx1nap9+
vxnD2CXnpoI4GwfrhBxvgZKYfiwgUaMP5Pd/djb0rbEIOiR+k1rAota1WcDI7AfEtg1dUL6AJ+Oe
4o1w7n6xy/hRwR2YOoTwMP5gWn24JTS0e8nFV5lr+0YyY0yLD+OAPA/5HB2qMhBqPQUaBNMq4HVv
biff6Yoz2ECm2RF0K6qO134VvK8EBw+MVJm6yJdtyNyjr6OMc+Bby34prAPlN4QYQveWGAH8YGMM
Qn2HssLAnowE/n2HgJ9JrX7e3syzPeTBBIvA0xJAcCw2KRnIYLA/Ns7RnaV1KW69ltOQ8AN29xJx
I+GP+Vv2CmPMwnNQH8X22SO2S9gqMY9KbPWgNvKjgOybjihnGe2o79kQFostLjZr1lwbF0Sq7GiG
SIGIgXLKfsDMRru79R80wPwp8SNATnHrlNtNRBeth3MpwVGX6o4oYM03PwG1DGLoGSUYiDcJ40cF
8ybrk15CQnaUDTt85oyFNbLIaIM5D3Gn+ZREkGRpPl6upuAAc+dXaJZLdKvxTvIjXjBgI4FMfmxK
2JfyXW7ajVpSNHMGL54wXGODEMf/sVT5mM6QdPuWC2VTkXOQbts8Nv0P56J6I/7g++5Io0AsdbIN
i6V4gxePc6M29HC8Zn6oEH6vkxRpfZVPTbSsXtBgqVXSfQ4LU6btdsZHEHT5T/Tby6AZpSLluSoT
pGYpOZgAGf9UzGlC2CbGjugekggYaCN54ISF+2gIcxQrlNrUCh/zhePCJRXbxBaaib9UFnXbMwMl
k8YJe5txGbmpn+sH3qgGhpdUr+4XW/0XudDo8wtElblIIr1zoA7rYuIPAf+JiYJ91VyeO9PhQ80L
ROByogK2ewkA1HlEiSoaVocHuWUmc9sBbAn28kzGvdtJU8v20qbVkVn2GrcnRBm8aUXb6ILoKLbD
huXm0udda1YDlVYMnOw3hIF5/R6GX16GFylxaTNtXAN+tWNn9PctvWIFATARZRQNSe6wKfDoe7BF
VIyRx2keS/A6mXK8ww5z4oTHiAUgfAImsZ6hU93iWTXGomGqAPemEUe+M9tOvnciZ2m60wmQG1pe
eVIdbI5BQBLsJEx4aYp0KJGak2ok3R2ZgfdaPiyLm7Guy7R0SqYt+GL7NBZIv2Dz9wBlAnDhjwiK
H7Tz9aZV682oBSb9zZBbIbmhpri+FbwXeH5IlU3jH3C4hQrvnFIZyelQj9kkSZfWEiXzsgkONI7a
PviZ25ShZPLqQhw4RdErUafM/txtioctjAAeZE7ozr+zlGzdbujGzTczEWZsS4boYbvSDJAeoy0i
g1XF4hlrxSOS0kIVJx3kSf1tDH3Mc7BMZbGMGXGfRwWKNAphaNUgn41kQKoY5zdlecOc78dgN1hW
SAgkNeJUb9GY+V53n97yyXB71AlHk58nlYoUeyC7WzylTO95RfdQsrpfaYOwNkvT8U0tLmmbqgJO
Q0MRzkFLyUlZXCnwbRfaaIEBPcKa9jg1JJIL0ZKSXnFpJG9Zr2v+BkKVgs/CX0qPa/pKh6Uk9iLU
Ib64AhOSgqfQJe8htmqddRPHzFJZdtG9XqS7ltxh7rlBcDPMUB/ychrs9K6vm8Pl0ydGHItdAOAY
Mt4xk1hnhDkLxNJuTabxN+eos3638OH3TvwvfSSJfEemQifErgxX6N+OF96toUclFMN2Jb7CXDR/
xngxr+5QnWhIvPeIJmjKbTW0c6mtSEqU3W3ZA2MRa9QVZsr6HdtuYuyjLaRTCrOWpvIqmFll2CT6
f6DErqhVABjn2JnMIhWSuwPbenIGbocZwbF5rB+Im+zbttGhQSoyOKk3dCQz9+SlPjHsTkfWXMQC
qgFPYwm36VH5BVb/eI7/Ve4cQYKPchNpVVNGnk49NbOA3ctBWOQEHS4rf5F8BvAsS4anVw9iYKJ6
SGgDtap0v8WHq07Lkhw0Pk1RZikmeAxjLxHjLZ26apPfvWMQge5XNkn7ARUHvQmKlDsOlNByeaNp
+EGetpiIB4RH8enHkSCqrGSZ0Z0z/9FMvdYGQdp8ua0Ae+nhWgIh2xLRZj8TRMBdQSEWEC7c8/Rr
HTUArKziixj5GJ0oOP37TZWjetXPD0hs8mk+GUsMSYsIK+g5ocIlAwXf2X2pE9E00Rc6+z7EHqat
04B2Vnq+9LRpSh2MXsFhCu9lBAaWbDGWB9rwU31/p1WxUnroHZ0I2MjLg4Ad90SLiVh3xm9egE+4
1EPY5t7eF5xdKD7vxvwYuh25wkmwSfeWuia3OQSzRMWcnBiT5kYfQeOl/IxHd0fszf9UQ8h82oGc
QJSEHZMWi6T8f/KObcibbGI89tSen1s6DsRPpdMxmKchS7TSaoWyvgowvGf0nxqnSSjq1s9a+A7O
VKCNPLCTPBKyzAT7bR7Jqs9Jj57hDHsDEQwF/H+8htT+XgOWvirb/lmBOk4GOZbkqtNJsWiRkndi
pXZVUDU2Bw6HIkjcg1EiRQbHJB6MazpviOaSW1h+RbaMN/C/MXAnz9IEghgZ13GuuRBPURL8FXWF
hGnsDuqo1vNzOghnX9gHG06TXcyz68tpM44BYNQ28+ctiOsETuKuZxvLJC+BJwE0fQK0UiklDLG4
3wcpvbBWHuowC5g8pa+F3PmIyuYexgZ291hbDpBSf2QUSGKhQD02cirjTkNZ+5mdWqsNTY3ldvfN
LX77jC8e0UcONx11JM0xpcg7JApaYH9G+V5jT5DbpvhqnaVxFz7/8UFtUBNyhRRl7ED1il3qa391
sdzUhMX7r2h2XQC0mVdfoL5YdxC4j/NL4TMo9xuPlMuvrP5hlA3aPe0g/gM622LLD84jZcjF+o0s
pNVOrC2e1U/zliUHvthYVKKnFBvneD/Aod3bDJLGD4u3cYpclrWk63YSqcftBwhVnUygUfEgQMhd
PcnYQ3o1BLhi+hdcz8fur3oWhxb7310EszBFwUq7gVKAtMpV/zUsdOLIeyPSNc/ltOb2QoYugEQr
HjSYlRPYbh+4+gPp06O2yTEzHcJZj1d8fu0Ex9BqvIX1zhhTWwq9v3xubZ86rB4ghe4tteWrhGJc
AuhZNt7up5jZL1PAgYH2k4QbEXjdsw6GneCAwrAS58U6BOnQHwkQ9ThfSpQLT3IWE6l2tSbGqs7t
VbAtRIMmvpKNulGYprwzixq/5tt3eiyR26bCeGuv1l/cYCHazSjqXhMrIjYyvBmGrAptvEKAf106
9YozKPY4mRO45PIkPxEEkGhZ7Q3H7D0ayW809iw5MADyjMwgHYn4TEoWsu7shiP2uFcg0Mr7mFjb
dX2LCNhRyJrqj05Ore+Ac5PN6BCOONqy+OPtjihhSaptxQStc7L+CHUhqomHJ2zJWv/ZS9+d8ERn
jqWYi6tvxbw9VnKVRz9rP1nMPubMGsjKlYlrCTlKIRyiJibvopgWSRSLMTTGv6BrlHlKW1NPGZ69
XgwNXayhZbPx4P25b5202YhxRaUBSqMzerR9DI26+NeH3y41JHe6MY/9AzAEpxyiwod/C0gpt6In
JoPgzn2N0LlPnEfYyH3hT8rdctE9QXdLM5A1iA1zwKD1v2n5/Bq0OBBzW0bdBzoTlKVyjnxl8MGy
IKPcX8dY16NGr1ltVZSUTqVIFB3TlpitNgsCMVsQFRbIEpD3Kn0hnbIhPcfsrXrVrm1gy+oji+pt
NfQYJsc8IkzxWYIbisZNlBiTlS+wCsSk6j+qTVPN3lVPwuJHsh7OOKKM6qTZHCorT1+iR+yUHzfe
Icfi18ubh68FufZcSiE5JqsYO6Nira6rviT7kmZR8LZWWRAsQ3G/fbEw2hbX9OUJuPQH8Jd5YEqf
kjD4hW7v9RtL7xSXRJbh6QNfTAdrWYlSuE1Uojk0Fwl3PFynYJLkVDPk210RROpSA7RZhScCTgxP
HjXNZwTI6N8Y+83DqXAGr7fNQ6Ht3mampDaHbzNoUUfOo/TgxjnkPkom9uXl9dXbHMFGAxLE9hdy
r97a9PvvJij6yAd8VeAyKJkhJcRP0fSuuDNi4MnSEtRY9A+W+nLAWGTScYdBUnkyfn+HTFTpLqHf
sgwE/2EVfmW+CH6XD28wX2VbGUPw7J+AVXx4z2p7aMeSPHJqEI34P1w3dTl8oe3MVcTBau5fEuOx
N/bQZc11l/GY1ZeI9q+bKWw8QOWWkjcD2FWCHVr/43nk31HKCuScnnBAZYYiuJEAJMUybS8PMC2B
QFo6VngsER0vS5GiLmq53ntoJdtoqLcMOF6VUg5gBrfZ2Ys1COELe0h7QVnTo0IZscWWFAfVd8zJ
3olrJwtWR/1gc0z0p52PEVFLVsrBpgJ+rQ8mBzaD4DTMnGtzFPgR8DfVgG5Zfozjnt9iBgxoiQYS
mTiM6ezRhTBPdFqHNQXPI60TuyTwvF0iHKcRKSltsKtGcFYWve60D4ycA2RfeOx9/p1ItZn9oG08
D6/3JSFaew3i1BQUe89GOGPL5fwwg2toZ8OEuSH71ZpQQVED1PVHjO+jL27po7EG/0cl49DlnecG
E26rG1yTZ7RmreJ29q3MUVgcoER/nGbzPVgtCDg0t9t6QZWoLZBZ8b/3GaFJYTIAWC7xS4AZcmDL
Zy/FQp0QjY3sxBXgqVQJyX9QwRL6aPBhvHrFGQ6TvFKRBGH83f8o/Em3Osv0bYK6RWaKlJdxQ9K7
tI06XGFp3BSonUcTr6zpvXJ9I577b858uqGgtvk/0TQiDvLvbqZyaoLRDYwdHAmifsyskrdivT1E
7rCvgVVLXgLRcG4/KmE3KNWXhAZaGX/lAJkLnhmYmDsthgEd6HpFD7RP3FErnSCklslQIhqbJNnV
al8V2EfyL0b3xnZWdQb3hG2GV1OvKXFbOcVfkHFgawFkNa4GFbCHIV+C1DFU6TmWheypapetlk4g
uFwRmJ5EarTBGwJfykB4GwX2fSETXQb6E6a1qsyMC/gDMMgnF58tiRJd4SLCtDBlUHvjOcKALzOt
hMkm9qxOyu7eOAGPb+yylf3FvkaKDak6Ov5mzeuf4ZXllug2TpANnL7sszlXmHR2/b2uPfd2DNT3
BX2YRkz7kQcmusvi00b9FkJa8u6ij95qg+fZ8pUcCsCrlO9ieKw6l5jMRKvPZ0BJRPF5LbwR8Q+r
86MMV9ssaTADSPp6n8vEmelrVNY9BGGMSwjRkyNuWXOUdUXFrk4xB7JgUih9A9IvFnWpV52Eus05
Gc0ieevYdfig9EKDqg6nfQK9kUy5eOSspgpoqS4mSBXkwyWKX03woGaDD20JpwHsJGGSb0mcAZYg
Qe6ulIFlB82ClxM2VP6EvzrD+2kCJUHmvjCjRaqRqGbDnfpd3YXXMvlNxHoDV9tTMsacCC28b2EH
+WmJLg5J6oELUco6f6neGEH16yNKIfZA3zZUv/UIOBYL3O/Zk9m4uvh4uhU0sKHjBIMxb56mhWaU
S//mSwcEipKiUAB5GRjOcmqvo7Q5xrSudo0wqC0hXkWSwsV0oe/VdEnZBYN1kbxyByzAdxDZ0vdk
Q1zb8YA5gmFMfrWs4dvFmd5TBapyfH+xBuGSrXXFRy6TcxGFO8ca+oLTLuLP7Pkdvm6BcbBAWKTq
jTqbzKE12qeh40I0mi4B4fhwgSJ7AybGdlmfnzZbFTZHUmmZoWl9rKGDAm9rdX+1C/IqVvvgeKpQ
XV+sA9LM3A3Onfuyj1lSoe6i966WKe8ICDpUMkRXexfWavr21osuS5tRhCZ7J+KX8xxkEOreIcJt
FPQGZDu4Ipxvr/XCprR6p/6wcajuqCJdlU3wM7UXnj5mC07sXwSNBZ5ereVcgI9hqEguH4ryn2cP
43nO4Ld+uC4vfHMywYuE22WS63jATizy4zbNgwZME2naMPH2mU6S8PWesQoo8RD5ngO8KEq8gD6t
Z+4uQXZnzbAoadrkS+iw/uyUt6iWO2+dDocJ3nEykqqJN+pmMlKz5vcQC1g9W38TA5SnXxtl42Kz
gv4F1SzODc7J023ZlW3fyYq51elIG03kHhIO7eELp04m4eBITa9cLQ1z3oG4ZBYxQiPorqgzDtjH
GnTqdMKJ5THW65FmwWAdE29OA0I/oQeGoCkrIeyyh65CcvKzx+OtIfXEBXcuRlWiiHIsvby6IXXD
wKiJZuBjBTtagA9+ae9LLrsp2yWwFOUQfmIfCZHnkLmvbgTiAx++EXaNCjX1CPG9/VKkrCXs5yph
vEe9B7wXo/QDiYYbDmOJAyGrMEoIAtpGZ84hl6vraKghWRFmTt8XuD6PqFwMP0s1SbbOroSo8vz0
uyaWldhQ0scn/yDqzIB/m7ansY4006yESE940GzUKaZpa9uGapC+Bz8K6SgmgvT5STpaIf1S5c4T
w7wI4c2fibg/NvVEZufFYB9wliorgty7fDjXB18LJhXDlc+p/sKdKiUr87Oo/luvNXclSjh1Sm+z
DpRjYTMhxG+cHpS3rfPLZkHEo5mxsnB3lMkdgOXdkJk0NRzYXQEE/DGQbuewEaG69EspEk0+bAdC
LmTcnvS5XhC1rwgdtid/szA07yiygzYy33JvmFoaQC6OdqFM1o9FNub7EeBE6NWAQvqqEc4WGWDF
QDdzB29x4uUjvDd6ofPp72Zdo/nKGEXhCM1BY36UrdZyvuDcT/77wrnsL8b4PryHp7W4yL9MK3/6
/GhOxzA81c2gTpYWDN9YPpdmkUyjYcaRwPlSGBbyBCtC6ATOtSkgcM/xGrhX6Wo/LfZS3drbj4Ak
uiJ7yvkA7LSOKPSPv19eh5n0a1A3hYI4P17k37F3BWtujVOBLv/7kJPezWjYFL3XMBIAMqT4Pye2
nQLBxuBkOvr3JWzca+jNkpk8bzp+vS8hgdotfALonvcdosUbwyUUHY99benKkbHjlT5++LNDRXWz
avkFOUNyynHg6kiOp2V6HWQjBKbh4pW7LzNEdluukkD4WHn32VL6K7tdtt1CoFBy0SgpUDZu/HHO
V09VKl6Z2p82fyXGtpi96vngg69H8/HK5L6z4pE+M+M4LOST+Gn9gsUkFGsxbJAs2/8145Dqip6T
rWPmEr17FatnmzN74kgxn8AQzfg8xgL9GmZx5KEzSS6JI60M821f6l0Q5mFiCqGJeMqrL+Uz39CS
ETxH5pi/qz0Ko6yyd3NHRShE1ljAQhkXPDuwGcNswbW8IAdhFHSI7Y/Aps7+65fz1niPINLQdlZU
pgaFuQqZNo3ZMYM5OKnLGmW8LvH6bBmR5v8wsJgM6Weg0Nykj4o6ysFzJ3MAjVy2BrRwCHfDgtS+
hHRbBrzKnIh4ElOoSJXr8+8BOZOoJpbBdLRrC3Z7MbxFpvEc2Pw1eW0OEyPJioF8dm1gp4LZ5QE1
b1hIIzS7u7xv7RsKgtPuBb9tJN6+K5uX+Y3xrj79ZR7sy5YxBHUpKpJ2Y4HTKua2v9Pl3u1TNCti
gkEjK+I/67q/gtf7Gu8yutUlfpVx7w8i0NznniOwUQEMbaKYiDt+FhBrAP6SwGgCmngduO9uZJKJ
cmk/1J1QQt7GCjEj4Vil68zQJeRLc2lBrt8kDubj1l0CivFn7E/iKmdegEU4oL7X3OzCIsx/mUTy
qjgvA+p4ybcqZDZZRlNUUOB9vQ71MvMVSu6HZjLNzUIoImSOj7OA1G/3qSxRjsAFwRqaMVJ1JIg6
h/P7qiTbvMxqT+835mzZtLYHywmlajxQWWLOjmNUwUXfJ9zXjrKmANH5HnR1g3Ec3D7FHNLEYpKv
wgrlcpO+cDaIHmImbo43jHmVVSHYjLgB4c7VTgULm0xBxqs4z+vltiZQ/8hZWP97SGIf7YlxWJDs
C9sT/8nRyiPLDOOn+RT3ly9eU9+UaWrS0ZvEKI9OrBcekvtbksM/Vm8WqpsJ9R+F7380jzYMtHUD
oYwMX6KWmc2XVTAFYTzoHWfu9KL4nd0lai7N0aNtFLKPN3HIcnihxTA9qlDOJjtGEaToSXKxI9uv
hDbjoVbN06672eICZKoWcr8ePXzC4XKL/LLMGL+D6dMzyX1Pd6TbTPaSt9zFbMTXakkXAk7GpSXX
A0+rX7x0prR9RfJF2K/yXYQ62IKFFo6RSjekuFsoZHDYvD9kjEKmG1TmkDNi0iJg9fT7XM22s+Gv
NokWAmtvtOAGBqloORnvyQsM9c2YbYuWIbhj0xkExR2cYsZVrhma7/oeMUdW6UgO1/DUHIXOjYGy
WyBgdXFQaxKkNsrJzaelLbLBatV1w23yctvh4Sw1C/04/rZi6FoILQ7n8UeocV0zs/2fj1VrcvM2
ILD/IJAn0R3cFNeI+5GqGB1tPO7APz9g9FteTmmx1ELetvM+XVT13bXxmU6rXeG/iA4ZxibVd6Hi
x6jsF033IPnHGRrplnqpCm8i7eKQFDvwXsb9TqSlPlFYqCTQjygTbReNMssgCMAFpPbvV2xCFa2U
U7HdvRGSkbYreJXCVA6oBUNWxYWV9tAfPm3jta/8Y7f3JuzSedbAb9wC3vPQ1AaWJPDZGlwueAVR
VP4d/BBtRrtAA1SYLZwP6e13hDMiQ+Iir3KZzs3nnUNlsav1neYvkH8MXWPeTohCk/pQuOEIsmNU
xE1QNKpbfEKRk3PeXTagFiYyaTDs6xu4C7al5u8DnhdBrBzL7hb/8anqFCPR6WKZijF25dmDEWta
8tDl9BCKO9Eq7oDRWwblIl9HgJ2zYomVgydBBC5iT4kfK+7H2rcvkvycWZZVTwhOvZW6+tg/BX8y
uxnXsH0p8mObTYwZuDtjT8aW/wjxiGUsx+syAOs4+UTGdUTqvPwuKBIa0rmNCfwAzYtvb2oUvc5m
0apyAJA3ZH6HJX0l6Hp7ttA2/7UimP/ebFVNX5q1X5WMZ/tr9lDWwfKY2DTzckkJhPECA219Mq48
gdbYhEMOHP1eu2hGXV8wQ63RFrafslEJ63e88bGVtnm1xvjH+JDuQmV8IjtEDtkL+CsUb+Q3KOvb
UxkVYi/GoLshMGUQsaGizx4oEeVYj7sj2FvkVGPSVrwLfrN0476uXobyU+AciOSLobGDd306qCDk
O2xRPpjDYRmNpqi6LL+Xv+wxdBfhWKb+S3bNyCcZ8SwdRZ+xtqIU24H15xWvPz9DoUF4ArGChJBc
v4uROKvSZ5ZTwvrEzf2mKU/qEoK84bIxvwJx4ZviLYKWNgtsLmFbew4Uew5OF2Kr3FZXcKj3PmBk
+V4FkXhULMinHX/snsCfCj/FoipcXcesAkjjYFLY8i/lBm+FDqRXhX4QjRZRETljUw0aebYhZ0Tn
mztp8sSfYukn0u/0seVRgmaOF9aXqux1sI1xSzqgLYWCpTaLG0YB/JSOFbtbwv9VW1J4zzyFQIdv
yKKeNWM/lce3tuk0nIsylzYviOxTlIYrFqJKdlE2OEc1kSWVk0f+e8j6rJN3SpcBQduT13+A9tkq
xwzNUcTfDlb+Aux6EbSWP0BvghLHi9CioTryNjBAB00ypporXl5SugLlscB64yQI/nGTWCN5eJIm
2Zs70HSIDrk8CPuhZY/EbXmHNi5WihUTYfDvymIFV0llZrCY94jvehtavYRmfKJufyjgDH9sCw6z
+7fc13L47IyT7PVSiX0wodPZn0iEpZaAubbZDRZX+pSzZZz/OpCzGDZTyZUQ95rc7MSDyaUgvCRE
vQMHaoLsyhCiSrd2oAQ+bCsJOdE2zRPKOc8GfecssnDMWbiu8UAaCVwKuOBPhcSVjuvnS0MwKMxs
MdcPM/a6pWsGTbUr9DMVjI9lHrAER4PPwn9sb2cawXi4LZ04w/GevBP2La+u04bZalRQLtFhhY6b
IvPMo4dBMq0jag/ScaGKDQ7LBZxjrZUvYdGi0zpxB30UySCUpKEobgJxJScMyv8DytWXUL1Ieuvu
m12KQcBxf9zVx7MV6/aPKIH5Ph6Ns4peT/tZlGlRRBhUQn0i5OiVBUHd+8FHGPyeoREe0PK2VDI/
hKM2DosDtJ0bppw0/lN6B7XCuiF7uIKwytRGHR5FAXBHxl1p3esLk/hpyYOCIWsrEqkWRy1tttw/
NK/4Ad+0wzp4xhJQDKtddfR1vUNaLbH5w6ARUhk/rPp727Vr0a/sWajWoh9sLNtMPeND10JWdI7Q
UffPDGlgqzxvS8kZm+tjBWQdy4Ks4vE2hNCZ+ixyDL8aW44RzV8FB5zPNhiLS0BxKPW7TIqIQpIb
NwZmcdfAk/ae2l+kb8QicPSdiPQFa1yws3WV/NXq6i6b2i+UPgDW5lVGlrTFJTxq7H5nchDhsVy5
mS2AGgkHOp3HlwfQa6WMotyJSMfp0RYv4b5Nf84Asc+dC2t4/KGKJ9A1AQcgrgWupomZ202YYvmv
BGIl74XNRpcwhMWa/m8N/i07tcQPRXV9Nqhoio7ly8P+In+S3eUPMEsDeK3HztyduJwl+N19aKpD
Hkat+1GqE6JJ1t+RsMogNcZRpFqNXDrBXykHLIwqwp8CZI7XO+FieSW71s9kP6KOR/KOwVpcNO0z
9/az/LYgBfbe6P1gYgTOXb9QeVXHJ6AeC0NCyVWJvciG/sbFgU9uHKvrpqFotl9L+ByEB2s/dj2y
1OolZhjw1k/S5zzr+Spp9hBZmY1UEeKYnjlbLhGESpj7sIuMwaVZQ/vbxmHtgpNaDgxwmndv3rH/
4G6xVUWl9rGqPmnD9sCNuwGVLBpa1swaH/+/eBEFdYoYnU6cL6eD+kEyduLOmtwrIaULtLBqc3OJ
IRevMz/5wENvZophXlKM7gGPPE/zADsnofobWuWCT2wN3zTKLy85MUgl5MT6Re3f4t1xZrx1zWM8
89P82AcPIs6bvp67hBkST0DRnTN4VA6CMRqUXq4tesXnEB69GUE1Oh8/H33NJ/y5cP5xkFbaP7lN
n9r9h6iEXnqHOCJyuLY6GgrRfc99szx7TE1/XJ78SjErU1DBQnABsQOV8ld1EIDfI8j9C5c+uClJ
V8LrsLTJARZArqt/n/p9398nm28xaToH94SLipUEk10vkxMOEZ6os1Yv/uwUqj505DkUaGMuoRlN
3KtuoTFnBlE6p0qpyWuqAMhoQf/z8ryiqpf/N+cDeAtqBsaNwdvD/Ym8gTVdzd/klQg66pTnJ4x1
VzyVmFa/cjKIbuo4f+Iq7Zx6RMpUGMu0mL7C3LFaJuE+Q5VjhTmvPUrZ6aeoVPCwEFR0LAfh9lfs
GsgODkReXA2HhLEU3STjDG7sXGnfupsMsogDVVBKCAU86xuCjwMJSzHSZhGXA0ezjaKFNgnDWVux
XzzeBRdTWPj9Rno3+EeEV2R51fMQYxRtZufns5jD+/mN8cVcgTos3pZzK9nJmymFob5OTB9w8pHc
nDnLtvz7R8Dm7rVOdn/QPgDhJTviVRrSabvjh5JzqncytbarzU3wWXpQfPI+SrVB99eoUcBap6IP
5Z5pq3OVQdiAZ/WuCxhML2AJkE8qjZ0oMu4mzZd3/guAF3bMVE5Uc696UTkqTHI7hrZ23ieHR0uF
CzZHOdjfJIviiHyH96Rmt/PNBxdiwEx+Ir9WC6+KS84lsVuzXkH21chll09hXZm+VKGWWW06pO3x
0ZDY0y2ACODFTToHud/6Rd1Yte6ECc0JGW4nRr1HUtcHZUUkFPLFgh36j14eVzbhNx3sOIAFTdRB
f4uwQ0bwRHi5uJUHbgqtSOAymYyrPVENP3Tjnxj5tss7xm9yu+9hNBwHE013KffPLeju/VVuTpKt
49eqJ9OLBxak9MAB8f3aJnl/1Kv2oVG+oME5jSalPLKgNj7Ey9GpAKzD16J48Qavd+pC9r4FUzME
5fOFmMXzn5rLZiZpzQ6buUvp0xAlfISFwOOozB2n++z6cs1FWnv8Cl/Jkhyqm4e1TdY1RlS89L1z
YruUK/GDTSFJnTeLiVkl7jhT0tg1ZIQfBvxZXNPoYZHaZW1igEOk/fM5AxysneiGtn6/0pKlv2u7
oARH2C+mTMcZ5oTqTmgbNztanVmPVzZbkuuA5ThnPCuEnE8DqBXHLE0NehU1y4V93M559ukwwMCq
catMFgYaJ/eaQ77Lu0Mg4rd0E+u1Ts7idhs2joyGKCe1aIVCYkcLATd3IXmFqauxip6rf+tPIif5
riWyvDmgRl8kWTu5gmHeC8zNzU75mYcqHqFofMo97DAcLwgDOGWMkMNkEtxf07lUoFgClsGAlvSB
de4P9EjEApxcC0vsVEy0Kq5YFhkbYEHgG98TGgYgf/E2i5uR+2PJZC1pZIT4W9336iy4jLw5xpkF
hckqDeKDGS2mECGN02UpI0uHBSUfjucvfZN/jrBmxvEBaz2VKCnQw7szar3boVPoCtjydBv47ShX
Idbkc80JAlAMS4Qw69JNnO4hLGWDNEE5L/Z7IDdSkTdZSerSh+rfAjVNhg+LSn/lQZoQbcQLcOuh
sR6LVjjdBEFdRWJNikLoTB5MLQafX6Q/FpxSNu2x7Px8qVGWmjcsmH1dOGUwyWl2fdWeeOm5LBvW
k1NnVDIsW/S9llKZDryNYtTkelbhKktR8bbUvWbhkHFUG2SWmOwFp40aElYwJ89/xGJ7hTvaKmU+
khTpNt91/aD2/tVx+AbPQYw+kwLTP4z4wWGuPcQxg8wh46HW8qaEhOX8zSNamoxJI1ELLQ784S4s
Ru9hHeWQO4pCF4W3CpRouescVTF+nIB0nBP9zN8XoWjre4m7UMsxzqajCvzdBncb6USL+Jo0MVt4
/wQlIg2d3o1CPw4gURvWBRtfp2yoUtkZWVuXIGEKz6TgZqRmRErh1FH3WNbCuQ8qeuzumdZm8PH5
nxad5jWeJjo46BxHTAZp6uJt0hDpiQHFP0aDaHX0MQ+mulswGZ0nnyQ1guZ1zek3zJxSe1gom226
jFV9FcUYC5Kq0e65rhyz54rxiepXEAtrLKZuEBX3CzZTEWRtm/pp3S7eaX175oM96QctWmIBgrnQ
m9nv3aX7rqOpe9yhZtVrnyZQ6RKhdRAJHBBN7CD2QoRdTi1rEUUDHvFntH6L3jGKjoD/eH3dtAE9
QQDHM9tuyxfFUR0ChsgCpx6JW5kKi7ijsNTZnIZrIBuJ2Uz6OgbhWXDeS5UVO5t/hNmaUO6RFCIE
0g22bYfLCR59Q6n4PCI3u4zZYH+YWEZlsLaBhY2r09NAYmLnu/eHIlmhqlmGVUTmVdxrcj/V2RpZ
aXWCfMF6hSjEXATOSVS5dMfNd0E2Skv2aJp8evuGDchrmbFefS/TF4sRt4l48mNkLrccOlAOB+Cl
7qzbwrzvHpKmZWIerH/vgpq7vf7KuhyXmjQvIirIrjgkiZBqJEIeyx/VgnOQh6eHX5MM2JtOeWjr
3j99rASu2vLzKfSQkjckjVIaaK+GCxaLvTD7GFVlNo5kQSKAham2XtzehWie2Nid5sSJiIW1lu5D
RJxwqaz4Jkav+7y/AlTrl1E/AlSdLovkUOxKqKx1odmEQVU7cg17kO0DIM0aGPtSSbS9CAg1Kcih
1i1X6SItzE3hso3gBCl3JAaldEUN89nTinJTTryGhJHrvpWX3XovWSqUUEoH1CI0V+ZVWJmS+2Zr
LnSo+FGrOFHpik/kM/GIZlSrQby3l5vmk57gkTmGn+XuT5g4GJ0Ybe+GeJuRzm4THWNEuE4H5AQc
kyICAp14bSr65z9f4oloW6M74TPFBS2M1fbmqN7Pw+X/tL4z02mHMi3Fuf+nN0rng25Ib/wI1zqB
tzD0M59pDG/64lGWMSe6wOmLFavrsuM2Lahg9/67CcQjquOA142AqU6Ko2cxvdm5qEkmf2Wnzpeg
Hir5bo+RBRC1UqdrSM0gb3cL2yF843LVfB9Z0M3qsw2d+TivEBZQm78Vv7x1GpvxNmAcwVWoLpfm
d64+Bwae70O+19cIt+lWv5rY0UgQ/lKXX6TmJWL+GWtd/EnPMfJTc0zwMQBig67/2JC7vLLF0Kdh
o2UDMTou/mJ5QbtAdjotm8GoUo9a+gSk5sEhkoYt7EAysORiNlD+Gjlup5Y4S4BoyiIxGCwYRySf
9fxDHlUfdTOPn/5UKPGwmnYhPwBwyvzCzcryN00BqkV3LBREB7rAYspZ2KBjEa6tNiFPIng9QrW6
RJ7QHlU8sKnXc6ifmm5FNHK5elKtN2gmKDinInT85FrQMIxLLqcgkU6SJtYNMlUmiolpcFndj9d3
HFdtGVCvDIdbkMUFxTOCP86/8NvEqTMcUlK9gXzZ/KHt38k9IAa2YpynWcpEhxjLGjmX73dHpROl
W45JECSzdkKN/ebH+PDmln9wzB35ET4XAsPpSfm55L8JKMKkLGjAc+SStYAN4fEWQnKjdSdU3kZd
0j1qDASH/fiUHVl1lb+cTxgiPd80hFxb3PcKMxfTdrWdzqY0bFbDwbsaKVgA7od5/69foDh+8LjD
4z634y/lJk42A/J38vS0mOWGjfbjZgbkreTERyUz4DEm8emzkjEv0ywyK7iNCJA9qcnxgpKjgKfI
MdIcIaJJLjBh/ScYVPRFW88DVtTPpdZeUnCaOQy87bo02l5VMRBGSgSdrbiTBRsiN/C8gS7aTnPo
gtiZisCeJQGBX20WvkisgXFCQMiFaJaPXzDR7C0fsDflMirbxvP5TBDQA3onaZklD/FAMdwIX22T
AcpYwHwM8/2SoOZxWT9SP54LnP+KEWKMmxp1dmqJW6AsDvgZml4Pqtg1n589rHygBi/HUkzvHcLl
RvOVtTv/7T/P0rx+PmAE4yFZWCP3G+Mo1UDkvw3r5jl4dMwPNAq8Onlte2gLd7/GKu1XUa1vCDA3
kpH+YERZNE5Bk9R1qPLjknUwARHiK/8IZvKYruLukvV5k20YuxLemmFoOZLlx/u1RMf4AtqomUNA
zlWeUyuV6KI5QijDm1QZbq8fUqBb/YXQMOpbMwph2B4751KVhraUWhj0jLjb+QRnJM9k8vOeFu/c
aznSApSR73R/4QxDoAN/fP3V9PlbQWSSAn2zyk2vyuazfrpWe4b1qxaQeCEyNdEujwnq6noGbu9/
H1g7G1ykwG/0hh+5OgI+nlhLJiR/oBc5fGXuHcxVw9rQwOKrYYIsMIm7UqlD2Ffk83mgBCB3DNg8
a2HIu7ydPuJdwn4i6pCxJo20m5kb9KiFusxFOJBG+BIkTSAyDO6ziSKXVZF93navGfdSPwcwlAf7
K2FphnBRVfSqpnIm9ZTZ+eG8NLHpggz4W5RbwC58TLkWP6HSuLIi8dYsyXBjHRS57p6I5uLXDtCY
lMjU+HuiNjHTWJXyWPA/wQj++JR0mn7SG6JbA9Qai3ro2IpPjSV8KiQhhbuhh4ZneAB+zpjH/chi
8PdnfzpG+TJHsXdzqvPt8io1+5oLnk/JkLAcCsFg98RPsRDpEVhXP0/JzFmORb2eu6SFheiRAN0l
FRzHhTF44N6cpqnq0b4Rmlojh09SI/NKTcrvVm7LkZUJ1SKBekXYv3DJen8O4NnhiJCVLh9yZjV+
FOeGp/YkFdaQ57WwJjB96EJ3GX4UqQbr8mpbgY2+W4ponicO2+OdPRrCmqvY7vQww+2iiplO9nUf
xbWHWqWNcsALgM7tZoKnz7lS8tTOcd2qfy01qWvgmhKwAFyEQk7Ep7RuOepP4nk7n4rrLLCR2ACP
RpsYp1SfvQdpDm0EUl6tRlLaRRC+sMziOMso2LVVoy+X+V+PiUDbiqYU4VMjLtSgLnNNvnnhe80O
45ZmyZqxX9NeVh5Yb8p0Dw0sQZz/fr6/8cKzOJxIlHQTksdm2aMEoJRUKjwr8gvqIE2pxzQmY+u+
T/iKj3+2ibbav2AxlPMbY6VaUmTClq5grGMMuhrU91rgcXeZ66ctAQtjuvR/UYiOhrq6VZm0kssc
WaDgGf1/JHD7qSqnZ+rZSwCJfilbE9Zqa60IvTrqUsY1WBcaxmM6D/YrzrLI0aZP10Qp0bq64FA8
llhGnrLxoZvUQVomt9HvrqXi96udbpXAAvgnCY7boHulhT2/3IwTGCZBPFiNfTRZxlM1tXcF1FJG
L2QRJzcR4W9l8MVEEZEwUqEXHvUEPnqXqZPVm9W1HzNspacHFiaEAEBQXMOHfZy5cLo9DJ9AqA7K
KvDF4s/d8tnwzaSJlfdC6GZ0/7kTDgbtCJeAf8+AKMmWrtr7yQsMq3CnKTkK4MGdqn3Zu6ApMrbp
rPh8u6qTrd8+Yp5YecWYDDgF+85YOpjUxwVPxxApkYmTDxWfUieBSxol5VxWMdhyseeekKUmIRE6
Q+34NJ8gKmc7Jt0NPGTJW3qn7TomLNYrpQaMa7AyaDm6Aa89seVtXM09MPSu2rzanCpR0IW5kRrv
yGGiR6Uee8plb0e79T9YiRM/nh1CHxbh5kV5w1cAJPysdvRC5C7RPnv2WvJqRAMgz6OizdOnXiHx
C9rIFi1/5nsb2EVfQdatZi9rAvOsxzffEfUac/FMA9eZQmzD90nZCgLHP/WXrMSBGQWZkGTsErti
zbfIhNIzqJfBHLHCeO7O57qKqUMXgbv64enbMpvZSp2sK5HeddyiOBePVz/uE9P3UpqdfaW4Gtfm
3kylTQKGnLaaGbcwq7gu4571SDtKqipAcbmrF81tWoKr2cTUww3u2jGaiQAw4dCq6ufbvGysvIpY
yw1ysN3MfiyZ3hduOKjWrnu68TNiZYVgkhQbkDjXZkcPlUttHaU+/fTRClNHkr+LJW7mf3u69jq/
Uuqjtzdrr9H3oZbvKeM4LiHI1RgBhIr04XQer6W+YjfOJtYd6nfBxkEzG2KSFxZ87UiLXB4clKpp
1ULjzE6ko1e2H4hmkzq1IEV2X2HcOVIwyme4mMHJfO2dPnR6sBEZaztYifWb2/uJC2KrLTaZCzsP
wZdj//lZd8Frk9gPI95ni6IhCWWI7IwMhC05TOBdAsPNtRSSphoY0jFIK8NScJm/93S4mvANBaB9
L0nfrzoypMZHqvBzWBn13fo8tLarRjhl3ED98DNNiyj1IK83+Wbd7d6SGCNjLd8SD2OrXmQVSQUA
fA6zD8eXheWkcsj43HswpfNavGOoUP/ahodMI+Fz86sQiY4hlWWHSQk+WMczkU2htLNlhRkrk0jY
lI2EAW0sJ/xOZKt66q4r9+H6rXfuC5M7Pti014y35D2nOPkz0L0c9MzOgFHkuhKmE+k7ex9YoWwF
NjhNUNGJDJMqq/ECR4aPuJ9/UFdOk1BGaGrYWdJW8452g1zw/q3Rg/ajMJf6C4Ap1c6h+J/B9T2D
aao3BlipycbetFM5VHl/bg+XI1xbDLTL0ae+34SvS5s2CdUWyBTjd8HsgF5E79U5GNSX6pWptNXB
940fmEGsjXG1GVu/0638FGiJQPZ/d8/A0hQI+eFB1pXi3OZ7K9LDFLiceNhfoo5wY0tG9j58TdLN
1wMuBFO8VOTrDzgVEz8k4CgYiUsXvd8z1pMkxIeXcXxhEsyhMTmDdJrYgZWOGVR8zNFFJDwQ6evn
PR2/+Rixkx2/0D45DBQ3zcFifQI/k479kLX7DsQ0D49wSszgYOMLV2PW3pt372/TUu5tD9YlxcvS
4UOC/xo6WIsh4vdUGbZl8wLgtMFvFXGAQVZAPbWFhr0Gr3/BvazADwofGG1yOwQMjejSBkWTl+zU
zdElDrpUaYAMHh9t2GYtjzx1GeXdixhrNyyj3lQtH+S+66MbGm4ABRoA8ovj+PBLKag2uk9AsZRn
vk5twWFANb0jUJNNMqnWayvDZdVYiM6D4adv+bjSDrO6xVCOpRP0Fc2VUZzlAJ8OUoLrm+S40WX5
Nsyi3j3oSNsHlLXIEa63frkh65KMKnm6FvC7MAhKdDHumMQKvsj4AOtaIz4nVAdjHlzsXuQt3Bcy
ley+VcUq224ApYYm/q87YdFpBt79znISv3c61Se7ggvc6OmLPz900k1l562GIY3Jr61VDd345WtH
aaYJIAre37/UQg9/WCLtABYzHqZ1ZYhJlQ/Yro3nG0UUFzdR9/DoLp1SRXCGe++Qdy1c15tzvkWd
PBjDlt4jjQCxIxExV740nClcNS3zBztfvWCjZ0ZHwQ2rcZ8oqRITqk+AaG4GW3hUtUvYb5hrh5h1
M1vowgZW7FBdGdO7xa0xUHQtqzHJEbodfY0ZOvAMuQrT/udgK8IFXSNzHk3WE/Aw5uKUzG8pxPvV
UVqoVvOwsQDUtxhYWhAEHWTBF0CIxQAXAp90g4jFGLAH2NHWbwpCkILtgeDJll1B2wWuuK6xCEoe
h7j6uRpHH/DINNr63YdveeFYQ0V17TB3AnVb/K4vguA/AJdJT0tBmhrFbN2srjzRkXpP6oqPnX2e
SfKgAWkS2WcOjWGUirhKHBpVijI2D1ztUOAnkpeyShy26/4kUatIghJTrgZWvw4+2cTON2liUYpG
lFDwFPdgsRTLSkNfjF89yFDMfEJqPfsTWt7+Gy12KAk8j+8+2ifIB5XhOXB9AZ2LPzSm+9g9+7K/
4pzbEwwEdlrRK0HNSceEqDL6wV1NmuzvQcstkWlCkP3ljswJppIA5oauMo/+ZtakgIdAdV1c+Vpx
i9XcQwQRncdo2GOArdQPdjsMyUMp4+pHs3Y7EY1J9krN7ouQom89JPw9R3f3WqSihJcsHv4w42n+
Xx61f4bV9o4ySNnwzXrOUAbzYWftKfjUpW8fCcng0bcoIwEjfsZKKL8u2F3AVHSyUd8TcBEGadHp
BszgV90HTZk0tuyxsZ7WgrnJHKNg/ZbGrsPg0LrEeGK3lGC5DkhnrMDgnlQwgDdOmawWrKaFSJ63
Q1PbKlfZjG2lh8lHhS3lx7PeOX6qYzex2n11WJFmV1W2zxogeArwOCAAzpTZo0xi4c0UJhilTFiY
X+qeM0cQe3FoYbhrKQEqxJRHKXAK4tb/z3ijI4scAjXRGOd3YpssVBQpMw7v+QIDpQfAqCkZ7xJR
1WFYqHelrLgeghqszxlGaJ/FOGXuH4I33SV409l2aQd8rbK+JcW7g1KC3MRUxvZeOuswFOgpkikj
0mZkBkMDQv4ydI1xBgj2etp9/oy+lt67PtjWHGVruRRdY/Rh4W9dna759Hy7dbSAHY4KuUF4EHm/
0EABUeSELOD9fVicD/AOUGSZmpKtpBk7wdgn5FovWMcqHXQUG4T3aXet/xVhXN/cjYUbK55cOIjS
F8+CD8iPBUx3Ii9npfMihdRu/VufTFljkkYe6z2Mx7LZOhR2L4ePRqRylxXEbAuhYTgbol+AENHt
cTJ2R49bnpzwlzx1AwwuzELJQ9pZiPpx22CiR3z4BkIdN5kAiW8i7NkKIJFCKegWPc5jx5cAEwTr
CrDYkjczFu302SdOCLoW1kTr/PiJgA5S8fsAtFRavDLGHYmqKW0ldmc6ael/qHcCATQQnixddJsu
dEVsOgLq241Xvgomg3UEJGAzDhQRf7RnX3FkFXzniXKrReXHNq4rAV1ol6Q2EugskQ0zWSJG6xvL
FflXvaXTem1OWvE46I2+XMij1bmeAlo3k5KhNGeqMB605s69DZ4jKsFLHRx4gWJsg3/6siiVc0G4
BkI9D9BTg/b+HzAqqmeb9vdnxOwwhc/amRUyiHdYwFYWI/X23fAvPyQ+h9Ajd3hfHrBhL+vGm9pe
my3Dd6YzWOrBnP82paK+YNsqh6LMelwNKhI77/G8JtgpIoNYo4E47XsCroe/ce16FLJWLH1V0xrq
K4BgPcqCz1Ui+TYzd6xfvW2uaEEzPiY70TBixnTODfFKuWxoyODswNsohKvNVfhoV2eTTrk3kftC
shJN0saNLRk1acAHKYDaF7BXupC7+0fZtRbIF1CnX26UD/OIfltQj3yA9FIbAqgqULF28kOi+Egl
FIMTNivbPo6ilGdVK6TKm0nkaUHNzs8KlETSP9Y8fXeazOp8G5Jzoy/fAOvRTL0hN6GoKBeIlmgX
gFzfovySvJukQjwr5xGz8pkd9b+L97Z5KFePxAZl0fB9P4cISoZIChcZBdnstqNd/4w5Xdx1+Syg
Lrv3lEyTGwdOcuvbjgjYalvzIf9ojDLCSQK7bW1v+6WwwwR2AE3MkZeIEH8oAT/VJVgQ1n6qZ6J+
96uxTK+8TAHnj3k5DymzVnwOFH94123fSXTH455N8Jof+h8jOy7okeB2YsFGEzdKjRte/s4zewKH
3Uj0lgvsl4/zedgB0cz9+wxYSRFdCB9ZRUM36ODWAbqbkC/xPnYjU+v34NOfmOmeUbCHjtLwOmHK
jPOMP2pXGhX0jdJ8nFUy3csqClEfhp9UvxW2AhGNBZDSqFchptUjcii7mBXr0toLrImqi+oVpLNE
1Kw7MB3HlMrbRUO8i3OhDAurF3ea+emqplB4P9TAEMd5WkP4jxuOgIzi+cDWcObLpmdCxQeJZeRh
XCNrFh20/deiAsm0hPvVcAAEYO9oUQrdb38/EMRq7cJYzpv8p6fpBC2A4LQcrIRgbA5xo12iq9GZ
zDSCpj5MdjESV9UXthRpl44FF6e1K++lABDs7jqJOgaKz1ZZ8VOtAjKU9qGJ2n2nsXo3CC0Rn0W9
5XO500+kKwbPZClUZJMkp8DR+ej9xLzypeQw8S0Iec9ZkZyd0u3MQsQZiIiT1yEA4VNYgRiTvzvH
JOMMaqLHC98Yfie9aHA2u/5wp8wx/cpnJnpU7z/0MXWB6LnEt1wAskMj2qEQ41L6Xkr+JAL3qT48
SBMPbmuIbwKj9QsfORWstU/I8mVweaTiGs3XXNtOl/5jzHnOarvwWL93ifNMPxOwyH+O4TmvTHlL
b/MkIymUaxTey4U+SwfPs/0LhF+XNwbz1oX1WOd/DlkDPE6IU3eQYA5btk39OCIY53qrQk399+9y
G8i6tlkcr1ixCti/GHBfp7UByzuyNZPxSC8Pj6uqCZQYB8G64fAtHrwLAHzSaCAH7eYALToEs7Vz
3XPLfzRQfDkZe+xKxmZRnIfXL+eP2g3GRwI0mN1OZ1IUp0ECsBN9/AwAQXdx+432AVUju0tKe+0D
bPE4iiI8MegOs20/Df7Hs+nKc+UjWl0zzL9HsCNpTVoKV0bpBgtURtlBPIYKnt49qnE+BNcd7IiV
zfRCc07a5Q2W8dT4NpPG/107n1Jmyr0R9n/yqno+cBMa/sjxLozE4kQ8JsgkT/datIuv3pQCtWxg
IGHXrQk2uBgkS/0h+qIr/5XZTSyv/FodryZ066jJuHo+e1UsGbAFXMUpdt7sgIXMyXD+djVtmyYL
JQiZbudJQz5Wbzoxa6ulYSV5wcDqLiPC3telCtaKrAw17uD9CR+YQb9N/MNxS8TIYgs0WKW3n38T
gfjtVtq81NI3oy7fWBdAr6JqSl6eBhDuLW3pWPakukc3wxyYjT+Rd98xjHzDp2xpX/hXNreEzfeZ
L60NAZFgig4KWmHCGM0pON1G4bAlYmj94B8YiY+5Bk+scLIpp6xgH1dZtDluGEaR2idCm0t/yv0N
5QevdyokUv5U97c98YezPZtgV99vXJVjGKs9mFTdC/eauhwhLbZzFZe1vQuuOqHlu38kLV0zLQ7P
BFtobEzBJclF0UdY763FkL26o9AYETibzoIldv5UyxCCTv4QIfmSyNMTrOQBCmtyYJYM5GIBQXQW
fsqoupA4l6QbURStN1/pg9crHcibHkt+oyvDFPmL0fwyh2exP9PyYUkHry9je+B1s6Pm/Xz68ixx
pI/miPkiztGwo8kVLiAPlz+a5d4Sar5R+nietgV378pblBYKwWd7yzP7469Zen+lhnPFKu6MhBWz
QTqz5oI8XEKPtBO0h/qWOLQEMgWNBKHft4b5z4SNgP9CqHBRfhvFdlAUShmJOL/rixruutYgRTyw
3mMPAbzZZZaHOAcVf1Ke/yzGbCpYwnws7IDMUetS1a906NhjDpDOr9PHTqpiCvR2sLF770CToa8V
NIq9UxrkiWehk2ARyiaWb1n8/p0jLKPeFxi7Js4BkD6WVfL7VtXlEJ/UKods+RVmRJhtaEKiATAQ
sNgfXmarKeF63oAtyPp6/RYjZJnWUn8D6X8hvD4Khnxochimzmson5fBgzLU+e3GClOeTYzqkvKn
QlobGC+0csA/V6S6jmWPmCdNpzoAXzYSuZ3kwg7u40wwgN0XcGLrA75tB3sH8UxM02H3B6lda4nm
6m9JUnUJNInFIeXlLwQethhdn8PcJAfP/mTTCwKghmJ9UnH1ez80bS9EiIlDoZscbia6Z165trgQ
eSQMoLgUOK81qioBvsEbUjVMK0Ir5gXEMARrfL9drYuIE6O4hWDyjWPN97UJ4f65QiGWngzLFEHP
GpLlB+qf2mhh02S1R30chiHn87Y9JUBfHyPWaJVEWQoH4fvB2KlLFrzk8jadk8km9e5/VRjE0tkL
KVTUoYqDHe37ChA0hclJy/CidDjs9xCUIx1hi3druem5URnQNDI5k2ydh5tXUJ5HCTiViGZgRjqa
r+mDwH6xhPwFR8sVegAfyjQb/Nmjss0fVYR8WBh1DXBOULk3XrdlWoldKZ7AXgyIlKhaA38XJ6hW
+33u5DMlKHbDVRx2Ilvsg++cXZNr3jeI5uZ9TJZ3ztQmVfM2ItpMAQOpJW7Kp2q8iFGsA5lMaYio
Kd2BJ5OSDx6uCou/XzUvz1Jkowrq1dkXactk0VsxfVmawunvFGedUvoIwgbHMLbPVVdwJS9q4jA4
zcyT2HHQYZOklLAZKqdszpDVLbMQ2IiT7hsI7RdeDMHRJc7Yv+zVp/g+kTaxNAZqYlP+BzIqF4yv
N5jNUwMcmNhcB+E0F5w29Y/nJSyNf42Ughi2tx7O9SURhADg3GS5k9smXaDbxV/KA2RomxYRYKgV
HDQgxtGVmCd5CgNbS/BMf9M8/K2oh4jkOqVNNu6vr+1b4l3oU1bFlu1px69tuL6lI44b+4XAkNcF
8J++4QZmhTsBMjKvDkSBzC68rJmeDi1/Qj1kV4zax/yIdl5SzU8uLgGAB1GqK0DK9LbWuoOrDCED
k/1+4+vqDWyuMPQh9XuNDVZV0FkcSuPOvDa6QZ0qXv7d0LUAcbGJylcnvoPyf0DKM5A9jCiMK6/c
KWz3I2o9yZeIw1enrDMcP06rhWdBOotcmFhCMo1MSXSDq/uCd4gcu5VcekbBqvozMZaZWYxldBMB
fscyUQiyQLa7369uduirjzUt+eSYahfhLdUhVTCaCtQYvRQxId/z7fkVl9XpegU6CJ95J2/dBr/8
jN+RkXOyxPwJCpqUW+iNbTdOLy2n/zJJu8xyVnYCY/SVp804X/NEa4egEejIyCQ9Y1CM4xtPlK8S
GNdiOoOQ+iYP8e9dKyUpOW8GQy6ypx0AQUc7/ymXcbDS4waggze/Cc8pKxeir3gI2wKso+wPRE63
6QTX1s5GlYvHS2nAk/adiT2cyJT+TDr3CQgx4Sj12Y3B4vGxPeEXciZFxV6raX7amT79Iy4t/396
Mxv31YmKoQVo3yCbCTNHph5+kUm+NwkiM+PmnggxSc5XvJGQGHH1u/0WieAUHOrhnXhyl7U79KNU
Ya2S8DCJWCNgZzF1TkdKO0FzWLm676kOQbASG+MW+DGGgECY6v+st19trqzI3Yi2yCmMSCZAWeDu
GasEzcMgBZZ0YtAPyxLVWAw5EW/IyNOZJmUl2U/tptSXgENPXF9M5SD2pGTrKk2oOYACrg+ChXq0
IzXiVx+blbFTLjBuTc7rQITOETRsy+mp7KkDD02loDbewa9bPDcLzeQMtF+TpPpXjmuZ+jvKXtJ1
Y4jqopZZSPoyXDpHveZNKOhXoYGZMb0CJRzFTGWDHhUNUnErIhuV3lxOdTzAKE1uMXJrN+hIq2Vq
pKcNnjxtqp30Y6WnzUmanB/MC0HNhPVFxRBgmeeE9dIlK2ZmApX6+FCs4lSZd/kl0QecWVOIa2x2
rndHvGrPgXm9NE+LWy09dZ6BP/p3ksKjdhvkfB/C5kxSi6yhvAUlBAtaBUgg8wZwfdamkpVIkxLH
390/WacsQcGKuUVXzuFFxWb9I2vTYcdL4IXCKH7C0go/GobRSYyhwYQcQ0lgUUgDiN9U3JzbyqBr
arrg0FXJrHYG+gFBfeQ4MlrN0ywMU8n4n4SXW1rfE/tZe/1PAZEbNoKI/OcsGgtxbd5vAHifGQgz
aEP4YUahS5rV9P9iPQUyMtzcpvbJMEcFLupoUJTRqdUw6fxav7qELzNboYin5gquoPZvTU3+GThG
Xndpmm1/+uUpeAF8a1QqR+UiGHU/sb8tePSgXC0zDKWIfERQL9wBuYu8GFZjJ3TehwqFjTDJEhgm
bi6vMV3WThVpJH9mC3YDeRM2Bf08epgHUPc3R9kPC/ssSO9kjAGGSs5PQ4nF1/YYy+Yk4u6CTgth
Nr50lmnKbAKDxvxrPSezqVOPX6UEJfHbItZfMyBA8CQ6gSKuQDqPbgj4bI15Zk5JdVn3y/XFLpDH
pngkSyL0xNynmN9Hljs4JmSoCmBubd0EoJHsaksZZRwk+gUvRCR31ueJWwCembxE1O9EBurZNEbY
tSeuszCMl4e9wvMWA4u6R5DsyUhxgXfCpmIbYu0OYzuR3osTff475vfYB8R2JFCAS8Y+O0FkstL4
Vx+B5ILeZKDbvm3oCN2nkaVDNGyTYo5+qTRs/QzsMqhfAQF1zD3VKrPhbQwlac9JlzldhqhAs6cQ
Pgqzq0n475LGv15vZpLi5sm0ArcU/SLMxoAajNdOp6Vmk1nI73umOAgQMX4NGVs7uYuT9i51gyeR
DKadcuO0y6AFRxGsAWFKCiaVXOPHrxkJCW+COy5iZSPgj08ih8bxXDa1bhepFjc8xX5hJsn7afZU
VQokAFfmQpuzaTO5B0jVTTRRviKykaYLSgl82IwnG8wGFTXpI352/8jIaHgURbf96+0HK8DV0VuU
ILw29gjW5flz4/L3SNM859eqc0YLZB90NAGcnnMb9a2vN7ZBkCFtfmVE3NyB7BEQ566FgEQ/gtH4
Cgw9ROYDRwwVu8pAhGkdY0JJ5X/E+vpuNgQSKMlgRLFttVQ/0h0ZfTAKfKpypqsG9UqOj61XrK58
eJC0gX5Lr/NQhpePMamwMA0uTtYeJw3aFJWNS7fvNs/y1Sjn//i7UdELbYbKXBSkHNyj4FfbwQvS
ru5j1/9QHHcR1VJqSGTESQu2syobzdJzBfNTj+XKsSvzXAo2vM9Gz1naH7Mzf8hq3bN/vDp0sOdN
XO/z3HXYnY2xzUMC1hve+YeniWUE7qaROov3T353wkBI7jKQPqzpBhDdXtPkso8Y+RJdxsu14xfV
vVaIqyjt4rYtxGVIU6asJjTAz8XNCC5rayj298C9kPRfL0n1X8/1cfVhohoCEjywJWouCLyKweER
/M3/6v2w2cqaiFFDDWnmwm271lLdXgk9B/NSzR4F7sH1TIxJ0v6OrRQD/Z9wZakiCaMi61bV4Mmb
1XgJsAnZ+vu396Nam8liCHVyneqz7u3hggopXjv1Nsai0Z4te4ztGLPlrmOFfWDIh7oKiszciEIM
zS+WMv1u93lRENtBDeQFgQt94wUYVEL+6gHqcIVsakxrAxOlPMP2WuAJNKp8xPD81xYMx5a6jM2L
UGuJQeh/ffUxEA+O5MOJXWOfX5djnEq043OAYu+dBDmJuFR7rywQF3lnzzWl6iV8lPvNiKNXK0c6
6DYKIk53dSDsdCsyQvpQlrI/cCJEHWTEVR2us6sYUXVcgeyqLpVS7a1rWALuF6wOtygGRUPM/gSl
VHvwefWd74oLmTU6ScVLI21UyB7fUHNsn9GpewwcA2tK0m8Lw2vbwEyLm/41dDfEh7zi51SHQdb5
skXpJrk4tpORO6BYtgnw8jA5J6B+CXGPl7okcE8yc4FXfhqWIQVUMSGEqAP3c5ktUUTHMUhEP8Xf
W8igGsfLxiT1y3Zr+R6PYY/X21Vq5u0xvARvgykHL4Bjj6AfgyR3MEIWQb3W12b7uXTJEfIE8zWb
Ni+vEU1uByytipI/Xm7o3mMXPOeKSEZIoEwQQ9GhZJM5hCv2rDMrVSN2Q35rzGov2j+LBoBlNqL/
1d1jVng4ch+F121tr/klMi7nve71Wwv11o5JRqsLXLMRhTN7D9gA/Gdzqsq0QyOiv1iXE+u1FyfX
uZFThVqFxlC50/AN1B3PQxmFiLgFoG+FfKUDTPDUdvjUxWAdO3wWEuXH7In+uW9BW3MVhj7hEv11
4AiSQzffhh/76ctePlEYLSYxU2dv+WJA/kw8ljrqtgkGnvHjdjSotTBGdTh5L1ZYMpNkkt7rbReQ
/USqZocLYJihrPjKaBXKURPk5O2X0/JqhWI46AUWwOviWCdVeNja4JuZBCJKZ/fRsnkMT1cXQvkI
xHFN9gJ4ddDU3Jyv3zKNwf5iiu+0fcahpnzLTcqDNz4TPcZEcCjPA6+u4xi4v1lju91RQL4BDjP5
q4le9B8N6f4535FfINCtgQpHeDfZy2Oad8DaV0fLPptNK4yGpPWhPbfUZMwjrE2rpKTZnRgfekt2
YQSQB8ZBVQe4odZSHYJ6etb02QIqXplebGyfvSG/AO7JW1Ae9kjuUKY5TbAaCBmbBwDy7VMoTdDC
QobC4ugdAy6dPWNyj/oHoWAMintwheV7IdhHb+qEeK2E2trkhlJOnajmkfrWYJT4J7koWFwjIO/5
gdUxW659LCN8PKuxQIHZcDfyGuU1MYlxlA5oSCioD7GkDFYj8ueQdvplehuzeyKViSd3GAyRftgc
BETslpcJG6uceog1Wxcky0X7Qv/GQnUKgbqeQOXz6qh5fwPh2B/8TnhLyfFQruUB+1FMyBYE5BD5
xeXUOph8GCXR2JmtrbKPYYu9aY1L/0sY5RhJv967l1P1z85uahb+qDpuaELY8P2Oju/RiSNjsDsJ
uve5uGS0jJq4YuiC4oEYM2+8T8Ir0FrxK6DTVVVBoL6xdUE3o6cXaZvjbQie4HjvzJcPVGZ/366a
NykMgZ9b1RKPb1LCw6LOu2j1whTNrmsEyfvhffcR6Nit2M7uAhZ/0fZdKRIiK9+k9P9QBa+ghVh/
1SBgG/hKYxia2Zeigx6MRsv3azFHEV9VgGzwGyvorUS0QLXaEDOHcdHXnY82Cz/5EzQvW3rbwVf9
aqwOIK72Ehe3X7AJ1Vq0pxgm6Yvmqpsib/0+3FUrO8AezrG6nBk3PGr8/9A1twgMkwcuhA9hYxnN
xXZmKP5cxhlqO+cbSRRoK5g5xoEW71MQnEOkDIkr37KYCZVxt6TrCj2/ksQjQOuq1TjgO7Jn6dJF
lGUejM9Z7EXfEMe72pljajkD8mdmhFhlnwlRyAmE3EIPUyfxV8yc2rLDZkYxNhpQ0MyKzA/cbXJg
3k63hJ9sI0LQorvgkjwtnR5h35YTTYvKsCpu1T+3GmvxFOWU0H0fiq42ct70MdoZvScNvd5Bn9bY
VkjOEy5tvq0Krvwd1fZT58+EMrzySlRWJPctMDi2Xy7qC/790feTjZIal83ihI/5YOq619QN6k1Y
mJt79JajkWxsnDazFgq26ANu4Y2J6fRoUauJOAJKGssxqhvH5Fzk21ajgk3RRSJyweQTiZH3Qj3h
tRRI9+8rVMdc76mxNt9aK6LV+oFpGKkneUtLsdhdG2nX59IvtywU5qw891Adyvw3MURYXwdhWCL1
6HwlB4cEynBGU0uYbjn9AkBPjF5Y1dyY5BNOaB/lGSBFXkUcc7mJlzTyHYh/Z4kwJVHWVCyz+Ka5
mrrVEsSd+o/NIuBLapni4ZntbuB2s8cVg039MzRGhrtrKFYxBE4t/RUoiyb3HZkcAnHTlX9z/gH2
jKuEV8IhOIYEDtMH+K68l4Sqr0ndeapsYQLc9CbwnlPKQ8zep1d8KrNiS1XAFLpeRuT6SyLcylgC
zOefaDfv1uiZ0usokIOqzzBToeyeYfg8vzUcXeoc1/D9Zvz2SZkTV92cJ/fzpPFfFP962bjnzEdw
ukxTJ6lTmirO6wBcz4c8gbMBQK6si9hKFs2A3RnNeVftAXSiCqEfCpE1J01cz7NrtwQX+gqPy3cP
blWLCEBA7SWhLvrEzoOC2A7qh1ILB+vtgAna7QTqQdeTTEn+bbtpMnPxhQJc1gPWdPO94dzTDW8B
GQvQc2W8dL8woLWrL1lziwlO+gR+iHi47pVgB+qG1HynwigRa56PDNqdT1eHe35HpUEjTKVPTuQR
eMxgRjGZxBbvNy7D4EglupLehbMzkUzcr9YhUq4IjCGnPZgbV0YbvLUyaFXA8uyIhCRe0sChKOsm
HojW1Z6666IK/c9Li4e9sWHbJSobWgj2pQODFrjMB/Av28Z+ZuUbTGlBIw8L8iDFTdl/Ol4ZXckD
T5z3iOraozHnqX7i5eR8MPmrjx0MHbEkgQFAEPMZjbMxORtECPOsuVFOX7WvFX3sONiqgbHmMeg2
0zq4Z2hABNLMJT/xfh093EVHImgLUbRqgxE1z+YU4u0gzKHJSVsMlFKewfIPiszxbkcxKWTyrRYO
GIeTAFWNb1fViDBp4NCICC9IhXjHWEnooqzirckvZRdbtJ9LP9jmuzodPXt+TbXk1pa4upIKUKvl
56HSpxzM5aH7yVc2C+/88/jFvmADMove1wgMkDEftasHN8O+mtTXIkmJZ+krgaOTDHsveWU409sS
mIdMVC3+AtlcBP2Jb0FBH18V2fQdEIVLtEJST50hoi2oloinnmivopVa9UDUH8z5i9BnCiXUeUjG
sTplVk01dEmaEFZ9fYOY5cNLcO6d+a3IwT2SNXPu/pZ/7mtlLo77ZDbUkymnQZ89WVKL2oLJzvk1
mOjuC1U1qCsXxv6Wf4P5gfQl1+3UEvuBXlao3sFa9rryfk3oecV1y0cqFLhqhg2rzgSOgaE7on2J
DOF+qwggCKcVKkU2ns2YVkDGmVtOo1Eh3seRaYecsd0wsnzgkW6zH7QnZCHoBxnI44uEqQkiiZYc
x1PkjXMRTNocAuXSat26smhdZEyM3dDWBd9BVxP6EuxQVh8b/dP6iJA2JevMJpxACEfWOTSco6or
moa7IQ0xFyO5nLIU+pMed72v5h4NfjQV1h7DhYI9u6lyLP/gOQRCM5l77J1HxX3lawbhM/BXEdTq
LVczsWl7axm0S+yArcLmwu/W6lRWXx8TF7YPbmvXbeNEjrD8MhIIiJWQzfGhSIA2tfxjBUUwzGOY
ZiFI7LtAXjOPWBxt7qpKxD/h5trDvU+QZ4vtcEhp7uBpnhLxl75qu/HNAogUJsZt4siY0e87aNn2
OXAefuEZp/mzuLKK2jMOJgjvIktRL7ptwuZ1ze9FSt2Q3FHa/dBx8VdDisI8ELjyj8eAyISAVAoD
B/o10In5lh43/TDsvAc7H9NSXsPA0NvXXWk1voEAxvOFzCZe+TDRU3zoIF0Wb1j7gHkx8vYS0a2d
ah6jIcKGbP49lAdTdAh3aCRpNoYGJVFbxLoPwCxCYf1kaBKJjnfHGuoPiSV3plQlHxf2KGm7zTOj
R2n5FfmxZRmnSaTGk92DDshRGDyXxvJGnSaxL9WQZ3HCPgjofIOc0e754EAJQ7MMU1G3aIWO+UE9
T+GWlCIIpT/HANYlTA5/A96OzthsdA+0kYMyK97WtD/5rwWCQ9EjZ6ONfihPGfgiIKJgZXerFEFs
8ChZQdk072HMjefe6aKYGy0/w1qGAbBWC6zZYQewjW5WSMS/0WX7NEwCgu3gej15JKjhS3TbrWzy
JXw482W0noG541o7Y2qytvYJliCLhENTkOU3vwMQx5lzOjHxCePVmxushumIh5VvbvshoblfN3V8
4Xe/4Yk/W8RW7yNWTUBJVZgu2JH+PGl7h9689Q/3VX5QfTffUS2Ges2KQoUMkmh2UxUUG65Nb2WH
MQnLlvXzfu8WqWRjxu8CvENNlGjcp3/nONJe21XFA3KnqZX+6XF/Vv+SEqpmuoXO4pIpVaXsHvH3
Lv9vFzdSV2N4IDr3rw9xv96hG3XoqLMdv7KBbpN3BjwIu6Bk8rpfHpsgE9w11sneIQBU2qeGKL1W
QNQpmaCgBo4G6wlnTrGtjBp9hAhFOgp9NjzsGcD0zd40rVkw7+AsPG8dF4V19tSt1OSmI2/wHPop
avttuZfYXb9XLJ3V2+Q25dHPX7QIRzYbPKC+KeXzACoh9WY7zl3nfeUBtDvudCO25r0IYW7f/cKk
5xyQIMvpJDknWT3ueJK1oAx+kRLWZvmjknJ/UyWeZLkan6GkqzkrahlqX9lKJEz0hevvXy2O8gIh
pCWL1NwGddfP3ZRBXYj5oC+7bIWTyV0O0l9V/iBmBbVntOn2ZlDddSSlhVria5MKg4CnSpjPFGwl
YKaxk1Bl9c1CtrrRwyuTYNoOlcFSgXwy+awsems6ryKaLjyWJ51lpO4tcsuHSAUmyq2v5ZxnHskA
T6dVbuQtk1HPzN0++Wj81aQLS9dE1aJX7VjHbR5JMRZJ76NYa88AU7McvxYIvjxvso6jQL4kAO3E
Z9Eec0jjdPoAR7kpW2Oz+7W3RxZtM3Z4qZpokUjSjlk+zxqDbz5p1WLCF8u+buoDlyQ6SRMG/uQM
IhKwruwzsOPPEl6Ej+Sfp5lrXf04NY2M45Z5nKNeGadZ9ae9X3VEo415i7fmJ+LLbFIOkHskKX45
YUWp0pIZ1GOr/nnLfwN/sQTjV51gJvTzlqbjSL920oCXUBbnmLTMkRQPDEtP4a9owLOpI7UAG9sv
09x8XJmBNB9Ix/2vWedNt6V691TJV04LgrvjFpNDTCZwKQX6aVli5vJn5ZzYFf21uJQtoBaGdYXe
DOcP0e+KenKETlOamzY6Dk3RYat9cOU2d60Vv+If3MYVH+6wFPNTDgCauDATeJpzXpQC1QQqiy4W
BDPAQR3JkyXWZ3wP0Oau9YfeqB75cE7/uMT7rfOA2jq02m3X6I4djunx2ipl7ygf52kWE0zobEez
LhMPBUU/igj4pT060UJ7+Dmj/726R4+bIaDIYwLxhPOvvYkoYENLz62ILo9ealwovweTu+QnZztp
DvHNIifmNRtht0VzW91OVB+jv7gej8WDOu0oyxr93jvrmiVh8U6SfFmPJ0qczyIEfVIdeZCiixtk
XbZ1M7My3lq/TMzWA5HeG0s5pOYlArSTzhd5AEOTLn+rzX+j+aPZlsWxkv+2hu/fl2rzEonol4St
FCbo6rCIECNHle5dtmHTFuymM1XnbqaKF2ogQWzQacLcXixM9Fe/TYOebcpzCXwf88e4oS9hpeor
TMZhptZpD8MHaWuaM9N8OZBWnmx1VANNHJZTH9lO2svblKGmnKwNU95RhQr1Y6g5hFmZBG2KlJ3I
Yr8h3Du4OwYni20juktmS1YkbnzAznw6EnLyBFUxb7Vx60BPnyPNR5kXmKB3Htlp4m+cT2HD8XEc
MzvvK0VrgA7IVmLMVY+LPFqKD+blNCyjeHgAZ3STUfLkRaa+CckCo4IBqAKw0WSbW7IXLpdHkUsk
f/L5xjazXi+T5jzcHJ956pw/fOKt+0i4d85ZL0tprIgn6Je3yp5U33lyZ2H/P4M+kAUTBNxgHh7H
pHf7IaQKSyCO+LTlsgINev+3oiA/UWfU2phfL8bWZ+UTL2mqIjk8+vDnTb3q+czg/H7EmbO6q+9a
SaGiIjoi/kS+OPIlVZVdbIg0dIbpYgPyTvAnIc6E0te3Ve4hCtSPvW2+Imn+JkQQeoi0tjGtlGEq
cpJ7uYdODEPBWfAekYbk/GGeFEkLs/LtySO7vvW7NUmnWzvUvssnhTKNdd3OX4QOGxl0fDAYjr9Y
PaVCYD9LJuH1Do5nLKMwCBO1/Z0OVTPW1Lr+6Ttanj/tV5XB0U7e/OXmF1iVbO8oGmqWardrlihc
2VHLQb3YIv9jqdiUDb2p8D3/yBRfki4kxzsZ1zBDsFlsWnmP9lGuRzTB7dMtWbkiD8RDR8zxtA3n
kyP8qw2R8OdtIVY0rAh9bTxkVSWK/9fn3wlGyEGOBmgv9kA5kH5jF+ku0Il25d/Sc6heUOH43M/7
FG6heeFMH5mfRRFYVbdFRudolnYTc2n2FIYdu83H3//du4y1/50+zQVnnhs1ZlDyUm7utRQ+dNN+
QW35fID3QXXO8Tp4kUdz6sA0TyTMuL4MGQzGn2K8Ed/eU/dJNuCND+YO5znjuO1zpVTkrFi09p3O
b2IcdGqWvJ88vQaeyTAwnkF3Juwkh9JEurvRRgDmN4FXEZPsGKmGLwhZ18vnPHjmRKvezgCCzgp9
vePfRCGxPzfoUIxyQ4E8Xv4tjuEEu4+tCiIS6RYNYsKz+7flJXwUphQwatkhvuVFYPEE6P+rDPUq
boGXnfTTinY8N/tXG+Qvj4UcGtKAr9YUJhF07nWe/KZg3x1RrGBwEejx0lbWY9aqZaFfR+twHfFM
2lav1a2sVD1jyXDru7zTk4ZwHPCiqYS0LO9oBRUW0lq0pfWyRQoQ+FPKmBMSDpYItupI2u4f/1Xc
zR1NCcpDVRfdNyz3aJfe/Q5Xhm0yidvnduA6taEoKhHQdmpq5Drl9HrYz7QKDqBWJccn/giZizjK
OFrZYv6AB4GOmJEac7BP6hdsmFOEyRgTjiJaypBys/+TBvw7aCPxVgIy6+9MhfAqjQkv03bJJoUT
xuNP7qOtf/Hq+wrYNrPjHcwTdX1dpatRY2H7lC+whSCNSp2irzhva/JBrd8gJHuqPdMw4V9VW3GI
ate9/xxtI4VLnJENXCQD29ylyYZQ7ZtQkdaNPxzUI55FI4xlwT1M6JsJf3RmJsSWVX0Bfe6716um
eVlJIRxcJajIc9VFucgKnCJz74DOCeES/NMYcyQTs/e8WBFpXr1p6RZvcXwCw6E4DvWj1nd5w3pb
hsi38CvodN4Hz0Kw5/ajMwVHCKcEsDGD6uZ2aLEzdW4/5LddnbFtUGG/tqOT1oQZpl1qme8VXpUn
I82zrHgGzCVJkUevJkJ8TaGVaZVQ4c8s2WW4Z2fklT59j6LAGPYNF974EKOJJL+BWdVcefYh9Lsi
Z5eroxy6HxJU3w39aNmXmf+PCaSZx+GuyKVyUWaWolLFWKxjGT7rez5OZe+u8+tWHKo+CnVUG3Bg
h/VT8wWNCJZKmaKF4xQpUpkL0w935c8kQPjZPZZiSSolKM/Zd8XRQqxNOFZVwTTOYdPE7DQhQ6Xf
UlR9khoBhJZu1T0+LxFRdoeVB51Sd1hl1tpCgdPkTUaGV6yDmOcPgxOhZ9smgWezV9SS/eZ+2zAx
NbjCyfZfLf7hkpn6HYly/ZzJrBwaZxQaHdqDrOp1dcVQo9Wy8+Xt6W5ot+aB4KjqzK2KZgN+DtfS
ZRX/lonTb3xqn2XFLdYcubf84y74eX7yiXnkADTb3sA2JrdCGNnrb5imdvinIbm6Dju6GswrMjUI
99Xo4ZHGq/8nf+uIlmBGcDiQ/07Ji1oHz80uLNwrvqbB929oC33XlDuqKFsnwFEpqjMpnckgI0ic
fF38WvuBqwc1ncOc3S6vQnwEUQ3hK8njI+Xy3U2DuY8ssLnA3oRiYBKs90QRZVmOWICK+IweDxVL
HVJmAlesE4tMBxY0W5aB6uaoJmA9Yyc+66GSagIfuXTC3K+rEVSrW37mfppuCAqEy1AU2qcGubsW
hlLDawUdMx6j7b7YUKmcCkh0P+yG5fhIe5yxKQSky2obK+f7PUYUo9CdiNQI7IGFOnYfarsehIpp
a83IVuyq8iB29xyI+6ZxoBAlRkR9tIuwPKQKxbwu4FUoAYkT/KAEto3AiQRhv0lQ+pj71/TxFu56
YoXh5rKU3SKsG4IRTNKAJjp61H/2QxzwjC2wnYH1Anu1SYAqjCcJC0diJglPJA+8Ehc5vLxz4dT3
+y89+O9RLdPufwtnaqgs3A/4y/uoHfg0IgKP/K9PNEXytreEH+cVocsnMPsX4gYk+X2cTsxOyfWF
YgufAgbJVujCIr4Lo6Tdigf7DKieLKIqrp/dzod6nPpHAF/uKJEWncTzaiTf1qX5d2CND2r9sTJ5
Lwqd8b93warohUHA9VgtpwR8bsFzQAzO3ezLkWE+nTyGFcMDXDgkefWw5mGD6WVSC71v1ZLbhPls
gmrmwcxGwzCwPIlOyYh2bEI4pwY642zA4v2f7eJ3aye5gFtRV04zwD00C7wo3uWDRt6yjsszXoGU
Ae5E99uRvMgMUcCJk0Ux8DZ3tsAALbLSwxPPkwplCIDFL8RnnIlSEK9Upod4f/+vq8ZUoKto/sEE
vSnZ0HC/rO//UWakT77Z5BTd/1yzNH5iqoNyZsiQiodUaafXlhpF8uGwYHbEkpf13BIVcawAv4jG
JiojJemRd7Ox6d5kOwoTFO5fgA26836PnTiCx01Ct+5pWxDbnLxye8m69jvJG5k3u1SrEtHns1sY
ibJ4xhX3Bu1Z5/7w1bL3fayPdm0xZB9Me51IvNjMOuK3nlLkcZaHlEL4lkFGZgZTRb2ROgxgr2g3
Hm9t2VstoyjhphNFWR+8FfOEEck3Kjdkd3ZFTQYzpILDVCLBHoIs/8CklEbp+MEnHsP1yjmUJWVz
UouAQdB6SSC8Y+4rMyiGzvGY2PQNQpByMiWr+bgcDtiLIe7zoj+o7xd4FUqCdUTauJqfNzWXyvUz
rlGGlk0OyoNK1ynXAOyf0/gUVMnOxGqs6Hu+YQPIIMYsWD5NBeQaj/OS7pbJP6NetsVZwl4DQDuq
4mNgea1sN6Ge2JABAT1MFy7gQpHFJP93TxWpDmye6Dlxct75uGHGF/PB5/tP9bS8+B8F4PWR5w/m
3JfaPD549iYW5L1Mge9nldk617/1sjmHr6jWeWyXkDd8EA5Gf7r4ztkQALI9T0u9YYnuS1o76oM6
01SQtOywweFto0NrUK3aSwxKaEwv+vdUIyNb9v03wMXc1CjrQ+L2M4Q5kK0ymr/HZTZbyPtGI9nn
yFKpeb3TOeKlvvj4VBK9n5kqTQEwwH2XUQVWBTFtDeq1CgA1i5BNxL99hi0CQNYf1KhjDrvuhkbr
lz630sh75ZlUdswJzZLSLLuyrC8c20rx4CMyEs9EM4bQUBu3ZwyGlDkw5DPGhiSZaw3NbkUwM+KT
oYZGoGK4Xj0SeCIMyqivtdAUzhqHowXgfas9qd6yJCPqGKaZeRIyg5Ex3B6OO2hZftu+yGBuWmmL
eT34+q+eHQLtm00uhpPaVeYqqvX2COlCVKDwwknW/Rt+1PVh1Cw/kqoQ+V+BLVrpo25/jcAOKDvP
ShSXXz9AMcpJgeO4B5Pg1HnRXEGmTryIzc14JJRc0HkCZwexQdXyO+SIJCV7elTLfHx9WBIfd+lj
MpxK9nSlz4gyUSEsy6c+AaDqBarwH4D0+hhy/JJSlu82vns4npkuTmth4tqs7Xdo/l3sqOoMlCK0
a0mxuzowNQJ8z/fGcrJmmh8IZsMmlLw1X4Pe5nXeIp1tb5nASkoU7JexpL1WlilDc7i6R+BNS6er
q6+RllXGJWEowOvuRomYSJA9SrkHoy/SzR/4l/k9ByUaoHUmIWtuHQlCPMnP/VXTGW2gff56Tqcy
ln7JW7CiXHWvL9en9d6gjyvF0nyS6GjMA/FJzOfUC9S1fyu1wVE81CsneXgyWsUOn+DVWdw0hbld
IBM///ICKuxuYyeTev4QkZ5LxIaQpGhB8znY+UUu2Jf1a19b1AMaMG0YhghOypdgkbmDm2SZCmJ9
Aa3ReUIZ139oQepbtT+jWpKDnTE8pnRz1TlRIgPtFGTVIYfaE3TC42Qgbl3bGMx2Uee2QnQN79Sw
fcVL2yw+zxjtEbxcpHbfF3efsP6nIOpk30GpbYuwhHvFvYpucyfG6Q5KyhfdxUw8G74ODQlxCZLx
Y0pHbyRsLei3f1j1McXgTeTmbW003kFVyaoeFM2qzFTaocqruxebyGHKo5yhq/Gp9rqfL7nlRsq2
cQzDPkbAmJrf/T2WXMYHBIwGjsGs38h8k0V9ehVgNROW1GsNEKmU6+rsxJrn3snGX0cr7HJDYiMd
vVQOvl4cO6ieW16bpdzD6mhoYOizpgY5az4nOTsf/nqnopNjlLr3Fx6EVccrr5kIogOxsBvZu+Yu
zkOJaZOSohO/WQS36sfYNmW/LoxuxMyplGPKOWHELeurHD9tVBAJmnEjYLhH0ORfGyZLae73HdnD
toJ2dzOLvmGZKI6CDYkkkkR1oQcLLxxh39Ff9F5kWETF+sjHCCHNH01zfJYzWJ+iagWG+DcmOE9t
Ee3vOQrVvDrZy7udetnSATY45EcRv8P0kdGQP3lMyJMS79cJXw5hxO/fn7u4/E6yluZ+U7RWp/9a
ZjBVFGMd1zaQ7L3VZwwI6O2nxoVIN31AZcgNBJoBz5XPAmsXPDDt8s/3QnUplF4H9bBVdfXBhru9
Yb9xnK5bzJN4TH4Z8bekLxmzj3sxElhoHBVylwhS3aNTuYquYN47ELDWxgoZi5l1DTBYp1u8sQmF
VRwh87Brp7wiUePE5VV6GkqXE3wEDyXSfJMbkqa58u6sDGqvYgdGis6xMqijQJPiVW5+wBMIW78L
10nkFaqWmPcDyX/Uxefw4G/o8wXoH4CFgJynYseNNFsCNOGL926SpcMwExIjjk606orIfjbq7UuG
5UKGjxSQKPA1V1tVkBdQd74ahjvJxEQX8HBWvX5aj2bJbgkGUIURg6Y3xrI62VejuAgD2vc/Kqkv
kFZYqQOj6AyCLr3TgvZc7Wk8wcQVuuh4c7oDnUMDdbZt0tYbz1v4EmJtggP2iD2npvDUG3APVt7t
jh3ytr62Ih4PPYFm0Jm/2bYE4+czKF+bj7rjJAebKi2NXArDb5WP0OCss1iRIwXsx/URpVMWSgtT
Nc+3DYY074dimBfJgtHG4RYhMQiwFz03c9LXzUkGHZdSBhaJTK1ZODnyO40SeFpQQW4Nv9ZF06be
sGN7GX9CzrACgLSd1GH8fe/tuR5PRpxsjQpPKX662s8ZmUqyHryC/wb6N7/H1Zq3XO9VRjNQTIHo
QgIK4JyiIFEw2hwBcpqZVb/oSJdNIU0bGnWmnRV+Zm7kykumUNQgU7qpC4XrgVAQPbyM43+ivZq8
AOo2tDmZHGrvBhfA8dMv49mEBXWrItJ9+sh91ir9LXUukD63GT3xvmZ/ZBNJu/o2rXDvw9awb+++
q8k9awOmKadnHgLfqjbmwOnz7LIzdMo7pXAQs9lgjJclImU2WV4QJ46J4nFwSnzEuxOE/eZddfmh
fcw6wMEyz9Lf0F8cXDw9PoblsKE3QRlJSnre9spPfkbL+8f+l8OkNSpQVTkOlI/pXOWYLmmfsg7S
stCwTQo5dZtzAt5Bp4VjscGIB3es0jK7MZx84Lf1lZZTJxemJu59WWyf9QSX7PFNl7ffbWovGhtw
gXWqC+UsRhkdTbThF3IqunhFB7loFC+K+9+YjkDhHdh5FQ+NvXkPiMu7HrA2gXRVkvJ8KHNi8Rq7
WELMrsExQYCCp3EQ9XmoEQYJCu0urkRcmIxWrY2sBBuBeR1SYRb0xkouFygwCTA89cwvYffAwz/l
PS0Rqx5tRmvYj8+RvmujCX6BBQP3bw7a+qGMHeg5kN795tYJ+wOplQ+1QZGVVVpWkYhNesFAzdJw
Ms0IrlJ7AyrjuSuHOzaTamENWUfbZExv3hbPFoBPYZabhhMzLNE5qKkDHB6B1DVrMSFhhsvbU7YP
YZ6eXyaQPXVmEEZJUA1P5B6wwtwf/9OaKsZX4YU3mcBiU9lsdoaZDW21HlGtNZFNbH3SB0amj31H
BtWgMUk20JKckpfl7zxDQ7a7+YRZg37MHLcDTtsScuocYIJnmIa6UGTZAhTF1J0360kMhmGDiaYb
4RYG6dLXqKy/MaRBi8wqw8PUrga0G8tnC7kQ7NXn2WMMY7wTHfplygFJFypI9LLVubxOcgHW9EH2
7QiorwBoPxd8ETb+htADEx8oBoFpxkV4QIPEl+MbSV+eQq+nEPQzFyp0SVtxhnaDIkfi2fOMOUIY
RNPmpy41RUyflVluTUJ67iD/OW2nv4BYYYCnigFcXBhp8yfLkIWRE9fZI7YH0MBj8Qt/3DCN5tuH
rLWgLG+U9A36OGjTpFd98zd8B0lEa/ya1IcvfMl911uRjYZ1cHVxY3cDILnH89LJL+fxZmjKpATl
3zh5OChUP2CHJo+VRlD2TkIIM92fPLmp1WC0/baSKOjw5Y/KWG4z2JiFByq7jUeIVUQenqNCtlAN
0on+oJrdw7bvjgQuMn5E1RGvE3arbDgGjr3lW81F49+60H1jKpycb6njojN8OgTE3d8CaEAwyoib
C64aqwuozOr+514TlTMQW/hZZ4O1gRKK+RqnWmEthciGxWyweJYq9kTTsh4kzWCM/s0b0qOU6JnM
Dk/VdjnLBx6odzR7dkK5tGWxhSfoIjo5G7A9Cw3Q8F6F6RqowwoPPtrMxYAOIhFaZ610XIeAyyue
vgOYQJEq2ikeBVP50XRRSr84yOlgJGDH2rLNPsK8QyOav0Jlhn8QoT4rBQcAlwgmmSyrhd+oaYwp
nVry1IGdmSXEuI0JBHfl+cC7RxLBi2iInkTrQhOU1TyyaD/b91vn2FlbNkrfl136pXj2p49zvxIV
h2pVsgPvVA0jlnyNSvnKZrZXNj6mnbgZTAEokx/aX3WTlP2BxIDLpddg5gwJnp06SHZq4XJ2c876
11YZNeeEzeFAMnNsWnvVu586kbI1fXpuK2KFxVuBcutwvN8ZFz5VSkyA2Ai3AOdLIS8lZYZGBgYq
6GOjFhwNWTaL7kIF1XtnFDWVznYjLeky7UGalOZcQVvkb6p4Tnsu3N5Xb5xvgrk2Fs5BGTHmaP5G
/QKzbnIoIqBOTyrgaNrOx6fMC/zx4atYbVRFyhDv4WVJTyzN0Y6Io3x2TAWXMB4V6OnGi9JxMVld
NB/JOnQQLCrMvfutjUJq6D0CYE5ViXP8WTVCFyuDb2VFePdQ263/jbgAGD8u9jmYwN2Zpjnv8MsI
yqvEIEjdGojuizspQ6BN3a7WHgfYava3tHL76gqf5TLYgV41ol00+BwXPpp+CGqcL8FtM8UuuRrf
uyzoDvc5FUbfW/PO4lmGfn5CZF7EOku1C4OzEMID9NXfmG/Qwtm2v6kUxgRuu3kdugrat3weVdQ+
1PHuPMjBQ7CI9gUSF1ox9TqA2MMoQUQSLUrdMolBMF+2XMYwDGiPcIn1tfZwNSFNeagZhYPjKizp
6vbT/bPZaD2uWD62nFd3oAdRet9naGRyU1edyty7yOaNI4n6CmXggjaw7LRp4ovr+k2dzSLvZgLw
aDTu0QMBC3MXZxiEz5JzgMC6mwezwEoF41g7fGICDMr36yBnKQaFtkr8Ncb9hAO1c/JqJlAjE2wC
XirNmQReYuCYp1Fo8uCALeVEtZvfVY52blysQrkTKKQ5ZRSVekMavBDp8vT0GsROZ9r07iJk8wm3
Ab9lg0iKCO/UVugvNaci6UKnlXMCbXOaNY3THK9IDna18nGttFUHTkjTMpQVkUrp2dzQwM60P7qD
krLvHw7dTWkvmczvs7sjde9kJaimq+lPXdRl+AFlMDEMlZBCkdz9XoStWPTx5TxkSVdwDh2U3N4o
SGUyWY1dnPOkZFia3b/3m8u//t10H7XKb4ogAjPu79JTY8GfKSsq8Iia8iM1v9i5tcaMOhqBL2Fy
XX+V2f+MUlRJnzz3FRcd502AwjlOFqlXKocb2PTpb0ljB4YFLUi64c2Z/uBJ5rFdujVB52r1zFU7
GUrkyebdpA04HpAGM7fTZgmR3KC35v4sIZxHO6Yunr/fM/JDTPSmM14aEBNG5xZ5tpmzrq/XpxPY
wO9bBA9MebHwZGMBVGx7/j47Y8wQT7/Zzd3HKi+UTGTnaIH2YaDGuzpJ3bGmNrIzsjFaQzsM9w8K
1m2i8OMXVIaGy3TvCZuNBqwPSHWCfBZi3Xu61HgPsM7vkrR6vpBIgCoSAfPvsq3VB8c+LXM8U65G
zKEyembqFiSa0+jmwVOUikHdXLQXqM/8pCumGBcctBi1bxpuZ6xoi3FK7SLqj/ifYZG/pmR8GQCY
SAEH7Y7H5djdqWlDFmHRsRetYZKE/iZJoz1je5Do04x9kqW+5I+gs4FsM2JUphk8VxaDgikHmtNf
FosgaXRsJup5XRwBJtLxoIytNPOqKrx3SINCsfepJ2TWd4283/kEvHhKXoZxyPeIiqxEEkLL3OwF
lroiS8h14qWNhg55hEHs/h2UKmYOWFzjQNtohUrqm2PTUDXpgQctiZJrjU6m/nulFbXmCWqg+X6P
hoduAIIx/3M8UObqdPXZHQt/l0GctJu+UJLNPZGO1sdyv9bVzdleMdtWOWEGypOzQRhdAOBx3FrW
4+W8URVS0cr4yJ1DGmPEygy9HEmNxrj6OhmLDY0fTjQPStTuE5fYeVIVgu7JOpWmw/vpwOs/wWtP
BrNXeqOBQW5qAbq/7xp3HCg+dejqFsJjFF2ig4L/b1oG3PryQOZlfZMzaqhtoFLQz15QxVul8Ukb
S/S+V6XTqhCg8MgrJ2MceZ/R+O5YELIGc9TB8SxFSNKsGXPMMEGrWz293Dxfy7pEaVvFY8RpEN1I
vpV82I8jgNs1Ze6w3pMDnMSl1cC7JHTqUng88xeC28M8X4UULTrCNFEhJaqlcpUSSC1m7eINl11Y
lDHEPN6st7oOkO5w4dUUpBMj9PPJ8KVYY/IRFtbeT1qDkfmvyQhipyVJ8OsztFcSioeBJdI4Y0OM
n82jJISJeEmWRQpTo2+hS7su+FkkFGlBogvv/p+fYLFkE2qmuJ1bRMQ8/abwQGI2oqc/cPG0IPoP
6DJkn8YdJK2gaCvUoaeqp3sI0iVfePxf0EzcByW7lnlqnq45VTq/W1edAK4sYiCOTM5nqSngeh4e
HzpAYu7ek7UeTr4r21k4x/XhIcsXleJdzO9kHIgm25h4Uekrs1H/E1r0J8t8jMu45N5kD/qnbGq6
BclFNiD4hnmz6P2LMvcFRloeoMaN89y3ZOzuPmH7gtYRMyQNs0VW8qqjUdK/j4T0Ff4OWiwzyMAF
GJ81wxHY6SzJbe86aFYBsxBlWU17jDQJlL2Aa3is5+K/2zV8A28N89pRR5UnLTHzTwzU/OYwpSpK
n3KyuaAMBjSyyb17XbQO31FvoRZ1g94pG0MmSxk4ZuLHO+bLfdCyN0vaY7keZWzbeh/sjqHrhHmp
cz0lSihc2P69eOZ3qni28qYCx9efM/nZvYs/8ZqWisIR5p4aGH4/7QQBD2GtMgWyFmfLXc2hVdpv
XXZtOPZpLBEPxtU6PHs5HjsaDW6YvWbhpatlgyP0+SIOKrfNCDCLZjQS8NBA4K6ZVojh/g2yYGKM
rfrilyHLviuwkPIqQ9oMVS9LmdrVsJ5IgIK/TWaLS/gNUL94UeIQFQA6j3mHc7f+aqaRkmZFifyy
NBJa6jIiTfnkUr109ztX2jm0p0Pee09STkutevFUvEI503beTSB6EXufgbLOPdlEetItgnXmPFu6
We71ruKky13TQF1ctbqGA0gzBnXWuwOT7E9VoazjZ6zSYDqvE1TBxdRj8brpjB1AvUcApww7AWf3
Z3V+KgdRVWffCrOLDLSlX/b+z13y3iiPzopPTX9s4B8zB6WZV8yOt3YfR939PsoNkcC+TUGhuzh6
9ayclb/gUMuYSnz/hRBb9byOQ8z29NnHvsFPYyX6Jx5ZkqFWGgtFQZWpewi4KoGSohjsKXj0lKLh
MVT3Z2auojqM03Bycb/SAOeRCGBFd/mN+mWg70WY/b4GGUlqq61m+BGzCD51INEqawWvKBY/W6yY
kAtgCsAtjksjyXrXhREy+2fSiFTtl4T0PaXRuES8m1ure7ehacXMQ7QMF9PVbhIoYrOpASke3Jiz
UqBeeCMufi7Hl9HEsm6pkzvTjqxx6XsA+jJfEANWtRd6sYEa+T6ig3DhkVkNWPX/P2Px4Fu5S6ZZ
mgoDgDyqRTn7KWOoIki1ja4L+hH7ljhxTpFZxA8qBXr1K6LGOeh3TxIhHspul0k4lfRdL/+znMIo
T5jWMQUb4Pjp77rsGmBzK9A4I1EMLzued/T6yi8JEGQif0NKS8BbAKtxzh8KJ1ud8hTu4Kzb6iYN
S6xjD3pio0OpdRYIJ/Tok3uugJNNiMlyjTmydg2PlH0+zypa55f07xK2lhEwsbGOK4Nfr3KtXAsf
4pvzOja0WwFdYf48mQ0zHBvB76NKK1cX+wEfa/jzCqV1sTBSf5OpUKAcT7kTsTDKd1oLQNju3D2U
m2pcCGF8myJUqJtH1veQtMFYAj58To23VuJSLN2clf2Brc001gr4QIAvhTehByEenQK7PAcBa2to
3giYP2grhmxjUwv8h/g6St4+1y+gOw4wnZx0hfuGj1LkFNvjwtruIucLKtzCY9BP3FS1NKZVxYQn
jvjLLO2xG7PLgVMHE+MYVfIkgDUMRUOYO/C8owGtuwXZwP0Wt8J60kkWGOOXWGAlarCPl83pUtVv
dDY4n3uNJ+0YXaziH9Ync8+R6rAt2zN9pKIykxnQDQFJrYaMlfF4eGS33S1aZRXGFShbWT2uzWFq
f4os7ChtY3Rm5eYO9Xo67561bxEHUxV6pJsgSLf+7Fe6Q6aSMzfPvtcU2YpRhZl//FDtcPfaKcMb
5k2c9nFBGb+OMS3YWk6vBv9gVPiEWa5jSEVMCR9xwr6qMhh1/i7rXLOjzhUOzVdY5rJ7uEUIrhXx
PxMrVfYRHeVjTi9gtjj5Zu32qV+wAs/b+HfAltOGf8XzcDWFOLSBy01DmX4IhqT2BTaKaHydo4bR
69qpT/UqLjJvXzAsCpCmEmJ+T/B/3LPfB0hBikQcuaC3afB6MoCFfaQPQiDXIEkspVv/eB7cjam2
H8B9rrfo+uJ68p95W3hqjjpgOsCLH6Eht7WVjl8dEVQdadQFk0XPWK2MJ35/gBiplh/N//TrZXIf
/pn52d4jmHlPE24LHN/9J3ZMe3ShDsrlisBA1OT3LB6E4DJiuL3PaVCzZy6KsbWZ5twCo9jSrxma
SfhF5eWfxHMsh4h/gth6SvftqKgx+kG0YoEM6jzFFaKeYfqrZsNjmrODtq6LEsezCRakdX1hSWoG
MuIa45KmSVtr0Jz15TQq/eSQJlEo1nabndGLV18Vwo91HG6duutGtPcwBX3Ru9oAOHf++Z3SK9Z3
narlSk2EzCAzCmiD049NN5Yjfoh/WsKwRb7grW2fWmN1JwTM2eGjA2ooilhnP2YjKLr8NAlbNTYD
YEt5USwOHIBgpCG7AsSmiVmkq7gB7eN6n++s5vnjOvEJFbuHyEso6My8IoxtbJEdhny7c0RM64+Y
doijor/i2e+C9Yu8ZR1hTZRGzfiX+tQwybT5c8fZkdMmo4YmcqKjT1uiyjj/lIlrJA5EGhB9NJr1
ZsDuY3m3BOSkSwh5HUbH67IcGQrkbB/WyRVLIlwAjuDxiFY3aNyQb0doNixYBTEwEohJ+/f0Lv5Y
SvE32VdA0HeKaiULHvgE1oC67lOxU1k3tHCLqUuxCY0WWZIXnc/MvJiFhYOu7GbL21OOOh8hWJv3
rTYcBnCWih/f+BgqIF8kXedC3eRLTdxs56eE66GF5NhJtQ8fbLS/ujnZWXcif31Cewi00qPM8HiW
QEh6GzLES1mrm23jTs7hNTVg8FYp85AlGNBCXvWN1CAeqbvidZpanLS1+t2DWeSH5fCCr4eZvxgW
6sCwn0mxYtQmex+t9fsR7v0trqhudok1TTxyyZf3nZDj7nfHFLtRClmiO75lo+MBA5klUb37mdDl
A6sHLGR1b5ogdQGoctqrrKqv53VsbyMURHwHL/qofODFnWhqZe6VroxQ/BMVFU4iS8QW0TkGdVv7
tzsx0kBE+bNmCo7ZL+ZqwpSMLrvusJSiP9Z7I4yFTLUcd+y6HtpuX7XqcyIdHdli2K+jnQwAFFWO
6nwI/krSkZa0nbFNS2hb4hABAxf9B3S39YeXP2ps/Btr8yDpzzinsxbW0U/8LZ1w56jbxwmg2hl2
5O2A2/FEOWue6lS/KhnB/MNWIU8pLl1CycH2MbaAX/fGooaxKZWAYsB99gdbm1h4bScApwM2Snl3
8V5MIOMk+fqSYD3xV5krU5HGLFv8ViGXQEA0iEK2A7v9mZWyiEcfNf1gQrDn1NBjJiCAgWz9Ow1j
X85zmi9e3KaMNnOsY7zOHSY4iDVwc2UoQxUDKmvWfZqHPd8KmDx9K3YP8EM/+0epxE/FHvk72KvZ
TI9VDUQtpE53ORpA/rWGXbE3vh6MLr3YxaY3G5g4h63j/XyfN3PFmYhSZNKbFMBlEwD+UThPbgrn
BjJ2U01Sxujcl04BL3k4PS9/NjqLEOIKlQQPs7GbBU2LOMDiAZw+9pecW9SSVGbhtlb9PxeoOmKW
eozY87gU6COzBT3AhefL7J1f0Dl7Mv23wB6pMkF5AoLwZTadKrERgWqLZvRmvS6f++Slze8D5+ho
CWKoCF/ctVqTP20XcxwPkiIYnOFNnki88cqz4ZEvS+DDOGVRSJZhdD3cXRkBsNHjlN7aibZpnkm+
hV3mQuBtpYC+aYqjCtXaSycou3ZtHq6Iro4/4O5v3ay2KuaW1+W//jagzCz9AXvxLLCQGlKbN5v+
YcJ8dWe2QW7nAhWTxKeuG1tbZUGYZ2BYY+++AB3EAtahAPQZX+jajxRZQfnlf0GkNUGmG22Qn8Pd
ESqCtwMjgpGGRc65JSoT6/tZqwzriZH9DPWzk8Tcd7BpVRaLjiXvXFk0JhAnZRe48F0RowqUnJR4
Jr1wVwV3f5g2tLu9lQMcftr+pgQqyAzVsMgk3rz353EzXFWsrbbmPerUGO8cVUYrcR2H4I5YGnwR
riFFc7G4s6rV1R7zkQQeMan/YdkVmelzlxJ38XNd/D9D2Lx4Wu1C9NhaQ36UqmlVXhdqHuk6spUC
C1WKaxhzjJ+yo7LrnNveYyeXzDjzDKH0r164na9ho0cdaz9R8fxQ22n1fkolUPpyo8vbrX5HdIoT
lD+6dn/jaq8NR6mBpTNHxMmMD0S6THVgC31l28Vf3DDMAobH6kezq+Cw5kH+c9VsgMEpIpoj5RMB
eKSEksh+jQMX6NHaNocz+MMXiw86ORP5x6Xfakl4Q//Ves2Fd+IwT0HOxslsO/R8mg8nY71eDlvm
Z/FcytR1cI5xsOKJLxS7TCivRAr7qzQSAziU8OkfQ0OGqx9RVgoWNitGCY+3Pq4kxDs+VusHt7v5
WXtWluE1ShZcfxy7Ml9tqiu+YEUw1/eQLu3WgFElqNeR+wJ02RVyPlp6NrI+iAURqtVGc4PC8rpa
EjQmMZDx78s3ssLFvDDmVGUEmuAh0eQD/Wm5Aq767jvocryJpaZKOewtCD88qUa67R+6tYzjeztt
95S7VjFpiQ3xWoPrOqCGwbw4ohj1Yxe0KPUHVBVGofxRLzJYaGBuQ//KzvCsaCMT+M5KfR6x2kww
le5iVDRMtL5l4u3s9q3N3jPF97m26sprmtEKxTbBGD//Xxavwn1Ebl3Ad5XvB8hNokQK2i1sL+Ju
Tm8d+CtkVN4C1Rx5IMMHCPVx6BY19KkCqYxmSttG8y0AryzdQeAH+ryKRg2wW8q+i67gnol+vFVd
SnK15OZO/R298+ZL18qUtXzucKLJJe6650GmlzV/8LYsWdJhP0ee+l0GaNg2n5R7k9efxl0gOMuX
fi1HX+LEiWO4OCN3hCuPr4t2NeV9Vi6hPABRmaipYij5Sp24ijJYSxmOB5Tk1Q5WmqEWEVJvpiKq
qPbGYk8z5TdsAfc/HtSKTOjklGMGOe/LtTF9WUMHGUcwM08HnQewrJzvmDLFhtP5xS22bd6ukf/v
qh41VgypQtum7wLs2g41NCReDUvFnzECyQlmQswLWnAXKibNr3XCjgyUIsG1nd3j1vTzpj+JXcIs
7QTbir/YOYpI1ZZJMM/1p8rvF6a6rqKWd3rPDMzdtFWtk2kXErZbCrCFZIpQaU8s/JPSTsRo0Xhn
vmG6H9wzsz9FDq2VtbxMH38buyN2UAxlbHLi0lG8ZQjFaCv5Gu1W92EkcA2i8X/Aun3YmI7FDlYn
yWXS1ChxhpC6xdFxnLiL6mfXmFWDIyK1gEZqwMZQ/A79j4U9sizuPpUYy8qSK2W5nt6yInNW9etK
ebtQEzurPu0zmMJiLf3iHzdoF58+Jx/Mr1J09TU0FZN/iIygV7vgeKurGyFXZCUxj0FonK6zZKZf
0ewa19q5VxLcMvFbr4dAsU5eLIagrzrUle8G4QduhV7fHUNkeZnhmvKgxVfqli5qBAllFrg6jSLB
JfhTcCkrRWfMV5PLyWheExkykQZbSGrgRw/WncgbCsdKd/Pbp/pmR+Vcn5/2qRu/28dKge/j7PUP
0A4QK+4mi4c4Gaq2g7fW5bt2uwJc2m8ZZP7igZ1z/3tB3uhYGHxPX6eSXKMudHvg/Byt2C3HQtZL
qw37bqKIBOrYPCjCi0948TyBEkWpSEetJFmNHjL/LSE5UYt6elQgU04Y0qZ1p7EH5pj0uWKCcN/P
avhqKe9Yb3+Tk1Hq9Yx9anBSl4t4ddyMIJ6seES5EBdWz7Ga/rPerBwmWKP2TWbuNxjUv+e5ntfL
Q7/szgBJY2z7NVU6eIANNGM4W3XHa3RS3paPHdqSUmIO94+GDIVBwRFKW/EUZeduQwHobtJhZHNT
ebi142MhuSRZh0k6hWCuc3s7ZCdUZ6IzhSfkBD6p/XZY5qnzBVIrjZ065qfVIy71J7UqRcPJNHXU
wIKgjtDYCYxAsd63CrnYFhc92jhH1G7Zz5deCYlDJHp3CTvZPPETH29ru7fGK8UWiH8wMIjNgNea
EzMsmqfuhtbyrwJbteboeSMgayOTPH1FbhTaUmCK33/B2FGsQQKbzxHlGB+gwnGaXg==
`protect end_protected
