`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
itDJtG0nokOq+g5nZrt4q+F5Fy1Jemg4B6ey5i7F2FSeRYIPxILw+cFbsNviBXCjRO8lnY/3ULdr
i3uhMZHpTA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YJjlSwgasd6BkfJHKMvMRUwDBAusvpvUTWraoWtVSFID8URvpErs3RbJmLB5WxxpE/NcL8BwAYXt
tw09fxV17qMMD43oHl/sMQwTs/GUnqVpu9Yxy/hb9GTc3OuGJEW9Znrrh49lIIwSBUoAMzzLAxM9
8e4d6zGJATYD3lKdOVo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VItk4hdRXCAgy9JXpOWrI9hN458Jwtr0Sikxd+eECOXTHHpE2VKWodHMQB8v2krzwXkRuLizrgbI
U3GCQvqmr8TH4h2rgPzn7lXYADEkScMVedBjSbQrOI8rK6XL84fzULpov9aTlN1KRQmYzr8MkmRM
2VQyVTDYGR6lAwGjkdsRfQID7C5mp52temuGxoEVNgEocbP4q3FoZcms4qopwPLnfJq0ZJ7V/20v
rAGjWrPMJAb8TrzRcwhG5BlEm5HTJ8ZIeHONrKiJQejO+wsxYDCEVILH32bXRSvPnBPtXwudBziF
jaZ9/ap3bvurh2y1Y9yqtcp6f4l88MMBuoiA1w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ecoOvbn9tBAbS2crOl8xDHi6UsvPsq6QscC3BEr6llFvgwir8cPVxJa3nydCM43gDiTFC2ingt3B
fridbBAZsY6OWvrWSzlbrEJdpZ6w7SkI9PkiLwExYro0q741BiQXPQPmD1UyeBYiAPMHCCj3pr4x
NoAKjDgbDgGxWaA+vNk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IzvNZMQv5Ip/yTU4Nc6mulDml17D6lz/h4ra+0imPNCGv9Pj9HdmqxgtFNAF8ezWaypOcJZ2kExg
uPEVQfPvPRI117t26+CFoXZZ56R2aOlZvA0J74aZ5irfMZH+1zS26C4WF8J+QCIevXO5LqPcpbYo
OqhkgLZ27wGNRviOg6XmasAxKezUtwkDUWYvTrtjq2e9mfTAJRbCYPXHP1JUYPQ1JpMOPUDQaJ/9
/xj3gtmtvFcSlAqxmsfoyfP+lShLyuVnEcNJgIV7y+z4735mrlo2M9zyp2tvlnZzs1ZHUzc3KsyC
Jx41P/DBWf2L/ETFRNTWlRugVfWyCnPLd9EJOQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3248)
`protect data_block
Oce6+72E+2OIv4tK3R7ogAwQnU32i7WidTtvJ+hHgCaYyFSF188GEcfFCJkwTJn35n3MCYjGhTJY
JQjjJvTSmLmBidiRFSTOzygbQG0ahylwNgw6Dh3DTi5lTfWHVlCxGkmqYcY9z+A34x5/VFeB1Dt2
Z22V+ZrfbVEQXnAaTDtIzhEn0IBKkyP7KMUDc9Y1exaVeUs5AfIwpL4XBgG9KN0BlUzeE8gzMEg6
Gek4zOBNwi8Sh0PWkpYzv6vOdE4vCVc6cXH94hWvnTAWcD5b8bNDQa3Wj6MfSY/2eZQEaVpU17u3
Gzg7aigpS7zmAtNqkZGoZvtrESNDLR1/YZbohHdRsf5LtUduyvqGUPVM1Q4naNpDxEKPx1W3zuE+
q8gGNuF3xaCXdoP+qne0CEg1w/k7N9FZC6ajEHJCljjdQKB4JPyfH0khe+eBt4Hb1YXaX+iu3f+Z
t/y6w44yxt0fqrF90bO5MAJ2MQc/wrXZwc24TGvdmCjGLFunKc9YggeKx+X7uMDSQa67TBz7YtTb
X9lzd8uNCiES/gFY4k6NgMyDyGh/x8X43O7ubfyatr9FU8PMTzUVf+cMdo9qwzJSKZWPFgpZGONf
WSpZKtUmQf+GbKayDcReHIQ1RlCWnTk58k1ZoR34lh3r/C2ih8akCtPmK42xOKP/IeCkA1KlSsfP
n4172Q5T07kH4eaGKN9m1qEY0nZozKYc0jUaT1ev972cknzw0G7/yqM3Kn2a78+m8o66xwAZMIJz
oI3Aao5LqQR1OjPtmRtMC13NCLqDK89JOnhk79ziFyyER8seUBVvM7fKeHmabHiV2XYy3a9Q4sBD
6//5vY8og7e9VSLt3o2Ls/Fg996S7xT+kqy5/MsjlKSisfqV9PAjEbXBN8ItzraCJieq+fPILJTZ
KPeH4Q6Brv/P8YnbbutvtHNiHYGx2dgShhilcUUMjSsPncGmoam/hgMuU73Wy21PnHPtmxjDxn22
b5CaAGRMIzNcbieSq8jWjY9HgqD6G9mcm3ZujDjI8/4Pceph6tIppJVwaNroW7s21GprVuvLD/aT
fDRoA/CdlkkCN3Czx5Aq9oRNla430oYnv2nbh0ETUoqwrOQ8R2G4X3iNA2Ngx3o3rvrSuNwkWX5N
kXpjNWn62xuaypFMO6dSqUwjaO4Rt//HxhiwQgV8XVQnRrXSToileBJckkMS4WyeuhAGSdf+oHEB
GiOcifALtzTuVgab6+HGMxZXImLDABW0nl+8NJrO3Xx2kRcqltd9Z46fXy0HTFegtqsv/esL9e5C
FzE130D8G2KOsNXA7w6pRHX5TzM/eEp14EFwS/Uqf7RtbrZx9EpYghe8YevLD4XIPvfEOxUs3Hrf
PzrOYyuKx0N/81/xO/3vr/lRBFlTly5C2ULTpTfm6D6SJTUToAB6byK7s2Rt1aXcmNXEILI7YyY8
T7TUMyvY3QI/knGk8MYSr4Wlk/wluwf32Pd6WrF2Be+dh+IWK5TUFaD/bCw4+RQ8tkz8yCdDJfG3
/WbbjY2lqFxa1pSGA1IlUFNQAy808ejHqlqJtd/nUADcYoqgEtfrVANrYd76RHXwYAT7J9Bn3BHt
6/0auqRx+F9nw4trkrhb7SPrPrr2vvpDleksQkZ0tv3C0Vm0ispjZ2IeWz/PPWclcyv2y3XBuwKR
eXmOPyy/u9gtRB8B/H9m4ZbhCknDfsiUcVdb8TBu6nx2wHNBFX2mCHXI2GFmjWUkOdcRRu0Bikqm
kkBax2jdAqhsz68bJLRfTED5+N2iQEuclt96512Srj7etlmhlspejV50jOkPBoZOnmwneCCoJ/OR
dvysWMALH/SFG8+9yKMBSVWLpB7MAHZ8lS5mtNM4Lh5ywDkOgEsjWmhMIgvniZW4iwAylE4qmWf3
h0Kx5cYmaWSzy8Ya2uQLISHZYL2q/4JhP8rF7JOfmaBGfp6UFNu4cP+HITlndgbhd/3IJG/qNt0r
BAHi15HTU1nDbAfUAIpvFkKDtElphubqMMkPaqVLo82hMF9sIh4MHHK+saroOOEor6Sg/Wr4Kp1V
TU7CvfNcxlSpzDByiYNNyp30KRbBloO48IQhOsunnwyokuUHj7wPzrARykJLkD80CRbRf3zFQP7p
R+Iu4T9GmCwTmlwepYzXsxf+tz9K4s6eUYSQo9HNxyvHhEUdrDWa1T7AGuamviMmp0VIwuq2mKJK
driRpxE+6GfQz9PYhqx8D4UjQs/GenwlpPYnENE/GWknDS1dGHab7SxUCYmQxU70ej+dUYiK0GKT
Wom1+g/dN+yq39T+veQijOdb+QwJp8dRqVaoLIhvTKuP7gbhVWwZJBtn36kPu0W94AplcfCvz7US
0kS1Yi7HKs+OL7aGhNChdI84b6CU/jVH70UMyNeZ8V7+lm3R3pHzcR/x2kOLV6W7KYfCarHfw93d
BBtInk26ZzjQ8U0yoiYzRxrEZtCM+1g9n1Ik4vnpOWKJfFWfN8IGWqDlfLu54ml/XYLCxZkv6132
B8GBXSkaOfURbriAsMfIBRWowbUUj5bLg1O8MeNoSpO1HSTxWf5HpdgozX4rysFofGg40ndTDgRZ
un/MMT+zdqPiZRgLeE1cdmJ8ltRpZkRfQy5UKWlpeZEzkCZhGv6Z0S1Ui4KQ2oMWFCWiX5ZqBsKE
fyxCvZ0+Xmbni6vuwfFxIqUoS8aa3lpNkU47VLUTY0YFBUWLJmM1yyiRa5zvH1z3Wx/tpMUR5fMO
WGT8/VK3/zUuWkcamnaF1E8DZOAj+sJqewgB86bte0fqdlJW47y2J5p4dzj4q1Jki+FAfWPQbNT/
nrvyoCcaMCGvg5AtkZ6czyFR+PNuVE61zjCh9vIGqEvrsjarKVdWbxO78lbPxuD3MZUJ+N0pneRw
aMAz88K6CfUpB3uDkl/kSRtdIuxNsnoJr3Nbi7HNCrBKU70XMfH1oMEnaqxASccvDbgRSKNKqJKW
x/LS/fvEv6v4PiNlIn5lLurcfUErnl86BEUh61mENgrxTx5qfBiFay8qRLbsSTpVHVNBAOkWjawn
DVAVRAted0Q7cnW68DSqI4sjtm4peIq66uajV32JQs0D6inO1liCIGm33+6eVh+bkK+EXkCqRdOl
fcojzuaB6AIATVEGPiLVPw5S+23gdFGgsRdk76Rm8k2HOS1hXh6dNMXsuTMc9lu27xZzFLVt9EZb
1OgDQ8TcnFttX1nkoPM7EP3UXd6uJlvAp3htu4kDb6r9wRdf+qSgUOUt715GO+VbY6Fl7Js4+A06
tadUtiC6brQh2th4Gv/NorOOPEE9wHCeaWyC9+doG42vs85f7K1FboB2lIhqdBtk5m21xBJvFEr1
yjEJ7bLMR/pwbZhVQeE4KeHjQ1iIswBTSS05iwziUIKTC9COesdjzbpRn+XItzLaNbxSBwsjXYH1
ly/3cw+0052CtPoLX/LhMbggpKDVRzTpKRECgqrXqZd94rYceTHoQC4e/F8OzpySKYGmo5g8WBqv
COsQ94GEXVdasyt8vm1gApSqQklzbJ4sf1mtDEdOYwXWcsHw5plDNutc4MRMixsNFcB+b23gkC6b
6dw9uCbgzxmrSMcbdpFv+NgZ3BOj4hLLZ7o0aPDi+FhZxXPyyXPPQGixiLhgffjDOtk8B3ZAPfs9
bSxfJ6X9D8fMBrCRIU5MKXH+aTl3BRS/TKNT1D70XD1rpcZzPnEVWF5znZtOl8Yf0OK9kCPxPqdn
wp+pz5kC7himH+UNADZA+TAGuMAZhhQvZ+ywvA8ht3/zX1ebEbLVOeSHcHajjodLVOEWljrJhR13
BlPy07OYBXtNH1v31g/eymAQmpMCspgpsrrsOZ743LrmbUvwTBTBSFcl6pEiJA9uRq5LzH35FRmI
R4dzPRFuJymSkwetOZ0/LBDIsUc4M0Yz8dsJdJ15xCoFqogWX1xp/usI4SyuA1aXjeImJ4iHQcc4
AG0+TkGMhkeOLjiJbJTt0ld4FQCdomtumgEjveLhySCD2m5+PRZstmFSXQ3PDaslR8SYzm96GuWR
dKOXPXrRwVz2teY6OB88gi8lRk6gcQ0Lf2C/7ipWp0FIRP4CRh1tYvi9SS7ovahvaYZbg2HP7pJ7
mA8nZUKmqsH7housBdcMkgO5CBVieicCbwVYq/EChbjAYofp9r969cfdIM4Terpkbn9NE4RR94ow
xpJ+ovCBxiQdWkq930ixnUy675kYKdkYECaTt/g+RkZNOHKSNXKotC+xRwUEyvfjnsH124vaEWko
/2td90oezUg1FoaYqtQnBgFg+c0M/fZc6px9IaljCNaIlFw9J57yNZClmVK/7aBUz7k0PyOz/rs=
`protect end_protected
