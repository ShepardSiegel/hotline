`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WC9+6XJPw4YwDhmkAcl5rvV3mCDpkR5yp1q/3wOtRSPNteVHb3zTr/huVK0/lN/nduiKy6hIDi+m
CpHKukBSNQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lyr1RqADVdyooL0LRheuGz5ATptU7yo1VAhK6JQze59YYfIdFtIWnc09+IT0xjtTL0NEvveXMEPc
8iJtX1UlnHpi5psalGcimxqmdull1U09dKba6l1xEDRWqz62UBvykQGBkKcezaz+VsP7RYqUPCN7
+X27zkzw4opJTmFeZao=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aeB1YXqYJEG4WhSirqyUw0OaYFf515k0os2/mZ1thqosCMHMx9J7hzL2+MYPmrmAVXFw+U5c9P65
2mZcYgZ3nHrvcuiRBKAMf1QlqDy1RGif4Cl0qAygzCMDh8UJluzaWle1Re+IFAVxHYDp+zsBVDfH
ncdl0LXNTTw1q0dffmYei0JWWgiG+y2iH6ZvbgEH5ux3/tZx0yQjy99unY3sNRswSYwlMQf90bki
WeXw/9LnL/EdCGNsp+vhaVyryVU12Bb26AymNK9qigoN83QzOgnS9k6TiM0Cw+NdcPEvoByHYRbp
moblQ2eqOVJczBv2gWNU43JP1wvd67MxjpuFaQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EF4yjahengpCmtd2GxsHZvtfEfFevamVBWFuL7mrX7ww3o+l3KK6fTCuCx6IEWGFBTN2NXUICzXN
vtGpWEQV+oaT5aSNMB3qSX8iBc7w4QX3Mpl4fSbkmqaOnOTey259N3U2Q0720t7M95PRgBGQESwi
mpmXrqJXFQNloe300r8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tnqGB9q1p9Oua15rUXC752ntwLskXSTqkYwYjoSOe4zdMpy66VDiXKU3oGXTHHkSUM+30GQmyqgn
FZnJ1LWbkAya6Io4C2wKJhCHZWwAt2xxdELs+kow6uAsRUsCrI64uR2TXNAx6ewnrnlKmochX1hh
Mkt9Ys8HomwgDWfVpuZb99mAbdcgK9lJywTaCLekF7RKVvgi3JLWKBbIAJUHQezZdaYfVJy+LImh
GNs6FxqXtHw9cFZO9mwFwKs87IgZ8MCpv5j7QyRmsaj053z49qJAQqHuBvoPTC/3uF1QDtQ3PUhK
+o9cZ/C0WHiIkzc9yrr+J+ewO/zrkarOv65s4w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5568)
`protect data_block
JKyrdLS9piBuLn9uG0saFz5mB1vpbd4n4snlazpuT7ZHI4J45+Arld1E+A3dSXZHnRYASAcN1gG3
xX40XM02mYgjkRGucrjCdhp6k4TFm/05P15ER1aGHyF0TvN85umyGxH+OLBFpjiYduzkZri6kDjT
YjuQM6vFWgVJnhQgUHraffCg0M6dctRs8P4PyBv5wvND0GIQ0tTngSbd1ilc9c1lUbplIt5ymCBq
wOJ1HFTVHQuxlaembZnR2szq9MB2zIMVMPaTTaTS8AA2+OZc+BYmODoF3gEjRYcYBv6u0l/C2kBU
yrpy45mee36G0c8VMgOh0SjIA8nkptVBx9w2xNyTXOJAd9A70ZMb91YAogCHoHQLdv+KGqjW+sHe
uO2rc5dLF7sdzqk1I+v+QMPMgPIebX/fdn/PCFjTON0NNrLTxBsBqKwm52dpn5IMJFRcGWkt376P
IkB2OK5Srh6xwdjXycnzFUYS0zuFW04Qmxvz2O2uvLlC5s0W/DlOqGuTMYUVCmsaMrtuRllmAEEQ
5b9JBHVc0XKVj3uPvLb0WeRd9OUcoaBYx/iK/iZD0wewkKi5spCp6XarMXBf2uEejlmyTYzV9Z2J
DmlhKVCGFp3SrCYS2MPi8y8Cui2hCx7/Opwr5bV3KJWKE+GECnwuIIvJlUnYSsDLE/CkbQSNJcj0
PrOr9LM7SXj/aPHl7TIKMfTpyw460/Friv9ro09Zpjzp1mYm0cLwnvvL28U4UlNi+jVlLP/S38+y
itUwHtlLhui0lejseZ2w0WQwAumRWfezbthv+RoniUn1Qeux8TfMO5117NOfcHjJHC5JXAxBq074
IAGyWK9OpjKpg47fYe+st68Gn6YtHlcSR1zUkA144+unKF+isGamKGVT4bTC1//ObKIi3KWL/vvw
LIFvqENiM58mLfZKotgnzZQ5DxVQOkrhFYmAgiQUbOxmESFm8XF85vKVP3PjMR1mVovCQa3U29Fx
hOrotSnqMEsEHLhqHC+h0SfUW7Hr5fgcMiaDbPRBsVYIBS/ZuL7fDNuCCzuRXrW8xfIoX6e/yBOj
6lHaO3uKiOFF9BKNsbig8zBEuhUIILVZpvDwIUks6l8I6PEPFiIHIBfNWLtwjCgYZmqm5vS1Gacd
YS91tfLkRNtCBwnpqTQpt6b6tEBbcY+Q/4+DPHOEsrRqkSqPxWjtJmss6LDLuqgx1UgJkJVzECOy
LCyr04ABEoLhjH/Ia1VTTBMUNOv0JFRLxTOjo9/UIABjcAIoUBRkM4f0zc/Ica4+7uCB0s6K7JWu
qV7Jwrlr5G4NgfYOd9mLGPvQV+H3HI9A6vrvXxch/RJcvLGlgpZ+BcDEzLNETNV9dvdYr8Kbuf7S
AvGCJOQUsGJEUKsVsXTn3ksXodvNt71Zy2XU0ZgIw7EpoALmodYQFKM+I07Wh3lpDyBODaNAmm/j
gqFXdirhjoWXNpO4IGDMWHNbFrtnqURB24I4Qd8GvvlcEGyRNdLzV6QbKF/8LtSwPFieW32VTWXK
dYusRl6O3BjN9bh0oO+sdfgBzAEWD7VfN/Xji3ptcfoH7CJ7j4CtJSwFR+NMG5Tbuuxvn+4R+M4W
IcVIOzEmO2fVU6ZLsVTjRDh5ReNNQtmpFEWP8wkyE8b0fV1X+EbqJ/W4emMqlBbCZQcctardFF97
w/sN7lvafD9fl60lYQDEY9nTVxWqsR1zL9boUJ8Ah0FcNl271wt7UdQIrTn7PZ1M+3ifPnjbDhr/
h/af0qWXNAcZAmtBDId1MGE7efqSTzJf5ZdkkmFCADgGaUz6S+7pkf6ssdlUCCNkKsmVAqg+FsmF
lX2bO6KgFii652BR/u+vvCXFxuSLey0MIc0yf5TKM+U8yqnHiY3qGK4slvfMuLc/2M6thvZ8e9CL
kqHh4b0A6ukJ4Bdic4O5QpEEohyOWNdmTW40R1w7sJ08OAZzrXOUpW6hpGzC3AUVRC3DiCoEi1on
MBg6BgFwsp9pI3d6OWlLvf0rcvEIf8Vkur+Be+0eTpSFj55Ti8omUW14QIDzphUS27Z4i0Q4JdDX
OOHM4spke6oW48GB2cv8C1rZRsMgKQuJwJM3ZoERRJmSZAg6TdfxFfGAHqDJGCSkf9DdvxGEWlsY
CEnu3tzLj08kqufk11w+MZV6Q8wlTvQKmYQNzlXZlKHEVKDVW5KH3DUsE4k//ZBQDkYNKLIU/j20
QcDlU/Sjs+Ggo25lxnBvX/zz2jzND8a+M3hCFKJIu6nl9kyRZpjN/UkuuWavAhAeMKBUk/R/HBMi
ASvxRhbngkRE7Zs4MTODMStyTgwGg2tRGpLhqVL0FKFUNxCNO6OkligaIGFVug8PiU56DXZIQQtR
1ky1hCOiZdxPqjqOQo/GIpOq7YvtiyUwhKQMlJ7LUhj751FJ7omX5Amuv4N+ClrBbJtMDu03/+jE
Blax6lruolT/6o/vMeBG5lrNtptYghVmhoeagJr3CHQqvYw0NmriW9RETgWVs4m1XnlsI4Whp/Qu
0W1SECxqfZB0wdjztjPKXax7MGCSjRpF/vgiUm1ZV/GK2d/FZi8SxOZfrhZGJYGBuBuRg2AZodZv
3dTAqkJz5NkdPXBw1dRGp3Hk0rQrRg6iFAPA8nLmwEsH6XAX8RkxOmcBnO8cmB3I5DOC7XY/9D6D
EmTA6PbVqypklRW0E+EmyH5HDbtbSCvo3CePMw3gVCb/sa/M5DzzbxKtkmTDIAFKJs3LYmG9dxfL
F+nOtj4kEJQ0Tzh1ZjvtOEz0X5cyuw3Pn4OPVgCJZMB8Dc9FWw6Hh2M/4YKXoquyLp63DUPSC+5Z
H0qlkTStCd0tRecCcE9fQBD70kSQ5Ai/82Ahv3JYEddZNQMqyl4Cg5M0oG15XXE6l3YD2nHIpB5B
vg7ewOv9hXvAt/e9K6u6UmjW81K9FHig2sr45mHyiZJeIvpEUidL9wyO8NFcliL5mX48FWqJHxzQ
UuGkynnqHe1L7AXCKWOiSiUg760fCzLXZlH0ml8hwk/udhL8ouvGF/5He41Y3005H3MLQQ4XSqGU
PoafArz/sOdhxC6CReCOwjuOgy1aH2EezaZl5e4rurcKttOOgRKlCqoQ13bgUJ0nUwwO4kwsz3Iw
tdmPc0+JrdlPDZI1HN1ZFfw+B13vnFr8VMOxdBM+SO8sWbBREFjeWZDhppUYK0Y5JoqJ4pT7uHgk
5/1pbUpcZVvfuHE7eqVJ3O4ruNBiyRSZNPtFYaCPpxcR9ZgXbgWTKKNLcx8MX6ncCty+e7VYEdqa
v2DIk/Nv8228p8qDFVPy1QX+bpcA5pgZLDEJ3BEcT/q6aqcT+4wLINX/k6RLd8vHqJ/fjl0hew3f
eEHeBW+acJjfL6myTdNTdFAbZaobJq3805xDQd1ftkhRw78ShLUeJ2tcIdfqntEOLDBu2tmkZkt5
nJgXj3x5/RPCOf7O3KISkayF/rqeAcy8eFtS/GY/kseLUuIMXuwnTv4dAYwz2lAdahxbmpSM2WLZ
R7xrei0EhfymHw32YJoJstSnFCUP4VLJQOPChF08DJMqotdCYRfhcmbbqqn/EoJlbEaezaBrhw84
1V7eYi9WggzZecNUtMDK2lugh07ClsOgLuqz5MEHWFLXHvA7jlZaUIv2m8G0uDUHtF3M89omOoeR
dXk8g9pdO2Y5KppE+ffPhbdbVv/VKe7NoKcdA8qyiVlCxtFQM9ckiC7JERav1FX3yN3BgboJn06P
KC/tH3ZOgAPm3retJiaQDMfNo5Hx4yrb+kUHHp5M3jjBJfHA7u0blu8ZHnRO8RoXYbMga4Ra7cW5
tQzzehJlDjDA775Fbg4/oL3NhMXSlrAV2rIjCeTAiHjwypn3KoxlqqTDGxTIWVXtDOj4lAzDZQpl
YztqcDaHDW7oEQOQ+s/Jds89yKChoyO5avgGIMHqK3vnU8t9S1S0+p0oiiLUhXDydHfMNi6VoAe9
WsSIOXcToepRNFkyScvFqBUxAT6LEZV6D+mz26SowK2rH2V+1so1n/rRdZYWZRNqnuiBvhrFqgqY
TQVUwcCEbpnfm7WIssYrJwyxP9kWIiAwkkSFAdSjuU/vzKdtB+p53txWdjNL22vxJ7cChHUiBgNG
4SBiGLi4Fyk3607221AMSTjm2A/sOpLFzK/XZzfFodbvrjPFelAPYyAsWtdg7WrLFciQLxFV/HP9
g1Wuw9LXdlZ4MR03HSDk3IzUdpKX/LSPERpvLWLopDmSI5i4xLMEnEmTIuXoPcah+4/rycMD4UEB
/88SRp+ajmCWW5Xklxw8E4VgLdKcb+TAOunaFFsoM21flxGNiCikjyhJIBqmsA4q6U0BmyaK9pi9
2iZymkkP4gBQ5ARlTW7KDSehpf27pLyfefIuNFOIpgjxDZ7f8unsxPrvRVJ9lF/dCjjCfTiCkZ8V
nw2P31KzvV7/S1bA47BVLOahRqnD88feds/FVgaufC5tgdwj+uYuq3WbAX1SRYv/vy38rSts2UZT
AK6PXnWyLpBPM3L+Qk3DAMby7yvAMSvgeKfqwiUhpvSLnjX/SGsxk0waAwcIcaOtTSruYoYKWV6y
A4urxGXu8/+G10wTGq8Fa8Q4sQ+9CjnmqCIWYvLH8I9rDibGbJp9+h2XSrGpIWJC3lzVIrYXLufB
j5crq1OcheSLeoqvj09ZGboBuxFCQN249/Nd28OgufqbMdFz/jiPadMVwsm5FnpEuT9gEiADmj9u
pDJpIT2GLhqScn9D9zcEay7USEWgUxuPLPEq/PzU7GAF6uCENnraPG2gJNUi/V5wPEZpHE1arWJ5
RIbZt9quLqzqHlqg5GIZOA5IwyZBYj4bZzrkswl18bpfB+BPRU9V9dgsMTDmJolBxvB3Jnwu0TIb
OtIvDgyZUc6BBxSPK8rRJ+91EIVl3L9sCy/Waq6MrI1LjmVN2psiXIw1I3ciY5Conx8wd+YiF7AX
uxDb/uQijij4X/iz6n641s6pr+y8sGnG/f/vlKmTzy9CW7ypGTuHFvG8IX3wRMIqkDV3kblMVP0w
pIrpFWcABnAIyQQfFO+ueWaRHEOcZj1cdq3BmZyr4o19og0QRqKxY2z1+Jl8v+kPfEQDd8Sbz6Au
fISwOVCF0Kfx8POVkCeYysUSYPsp9R22AJIIeKSTgZzOoN8rN4Sd5ONdpgJgEb96V2HyDUVWmeEv
8iRQbd2X7/dTmbjQzPraR1ms3A9cUZ45i49QGuBe/Kc13eohnKPtx70cYQp3pO+pBbd6ElTB21rP
B7i1ruWsHwSITbp7KCDK9t+EHL+v2muX9yRJZX0q/Fjaz0ApXXliTy3o9dd+seCH3edEImK6Ofl3
sANpPIX1hKTP7CeXa9mGzyX6RnFAQUa2sraExuwGityhx3Dqb824P7iNm2JosPi/DORByYZv8x9e
LG1NkdC9bjvSCgLT2mRf5PBvjTbxqR0PNPcOhvnDDBaEP6osE2HRoZoBeKFxy4vGibjqp/vgZdo5
1nLkDfCV9NMyzHozQDXhOcwtHaftLhyJ+4CAOV9B0Zr/awFxxUhs3xucS1EBuIFJxesYbxivmkqu
BsCKcF1MwwGkpJN9MpMAdLfGvR/gQOTFo4tmFAokFw6GVbnTtpcDL8GyYmlHecPQ9zXHWP9AzED1
CsPeb6Tzj+Ld1W3G0pq9WL09YGFTrBTjB8qrhRlEqQJ7HdL4JWVTNZYHmecZ7WCpJNXlsZtNOMzj
ufgx4wCJiy5GbBYGk6AoiL5NxibOx2C4qx2OHbbaEyCWpKfSv3NfKfbW4lepOn0AI3gvWUbAhBt2
GLzurIE14mwbgQ9ttsOlJHZJ2UJK/RnhIzTN44VnJ2ZbGHhvAQ131NI3Y/S+H9g90b629Z8lyRmC
iT94AJq6lIQFEjUcHlm7QZ3mK8RnSO2S2xCF2XrA+XiEpz7alwIZ1Cg6jjwY9M7ExFbTeFbMO+U6
5nFjRqS4IorFp8rQCySGDp2lUq4HkGo6z6EqMH62Npk45oAw7LvKqWiu9w4nYhctVHyWLD7xIqD1
uppt6VE3vNPcTWEaj8PtaB2Ze9x2D29Oif31X/yq3w6N6l5UokX8MNbmyhQLwp4LVXT0QoBR4dvS
iNtgUZZUNvgJI1KqJiC/QLeDaDc9o43lDg6AL40Gpjsuz85zWKkBOX4sCmZL1j4jCzpsAdCkK+15
QlJgOeWawsU05whxNF4V0TXYqDP2W2y8jmhhUY5g+tvJoTb9LBGxM6GLukNRj/hBgh9XaKV02/pQ
hyRJN1hdQKHQDAItoCG4cWQShvx22bf4+PMj45WxZO6ON4+2mfjIxmkD4bbrmV2oUZSuUwjl0+JZ
TrBRhbn+iRCzNPf2+BzithWELowYa0kVqaTiQQFqVlfGRdNGX7KqSLuNHEiBJwcWZ/INBOp8guhT
gl8SLC80KaeRnqkdM/fDOCpC2ByFqKO/xqKUYDGli1jdU3HB9IW/OCJuyaLwJqWskf2aOe6EFje8
dh+mZJYvYdGaAak6vvTQBcVBiirZyMxNluIrVsx6EqiqOB7bNpYMKcJ6Cd+tVboL+edQybBfH5LQ
Yd9wBIp3rhc7PYl503GlkWSItk3oEOHoRbCWTHZGTf5JDRhc383+9yYZAWhhgYwQHR4V44ZQEUw7
7PQAseZZGZ8cFpdxYapC7Nmtn4wv4PTCBqtCgvx9aoxAxPq0DaZH38np3+lILflcDAwuu8o3gOt3
B0R3d/+X1nr3OGdygZXdU3rMRCdKrgmnJGamkRaSWV7Heahd5d62nOK8jjbDZCwtijQWQ+74SYb0
PRQvVZIGKUZq6QWa9JFo4SQrjflWkul1XY1baJkDBG1S9Dbw9+uCyFNekaV/+31Yt9cbYSJTNkd1
dvfxrItY0Vy62x6kcDUMXG4k0I5nF7MoYs+S/BnNEID72/q5lIBuFvVIqpAwNIMMeu/9UU2m2Ifw
NZJUSqqnU9i3Yx43I6R24j6LbVlR1q5CuCBvIeMuchHp10OhoaMh7a1L2bed4+3++SwRQ0KSUckW
Z3oMy6F/mbudvWdKRmM1dbRbbQ41O9HlrrAFr9xh+7+XxsogMVxd7L6CzBCeZvkWftu7iWFcfc09
+MMUPLqohM1ur6APBaHvaCvFbKjSH8xYG41ckP4FeUqvIWqmcK+ypDbl5QtNsMiMyDYg5NI16om9
JPFx8dKHCDhhMZ+YuPn8kWPo0NzRe5GMw7s7T+Q7gOnT/IZ2omR8psmf45vxCADKY6bmlUlAinR7
YmhG57bYzG0VbIc/0sf5erZc9QsluvBYV7kdyqQDenDYb6Qts2RqMk2Y9F2271rfz1UkZOcns51S
7lUODsqPAhhKCRo9PIvq7QMUacsCiZnQ5UMHtiUnODGWzXsdPlEr6oyqIiEoW4ZxmH1Ub6BzXO8K
jPzm7ekb35c0E/i0p/Bwxyos8r+lWK8aMn3rcuRqkFdgIQmdUfan
`protect end_protected
