`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KhvGZYsJq7NAqX7KQ32kcNhns9A/br7U1R6r37FT0lYUmHMQ7jmQ/+1x5jyp7BmuV1j88Vg9MjF9
1zN9hBjNow==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TBaW1iPJlfcW7rBizyMdUjSetPBdGPtrIRz+AVpGlSIBbdSNaWFCegcfv3EicMi0yWksULMs03M4
V+WSvJws2yjpLhEPf8Bch32X4/uFAblVwb1SPRw/0bV/AfLOfKDor7lQJbzxt4If4Hawpnf4p9k8
/ygE1grCSTQtfFglchY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lXCDwn2QHWBQqtBBKrevARZ0uoVMS3hNH9i9eaJmV9KA6qMv9mYYha5axdvBpfno6nKJ0+LNATfv
lFxMq/YWAtikVUG+W8ErxYn7Rd9mW24DZ4BJyumr0TfffjhnO9o8tvecsLZEsT1oeq4leqPBFSg8
+IOp9HXbf/uqClI18ShdPXBcQOW9CNphSYe1JMwqXFzWyK5+YvK8Kt7md08dvqBzjJWiQc+UpB0I
7jNMc2oteUbA4Yo/FSdc0YRyivN2lkvHiKBjql/XdfDmeDEES4L41s4PAuzQiJqBoLHjLJzOXbnA
bCaxuWJ6HdsqUhnt4X7WCydbyPF7jNG5gppVvQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dIe0PcVRnKlzA7UBdHnjOPz/wWx77WVJtLu1HuM4yEmdRwGOJdI679SAm4Z10m+h07/fZ4xFHviU
LcOPE0o06RGftFrpLcev230WkVKvCLbK744kEZIM8NlflwuCIvHn1yLmtnx4RbtcVhKIFbTilyw2
iZNva56wzI4H1J4dDQc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U6uxhxmCg/7wnHZoUW/k+EfaFIhouQPdusKGexVoiYtyrn3q5341KHF+VEvSerGnrOwW7igkETL3
p4zScVaP3jxXKwckGGDlMWklg7O8S6NS+FAJ2ZN2mFxKoaK6rEYdQiJRtYTTt/DY9QXSpZ9J63sS
EJ+RbOdDk7BQC83UU9gK2DGXDOnaV2r043Od3O4H3o/XO0f0WookNV1Rz9zDZZz8NDueMQA0gm4y
cZV6dsFY1oZ7M7JPjEkELNSrZnPDuqaua5wALn7E3JqX9KlYKNzafhBBDwRf83AIVSrYNj8T9Khn
V7d+6DOUQjfrWYtAZuYB4Vodrt3EtRO2bnghOQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23344)
`protect data_block
eDnX8OJaXW+GOUCyk0NZ6c2obbsZq3blmPHqdvFEcmOFtIir4N9ZWA+1tJ1MYsMrdDI0hzyp1ks4
Em8AuLS+XSEP68fevKs/TZExHQh0r3qrHG+Z6Yy6r1m3anC+yFk/huNZdMsptHwbyvk2rXdfcdCr
fri0ZJdtcjgpp6w5kudWqsfqqweQZyjZf7akYTcOzG5NcnavAv7QqqzTcEjd4QhOws+B1jLcPbBb
yDd58tfV+ScoKHjOEVrZtBT7FhML3qcib21oe9CT22Q/OPGnl9wxweQeSBU9igvgs+OdD6h71Oue
vHF2GOejdou1D0hEAULvIa/mtWi0xqCKWinYt9r82UZrYqeS0SN0ppjAjWF49xJ6myMxz630liag
gYSdAQviE89OV+N8DG37I1weghBfn5WoDxCHDY8B7k59+mUIUQDvNHTsl3k7zNgT8imY8F4+LQPm
AL2hK2c8EzWhP2Bskc9zcfYCuaGmy3ald3hU4KrPeMz7RN70Gycixah979/RojmwvdPHvCt5zw03
3F1QjlebUjNfhEE+yKOVvRkAauLbCv8BwF3M9Zxlf5COPIjMSNtHQQiVXmq4qAFt24gzGCjVP5jf
W+x/KprE/xwTpBXOOrJ5gigNWvC6SlfY1zHGOlxQrpgyE4v1AXEszWkPK761c+azQtSzZPAWEiWx
v5ctJIV+9yh+j+BzmOztBpD5Nhz+koASPO2UyQVcvhq4tXF3aemZqK5NgeA/GkGn9Zk/cLZqjrck
7Q7mPorurPzZW3zObgcchzE4bSGA/SpD1tAZ2L9MejLgjRZsAvin2lZBplFd9aAyCnQlsI27i+jR
YXWdNr1DHpKLIuwdZmD5tQ1TBFoQ1+Zgn2FDLFah4V85ZCuao0VY1e8PCjHyTdCzC3Z55uuCN9K6
wKqR9t+7HbM2pL2OvXDASd+sSinU44cCFQ89dryucwRkA+Zm6fFaVmXTQAcEc2bBrLDLH1tppAxx
I3T/nqab2nRG+ina58YzFkxavcqgEwMUopvIj/4j0p8frHavl4/k9z9/cYOpog91lgGpEVkDMn2S
CY09NtGaGks59bDLgxYCjzzYmfBRlEFgx8PLayQrHDxBzwtlwYBrQiNJogd4OQn1uZM6ptpnBXmm
ygkiIcN0mxgodNekYCBxr28Zm26ybNdCWgL4JS1qxGQljjsCsb07lRneIsMZ54fOntTgjw2ZJ3Vc
HJ0OpYDOiqo8PfuRZ4qqKjC/J0AI5mYmh4bGBE56P6iWhJiA3mciJXBR2vK2+BgtCgD/NGVhVn1n
1eQfJQ/hB7Da97BPob+J1yAlNK9J1kaMeZww58jj1SbqsYb7PdJr8tXWAkPY4Yiriwt3DXtsxCwT
UHpUi0R0wPbRTm5tw8bnCIBrCy8BHHjO7CZ6CLFBMlWQAUNfeENsYMMtbJQGF0a3Rm/xIESopio+
7sKhMFaF6/9wFl41wdkWQ0AOgI4HYN+lUduveh8zzLDbN+eD5bzNw5Harbof34A5Yr5RtXaI1Eyc
+nMcKjp/0NUuCptnAwHX1VPYMG6di0gm1yr3ujMWpThDMNyp/ghYxwrnVE7uo/MRAqmqj/YnhC/E
5nCLimDt4DVVX5OmMW/gLb72yUCbodyiGEnSAaVXWd3f+MEgieb61jX/mXIm/0OZfMNy9bDbeV6j
V5YNVmtyjOJU/gZVJG7o9/w8Q019OAp7dwKqkJYp2zHfumoDo4/FkwH016r9rMSaE9v11ngmAoN4
YW8YKJFJaG0y80ob7A4OuVq/SoIqdKnGzr9qUYKOoKDRrimAY0eQjIU1mUQxZJdrPkBzRF06ibkl
+4gyL0a4xBswMNOs1obLoa66m5gIfrBG9Z/xchW7s1CBii8U3iLsWYBC7rWcELN4hDNBL5k90wvc
R0qmu6VJzOyEwjUHOi3ogYD9vGQXxe7MPi/znPtbB0QDXY2K98qxVQzeAXCDxDjSinrdRBIlQ5E7
EMdNZuFB5+1y/JxHQ0irWdJ0u9yKd7RYJbNchGb3Oqh8FSIRH4TcjLJebe7AdDePgMwlQr0sQdY4
ijuIU1e70k7MtAUpa0QmbBAHkU1wCrL7DY7WT9Wsb6LL9i4Gs5OIT3hNrltckkmoPCuQQ8tpGCad
cxXq7zqbN7Fik5aaC5hn8MoUBVTpGtazJcBMs7G4vVM0m5HZgmd7wSq+6JQN0zOUs1NMHA1Fpju9
ZGLftIfGUuAy6puRsyz1o9SFaAczyP7HDVV4bscm6dPeZbO2KFGIRfIYH4uRuD+h7LzoDLrRJTmr
dDu/+Ys0ElHPnPSplEIBn/P3ltxhR4l/bQVbZlRP5dr8FsrDiJe3LZyCDKbIztMBR+4qGIagSgJt
W9tFKEB4/096Oso2WX2zMBgDAR+OutrCAp6kB4Cog4MHVvfla+7fKl8lE1FBl+4qomjEtO2HCSt5
JN+3Jtk5FgeA0QHLNtYysP92pfjr2sGLlqXvNkPnpo9X/JduHQUHw7k5ihXGUKIzuJFYR+rzZzNW
O+lkm+7864QXYERN+lQBbngMmJDo+VnlHtrGJ3T+40s29Hulre+qn+/S08WCbLFhKjQXZ8YW5WZs
fzYIbHsZsGpqjDCcGxKCYuwTLTIIDridwz79q6ottVtcZhDJPuKuISUsqg2SxFdNBhInuXa3AK9i
a9f+iCyzJNPX6A9IdBEKRxYhhX6uOND9ktocij7pC8pJZ1iJvYf7nKBUBIsp8sg2UddQkiHz9xur
WLwcXQ6NUm+1GOYwg3e/0iCpWKyjZl34hpCRd8o9yxFxkCW1tZKlj5qFocHxxQ0iOiOm/kQnekRD
7IuvQJPKjh53Y+bobYVU2XDBtgw9eq1GmBfvuagHIK7T1cTl3RvH/OKV33+guCsyhwQt4Q7vct00
ftq/ApL6qCcNvdfbDOGKpuTy/FIFZW/08fZPWRuAFHaQldIpI/N+GWvwbbsKqo4WhegoC5STvzBH
oOzfdv3xQfhv4Q2QOwEcWaNiTJdXc7hF2Juja2zDhDzS0JMZtGU1bL+3j72Qi3AJqmp3B3Zam9G7
EhLg4LWoelWYJQB+7PgTfzdWdi9wYa8T/LOiHoab/8Za0+/lghKsvOI+dwlyp1uWENgXqD4lDf3c
2JpRytXhH9F8yY/iTmgAgfR9mzhxptdZVMgOnA5uyn8I2JQoIIsVnCzCro9e2SrskLZ37zZC1KEE
fE01ZwTnOKr6TdTVaThSxaGhBFKU78LiPJNy0+49GpoAYqT7keXlLWN0HkZ/5y8+2jh/gK/0E+kI
5tx65kQRKXFsuUsmJtf2m9YKsYZXotFb2OhfCQiahJwXB9sT0KTQdR1/X09jcv/FTVoedcMmtU9f
LXcQWq/+AyaRVeAOc9TqvRrB3X85EKPsfQVUa+29OWXTGDiIf/tg3XZ2lcYnxjHoygxovCTPgY5d
lScykfTdgiZnsoHIkvMTZ9bi90PmwqmP7PdYl48a/fecIuLlxBt/sK6oxBfBiQCRfFMTYZXBfpgS
vDVU2pFm67wLmUflUQmeRrxzcNHi5yjspajms9gyn1iwRq2Ow1IxSX+wbeRruc5aug4PSDDzj7WF
JzUPzvxOmZ37FC1o6JmqLu8AlT3wdfhWdjAZfAp8CuzRJMYD/Ti2o4waLUkqv3uLjzV+0+Jcgpl+
s72J8qjz8HQOSbHCncZayhRfuAL1QJRn/PzBidhav4XFcgkkK5fBpmUvToFlQ/R2gcRBrba4GJbz
VgEuxf5eAk/Mm73z1AZt8ZLLNb/R4FG+n7QRjH6wVi9Rk0ZJrEQ76zHLy39NQ+BjRAToTunOn5fY
9tfEkqGJVgsSFe4oC/QPIOUXx3oSj3eZ7VqZOUouPUZVEL9+viDHNhh4+GAErNPJyz0HTtOuM1gG
VN6PfjzD6BqGNuvjF5h2eRGS2BMj3KRNEGQHSNiWeq9PcZLuGaZLesE4q/28Zdpd80gMnzU4eQEy
ewan3BVmMmt/s7Lh87+/5GqPkiVt9lU/11k0MS2pDXIjg+nXkbKSV5qFZfHAIxUp88MpW7Ms+0xw
+LmfyMVn6tEfkGvhUIUTRDtHF4ydxd8s7LMvMEaDP4WNseMOUsb8tC5si27aVwDEl9jg9257bANT
cEblYavXYd3yJ31/XASikgRpC25R9p/hKMD8OKTTcPAR90KQ17yha1MVKeVQKb7TqAbchQOmuG5Y
4gBWmNhTFbA/0RyHp1+Ac3uamUZKaFuaeE9Up0HyDEyaSAF+0YMQbbpdpARu6OIDVATiJI9np4L4
mY/gitiRb4fJoOskE7qGrTSeoF1QCO/0NeCoMoAravc+QyzQhMF+4oVzOc+h6jrCLoWacwKzKHLU
WIemr9KkUmrGJah0VNNgpFr5R1wA/8Jny7pXZM82Otpc0S5FWVfqO4z5KSvqTRq70SnGhFvYUiEP
UklUTaxkPa9J/UkYRWqxJ+e0SGP9OIgbl+cSdqV1sVhSQz9rITO/E4EL6mOTBWlu6QYY341d3BQj
KX9EIWXYAdD27d6hiwyCgJ26ITYfYC9RNjrHE/qIc5rZAfhCavrR9gnNUXfdLvY0z3P3TZqjnniS
GOU3Updvq3Mqz+pxWoTJfDK733rTzqM34z66yHxVPvM0EZ9jbDIyOK6iN91ee7T3QqaryZ4cSqUF
NV55zuwGwzhNiBaKA4eB0Iv62z6JysSujxr5Up0lMDprFPRSYqnduej7upfZAJElIcBiIkJa+smf
m9H2zbKaeVTWSIuINCEmv8gM6q7IEyM2Io1Rg+auUdVMR/V5aR6CZRx0E7TAuLea7twjZXys+5mt
1snrL/OTG4azvsSmIY/ONeGtIZ4sQAlZOe+/cfRn+0ZENMhX5YHbOarozsWZ1cXYUQAK+ErK9BxU
Nvn/yHWWncQ4galP/FZuAnoeJ0DsLeNJxa9stLIcdf//JGs83j56z6kmaPaadDhJlciDY8vhzlAq
wFCRoDcvi/2xR/pyNpNTwX4alXAddCxpupi4KNV94QtAkQQXuUG33Dv8FAyzL7f5jd7GIJ2yC3SQ
xqMpVfW8vENYW9elDk+OM0fwsFExwT+0OO9132ujhszcltvtCBqUlDLiryyiB6vju0lYqhlT2hnW
m8H+akuu8FitGAmCEy1ppEyouONoc/y9nyTB6Nq5d/XKeQWKhxhxMRMJxHK9ggcjw+1PY6pdIXkX
XKZ3b9gqpLnYcpB1N3dPLyclp+Sgw7PsecRMQ1aDW+yY8NJ1559hD3jMfRM7q2mz1sS2o3G7Ba/M
a6MISWOfN8mapvFMjZDYM6JQ9eItCk74FzdNTH11bN0YEMWOryO+QcJUO2vmXUq0WpHJ2wtjRkHI
sZXkml1s8zZ8xykytsxkLGP3vB+ia0PYDBQ+fcXYUgIEVIJc/wb1G+azlBFE3os+R0Alnek1OTjc
BPFY05P4sRPF0F43Y8tB93mBsyIQGisH60q7s1lmM0iV6n4CdcephhS3e6HdkUZypajXu9Te2pmn
NedVmwpGDmjOyeqeETBLzvaQRTFWzRRuoLH8FwDWccupjXaDtz0go3CGNMmwO1wD57TjaPZ8rnsj
XWGx1Z4D02RT1CB4Hn/h6bjbv1pAnluAL8+lQUpLMh2+DLBakiPgCt8x3D0T7B7YecntQ2Vl8vrU
DSjS0eFIIffOGJh/jXLzTKPOU++gPeztdTS+YgI4BQZrUEWPoWVufrKQQcqqt2TvJViDnV9Tli4s
jnWtSntxA4/FsYZVKt4/B6UCoZ9r9icUrKSGsWU5vXajc63ZcHvZKhEuH+eweclA3zIA1u8PVwGr
WGYKScZfF81a0pCtCkId4lTxHWx8zOi9UeXIaZYJfEsyNAAs78otkCwRMYPooiyKpxTTLaflSm4H
mWyGPvTlJYUQS5QqKe3bqRApj1b6YoVRzxXthAz23hmgOwLVHKwPF5+Akd4o++sw0IihMPIf9FBE
843EpFc2FRw8DlXIGFolcY1NeyN00PDngut8XAjJtbm3OWDkUuTCQNV/tVt3LWFQsps2EtQ3qP4s
uMvR743vq4YmAE2Meu4dHcRRXbOo4oRTst5wHHe+AlIia/XZrYiEABQ+iYV3UUjtq6qrCIcT1Nlf
Q1T5QFdOuVh9JoTcdFlklbiqjlRdRw9mj31wycvtF+N812l7TW7p3Dcck+rnKFsJfhXvNJX/uV1L
fO5GJbQi0CnFMWWX36g+utg/YuSSOwgI4pJiNSGxoEpzPn1X+h6nFG6llW/zRqRw3duOiPlG3Ous
sDUVsLWxNkjse3q5SbmqutgANn6Yj+p8ZP1R1RcuxqBxH9Sk6o7j0tyf/k5KopdAdeD4LF1Ad9sH
bx7KgqlXI/XgPuqXQT/ypDt2509BOTuUPRc44sGdiClQWCH7FpuCr6k5r1vRlHZDXLUnV5JDGZTE
3FB8Z1PpfVd7GGQrimKTMYxKdhQlx3vaZz4b2f8vty135aAIn1M1CffUAhWFduOsnwnO0+lWWuwr
/hMJR95d3BI+8Lm0AIT97+yrXNok4U24d/oeKOgdfDaND96Aa99RfrVhdfl1Otl9Obls+/uhwQCm
c5h6AF+7YuA9etAKADVBu9sBzuaTNwSlf2JpfjolqE9jOTDIZkNVzbibw/7x0hxP+mClrF9z8xhJ
WfH581h02yoLATN/goEbDHIKsDVCz1nLVwp1ogXaLIz+AAsYJ58rtTKjo87NBArbqWlU/YYFh1Wp
nYJFpGagW2IyrnAi3dtz9Rv3kh+K6JcOnjJPZM9GKVAuCj1L0iNe1z1SNCVGmVmN6QkKTEHjaxBi
fadWYS+/11O1VTHoj7a/AU8eDJmmih8/lVcWLIK0tdIPU72MUBvA/NsM9uHQZ8/KQLGq5gBOinSZ
JqqJH7+7t3ty+bUG3D7jpVFNM/GOJTw1OihfDq7Rflcp6SfG+w1vrp6PfMP8jnaxbMtpDZmskE8l
RW76+6r46pioU0uy7jAO/myXy5PGUXgPXplncJ5DA63crXc0ho+7JEHOc/OmMFm7Z4T83digpZXu
Y7gMepSHLakVp8EBunWdZP9Mwnm+7rtTj5VMYp/TQWemjZKjS5fCKUX58XDuZv7MhbGIJQrqXcO8
wDd6kOwT8H8UHKI4b6E//a6cdRBgxeoAUCNtZnLVgtU9MbjHTsU01hw83m4MSgBNV/bpS6MF5+lU
+cpwt4nuKQV8evBNq2HSop8f9jCwhTgbZTyDbMhJJNsonr+8mFRccGdyi16pMfGc8iQaPXu8//2t
fC/IQDMALyqIyKiU4mCE1lNOmkvcs8IDPTS2j/6l4oESmzOBTtHmqCuBRY2YpGViiPV8kAznOYOO
6A2nWhGZeAWE4l6lPo+GtoVmPT+BMxlwuEYP1b7ubvQNnKnznECdOYZ3bzQl3c7bfEPsShgh/sif
88uXD3xE/MjIUWW3kK5SfrpuJa2vHgSKJfvwRTBBCESts1gpIPgWxchXT/ZdHjF5YZNweNRGG1HN
IcEV5pmhy+8QXuAhRpGgIPC+haEm+GW34SBe6tpLKHm8E5eG7wZ0eClOfP/V0oAgtqwpYxI11ftY
7+hb8xB6QsobyU//4uDiBZa6mQRouYGEfqWWKhfyGB46kJUbb5AXpuXTW5s26olHg2rJMXq7/HuK
IaqYTxw/PcZhcd8E+rBKSyDm0mUs2OJE6H/2yYkIhlfFrWm9suoHg5Cd3TQrDWh2cLKW5PMJzxmV
tlFvistSxuBrAVAac9P3ZuyuwYDqDks2gh4w9pjJ9OoroenG3qyBkDonsq1OpEP53DDeS7bgnzb+
369q3xQwhBm7bhK8OqMidJ0zcb0wcdq5hqOUdhSN7fUtb3LxHHbt3Up7i7g3HuKFNETRmmDyZikd
0NYT7Ri9qsgmtFQgiUvU2KbGr7+c6aMa39eMcel38AwS2/6k0SHy5zXBH/3Hw1htItbTOHscTNBq
ZW93Hfbtg4S01j0efvFnR311m8y/8qJr+TMiLykUJ2lQzdh68RQwJEYGh6SNjugQ9AjWVJW3WuMz
F15x1ldeVuQ8NJ05wZhJsXtUIK5YiZx9AmEs4HAyZCCKtBxVnQL6craIb49zaB/oHDn2aPAVj8Df
feTI5OzioSqA1jjidzYBcJqeokEGbtr2J1xQOcB9LgFayUjlBg3MObLQ6UMvG4g+2HxNJ08C4n6c
tgk+KQcoDd2u4bmeywLCSy5CEchOfaT5CiEZndiJH/Cy2YWNRoiD4FygA/i8M06soZkD96BrmGip
HV2Uqmi4yFxakiaYa1zLCLVA14V9OdK1KSkTSPJns+JTeLhGEXa09d+jzgvFgNDy+6+aDxz21Ut8
OYN8EvWoG5e8oRUn5CXruy3/TlhjPtdastD/NzAISCKq97DgXpO+uNfHg35hVY4vZFHIVwuzXFHs
JUgE9jrCDIKkz3MikpLXycBuaruSrOzsy/JFCnl3t2xAbWiSJfMb0YHNr7fg3TzJPRoGcCE2tavb
M2dwYrsKYpGyflYmQ3Pi4EsMNo57Y30vgNHXG9TD+ilAJSKNutAwSUYsGxch2kiDnP68TJvQUWIJ
eRKkjVzKEiIZ4bMB0V06EixIEv0xglg+qt3oxkehfzNC6e3pFaCAy0lc3kaw3+kivOhnF2/ziU6r
8+GmO22ZqgOAWWwPyVxaI8oHnsRTAEyPTbueFSvi3bthM6DCW3lRvtENmgHEntrSdehXoIjukpAW
5kz/DVJlHqRS4Alk0GoB3MtQj53Jvo3nL00mvCRZ8uicyAgmFydprCGGIjyGOLaD3nx0cFgvnKnl
+W3+4SChe92O1/P9mpDyY3QP5hDWliAhmKqSyeLLiE7eS5QBUviWZj97l8rcTbZxU/AUPcT4mEh1
pTZO4HTyjWiIN8jUZdMbn4qJA1j9CMg2FtVBGwnBNo7yzZgw5KDZrughbMbqhOusLq5ojc+qNbpE
KnJJfV4ktXMvg+sA66oNA2NrG0zfeUJMCHquFRa9yKLqRfyK1OrjbOn+pYwodhH3IoS3nzlzQ3pB
+3MA3KejaGmsT1oZ2dP9BdYylFO0lea9+UF1E8zBTttvmXAD2+z4dq2fPidko31Amk94l1cYO19c
qs4j63qy/URRq4Dv6kHqI4pT70roZDyA5HMV9Axu22tGz/4GkwELlCrSErynIzvgoDzX2dHENAvA
h2mthGZE1OSmFlrOYoGItW9qOh+v2zcqOLpgNe/kArU/F4H27uKVFhf+s3yC2Bs9zhMvr23y06LD
PUI2r/B534+ClkXd2omZNGWGlU+RKBDkQShMIDY/wyZ9rKM16QHPnRAHpvo3Vl3txzpoU0CUtbaq
hQKb/vEVGu0dTAsYIcbAK7jP3VO8H9+0Qb1DexpNuEb0pZlUE4gGkwOUuPu+zVNPLBJi6Ha7yhqt
lhiIDSQPzfmlU90qbIqNK0HtvAPZSCerN5ol+Q6zMM69W1j887UfhQP4r0zezcMmNm1BWeADkHMV
3vCmrOxmF1+XgenZiRinCw2Ef1i5DX7lFuqdpwPIYGT6S/3Y/nc6EIwT4Oh/PN852x8JLdD5LA55
473FsrDWtUcP9Zih5UCZRBhWCmhsqOLe0I2Fu/0AulDK1+KuWnyYKsIGorAxlYPFUjOdcrS/G7js
nU0/Q57vrKU9bgcPFHIUpWuNdgPj4H8q/e0emSGgSf0WWlAa7D04N9NyYbpE82OIA9cAiddRcvr0
/5bueyUOxW+u/tjKjRE0mwyh4BbMOTMIl6Khj/o6STEpCh37ekM7lAHWldCrn8Uw0ku65Gp8o8FT
q2FQM6UYjomIZVnDtelRWYnpn5gMrtVQAuv4Rq6WpJmEDxWUkjtgmjprjNrnvHf4hu1N2feej6rC
8orKKS24ygj2MJnjwzTOGcDQ85btbyRNKNFUpKoNug4S9T7007c2nmMxqKzzUhfOsp7pJu0t2YYN
movIUafnFaE0tB2IVzAJAKEx88/oFrKRsYzlIQkvESvZOj06qdGoh5UkM21ls4vXvXHdcfH0FUV1
7FYQrf07KF/dE/G/L4783r7wUBdDd2RNadVulku09EK8ZLFgxHsTqFLIbfovR8BsqXGzzVPc/HKu
GF8Q9inw2QlN+1xcM/7R8Yw5XubV+ndbggEPNS2nXsuoHJk/2d46sJIVwgszp53Ezin8eep6tYLP
b23NIdKuGxpogueb7UJROG7WISP4zPipRcpVjeOsJgoNWB1PIgPCOoZAMVLPdTX+w4NbqGWJk+5y
+Jjc6NsU88w9kO/xHl2jy0hh58L7+YeXvPLg1VxvqfucvYXqPRANK5zQftazdLXsW8lI1tFsKHqI
yjrz8q3yApdXQIrn/dGYOqiN1qU3Lw/icnLdDdE7sLcgmE7H9Iyg4zKIbIzciwbkutVAGNn4uxUU
HHfSaX0Y+aY+zs/zy1Ku1haZFmJj+q14d77uEeJYAaBXjvsKvRSCQM60LJakOxSYMVLwyu56m6QP
w0/V0NloP1ujF55LKdnhI3O7QmFpf+HlXrdZn4f5zH1WDNYjhgnA+jdGsOdBHrY8UPUco7o1SZPa
iD9XaVDcYco/xze/MOYeIjmpLNrk/w49c/wWWzvrPTFzAbtpku9WiTcZ3rqOiyyOKeAKfCA6aa8z
CF2cyG4h79LTrgcYDrmbTE66D704EcBZxRxM7FNcISIPlZbHyRV876Uk4wlhkuSgC7at9yuy9KkI
piwSOvghXOFcgevD6VeN47Nt6RdfMeasI85BSJuRKVEVv/RbIc7C3pLF829AtQvqQBo5p+5k1R5g
QvMXh9jm9TRSXmFdQj6caWA6R2YtiWP9+dXyEEuGQZvNWTv8A6XG03xCer4BwvUeQvH4B95uWhw0
KOmXEN55uP3Smgl8GZrW0QfRaSdfN/bscwdGZ7VB5h2m0HFInS5Zh+IS/kZsF5FK9gPJz9MFySHL
eopI5+vUsrmk4mukyMqSjv7r8kVIDzsl/eVhCbUBLa3MJjqEbAUlJ7oiUg0WyMp+iTVJ7/Zn2XwT
2rWJ4AYUNUjiHEvXLAxgpyFqTaCZjD09pR5rFvHtcIkiSPQClESmUM5CBqlCR0YmVxUOqZlOYekb
X+UEpkW4QtKhx1fIjK8hLVwYjNdktd3gWgGXyiR08jUigO4H0BX6zPEBiXIHqS9hR8lH9aCtA7ht
RM6rvjsDD7IqFBDgyqAwM2rcQLe3zP3kBwqxskywO9LD7ruKXx5Q5NR2M02XsfZEOot73TU2V6ja
5M1FEakKcm1a+B66J5pdAGps9dkyLK318VcFJLS/XSTYWBGkXivtJFaHOIJPwk5iItX9zCCh4zyj
VUp7MUbmc7OZjXtLdcx0Jn3br8syWi28MhuZdChWGgIZvYCuXnZs9zuHyg6c1+1fDtaKGtzRuGcV
KaIMGTpmts6aDMNVyHSQcq4bTA2cTF+zPG8sF+TNSLRnRJ08xXusyoOvBGupjWWbPzObcsk4EisQ
bQRZnJ/q4Gp9JBZJZFUYlI753fHLr88n4zSK3A1aq072JN6fMoWbDTEu4ehWhOzyr6KX1LQOhMFE
UPXVTkaPmSuiRMZvXIbdmGCpwjxjckOVrfJMoWEH0vkFEvCO2cGrgbj4sSnQ3NdUPytrQesYnNtn
EbmEJfrIZpC9Cb9PyUZie8MxKr/EIUmwp+LcSqFTpmydAxfUJS1Hwo3DgbxtLIE1KbSj8gsaimpX
soRzzkA6nf7XqV815vr2n0UQTTuEY/+4LesA55EIlckWmxP5y0N5UNlhtVdci4F6Gz9eICU4/1oE
QEFxetA1/9Q3O0eqH0Mn7THoNWE9dx+nVZa/jM9Fn9X0DgQyNNQGNsAzjo7IDV+m4GH7RLc+A0Z+
ldX2GEMt4YAgfLV+n13UdIhS99t9CQx4JNLr/SHwEdRFPrFXz7NxXSBVhHI9snAa2WsTg5TMUPHj
BsQTpPxppf1eFct94ai1HtLo41rcXH4BGBZZSYpGiZngPEZefKMzqlGuN+b4/P3LO0gQv9QU2AxP
pue3YV+tzuyAsrLqeqPOSultrY3alo4ce4LwOqrb1k3UoA5gsMhwMUVmCvKXWclzZkq3/MLyEdPN
y6B2jjSfjXoJwlBWc3zJ/cbnZNmtSWgUlotezPodvvP7RnSOMSBR7zltt83J8uG4AaAUCqoBJPtL
pjjeZuZYH+yJEqq2pFr06isWhTwUHOhk+MDldCPuK74Cdrl5FySR6DdvDKYJZ0EW9I0xonaFltrD
UP9sD9WnJ3N5Dfc30yXkiCuidxuZiSKy2HjtV1onO0RSesmJqkRyeV3ypLgQxkhqDlYgPjN0Yjhu
tQzp/Hb40s70EJhWmiQ+XWDyWW53FRuf0bMBL6F3We364UUtpncebX5qYWCNxUSz07wltMxK30HL
zVqraYtTq6HvKACiMNWRrq2WKO2Q2NGC/Q2Ffgp+MdAKXIXZk8D1rnhxFUBMDnWSAtoRKdf88crv
ndaFR/y5NbUOhG29uA60W+KRHhvqVPChSYXoZWmigu/J8RePoI+t7uNgbIAz5ulBnFasK/Y+GtFx
nw14lvZSVzlcwCSC06gRyCYQPPjlfIbRQWtmxyZDM94xO8KhZujgXDvsSYyPHcsOnzsg3MR+o6G4
iFgO2Wr6m0pzthddY1kRyYWa8EE5M4OYXd3SuUJ1hhKBeda+zIbbAkKTkzTM9KNc3G8bMWy2YxyX
rsFkIJT3+nYiH+vTdTvUCDcKCu6EEQrzoxUpTfEP5+uYK00xNMd5w3Sqvjy6uZA/x+hN7yXgE8D6
Yjy3ciSkI5u9FreZIPLL2QNaLsA/FsqDWfrTSFPy8/ulA8R9UDtn54j5c72IaPkJfUkY0K1fmx1F
UdH3J6ewham2jHIemxROtxsaR0HeYO7tMVLeXrtsEggmXNhsoe4cWn2BKYtsR2QCAWdll5lwV3nw
i6rpAAYBfl29c7Ltoo3fwq9IN6BTqJyGobCr32f6O1ffVhOn4D0sdRtwmXVpEDdQLRDt2FzqWS1P
Kv17aNUV4k3gbYnqtU59WU1yG0BKZWhpLnotsLla6iv9Bh+YYzpp7N7orzliiJI8o2wWaD2KkN6l
Ggs8nnm6U69di6QU3ZCh5BYoxBRCkDYnMWN56oR/XvWceYUYO6CF5jkIm5xFYyXGKNhqxbBM6TfR
2Wm9duiH2rdN3UBlBhf4u0zRLZw78GkFUgrKqz+uaisRFL2osWWlZQ0kFxy5lbLNVscmOOnMCakF
WHm0KR45focXgGevwcFXl3R0fgnXLyOq3ytUY3UpQ6GxE209ypgQVlQg7XqIbQM9LHrOkei50kZR
LI2J+sisZ2lyuTl2lPvX+RKYDgIrpk6DORUpmOS5nDUiauDUiWd08qcTm6RxomnpB1W2lhz1bJrT
g70lcn8p2d4rh5Uo7NsV5L2hpbrgYVMQ6CRO+5m6RNQaYelnPvADkociJ0TWneASFm8gv4iDvOUR
pqC0a/LJzvbwiCDD69+yH0l5o2EK8QZyVhF4Nr5rEsu9DeQsJS9gEWcg2/FJ3m4YpOexUS6+7fI8
CLQKQs3CZXmUPDkh8bX9r41Yapv3SvOiZNtm5NnulQ+6URQI2TxYNfzM8EWxUDYWkoBXEK0L1f3F
tBT3oNplyF15U3Om/vEYUWa8pOz6JnLHCxcW/1sZFrG+fPYSrPH9AUxqRmxg2LaLRanZBI3nRcKC
Y1sBRtN69FXljRJPe8h5p2bvsB69KMB17BMFioVyMYVtLmFBu1HGoj5mGKVoU5PkPyjQMsFAOjpo
q82lLpUAJSR7oDCHqKaFC7/H+Knwc994ntqDch/appuOkFeRv4Lbpcis9ctbF94DSNjFUu5Zv6p/
Ca0LY3LfHy6AqdypUjKm3Jka9pb7H/Mk4oUO6loJBbSOOhdp65RixMwdwQgJqOWwMWowRdgE4UpA
DvUuqYaOHfiEGiiTjL6a1yUDIu7u6NCaFomm0J4Ek68H9IU79TADn0q8Pl4TPWQSCXB83C1qSU92
Z30dDyBiOunethzaz1iaAv28iYliZrz3HIqkpb2OPsOsX0ymCnRVcT36GQ2eTiVEAjbCdr3dkiVO
zktyQWaVBvMCPI4xwbWaCPcukYXax9ltedStRdPvUOH7Ioay6AvNVrKjiVJTTH9qm9aB0x2i0sSJ
LcZSruYr5UKzI/TT2CYK3zgXkUDp+kDD3A2TiNga/ef40nD++o4I0NlwbCqHV5wERfeZqCtVNBMr
vgUlOnW5Pkp5aPUYYHZE9QdBJSmL0FBhF/kf7c8/B1j3qb3XGmoqV0fpM+s76kjc4IPyQvslSw7Z
mGDfClV0X5pLMTvfrdhNul12v32hITVb2WeLg1Qf/2EnBv2DpKBleqyxIbWd2GyFTzKmggXdp9vr
U8A8/qX77lcDt3pL9pd6itIkk+SPYkmwn/p0kO5xwZtqcjeJvbiUt8Wll25/7ERBEiu9iex49zak
ROJ4EiCPMYAOQT/9DnMaWneN9kPQQTF/zNq5adcAH5MKrKAKVtsmUrlAapQqBgbW5CYY0i+ZM6Sb
Y67MQX6X/yXdpJXBrUZvzNEp2BlcOgTQNLiGL10xDYrB+2f1RRwt8+83jqkJanW4sk+qEMDMZSAQ
hofHdvlJrkWyMpgyC4N6aRDNcgc5pojyEePczk/q4QVp6EmBcOBMn7D+9n0MuyrC8umV73eO78lv
c12GbYECAdbkmGeLfb5wJk+6G/eAP99NObxY0aJeBw9y3wl0TM7pXNv1vqrq0zGmCp3Wrvjm5C4k
6OWRRMLz7CKhWFj+XVND0IVfLXaSNIBYBN2PMqljVV79my17+OK5ilkKywseERlQoGufohCugNfm
L/yywQgmKsT4RKCOtBX4Q/NfYlrzPapGnw0Ymi5HU2Zwe0ClU+af7ESG5S41+FfJPfe0ywtCUSBb
A/jJHFM6S6YHGCrzQYxXEUgLb8qxkR4rHfkxhceCVaq88zIGrMW7PCFybEAChGs1YnaTJOjaU/fx
fXU6O2mjB8N9U5VsZjXW7fwfA165dFnoiGDZj9htiVyDXSAhYzVm41YunEaivRh7zS+YySDIse2g
lPwCRwXZoOFWjQGlRYsHn5Ykv7MFhAVcxvj03VkuLIzNPC68Sbd0+62b9M5v0hPsVUdFC0ikRfUf
CdK7qurjD65qohoPlA7zZOqqyzcEG9cCk19FbRgcmyCrmHilGWxrsf7ycnsXZpFaZFRq5ziPayqM
gFjcJHBupJTdBtyo8Z2SKEsKEeWWks13RnRpLjyiPOoHOq1L0qKIcNpzaE6mJGTQuQ3YAFpSAxTh
fVctjGH8Gh2OFr+GHtCe8KtHTciSFRvnjRyWPC+qtr2kdjhGok3cxuQGvPobVxk6E/kvU1V5uQZw
fdx0ikweeIWc0xxmBQ6afeotUxRLv/i/hdiDR9y/5RKltsvW2IBLGX+gMxzq7ZbIlObHd5YsymMd
+IIrSrPwAKSU7ib7IMbUj2ZOJWHlaeEneBj63yNI6OeJm1xBcPyVRDYPcXFr2X3WgKDehZKrJIXP
gl00J591W1L/L0xQelPaV+aYvU0iSDyx8+Ah2aGttX2fyePqMCza2NH+vvYvbycEdqa9UJkxmfN4
NXFjwAJVDmyb1o7tNg/ZaCI+zkRhTqI4PjtoR3+PwMLlcz4cJwMc2+ZgcvpB+cgrrN9Uq8VZcWWF
+SySoNhcluuzbVjMKKuEvg6NWa+2Tpl7URDUubnZpkGin9WKlxCnMi6bMGi1FiNvTLqHXOGSs+Oo
Spx3+hLUkKz/s6yRvuExfQVxm99L3GJupRmkw8fLJ+O2dLGGxR/eaHLH2H9WAMWXJGhOa4cb5h2b
xI/GTXMDd+e98mvPyW0y10QgYdCo0doLi0Kee9mp+lxKnwFU77LUfZM3tpyVZnoCFhzu47nrBWf+
gkFH6bpwd12wzvPGJ8nRkF6DpsITM4hTgpG5S5Dug/uCN9z2DJKjdwm7Htz3vZVa24IEmB1np/vK
Sm+Y+x63DjBKRKrTex9IDvHrbbOxtBGwZPI6K6807TZoQTogOIaRHLIgy2OSYmXGp34ibEPB7Ccd
nUO6+Hxflsa+vam08GES3gv+M/kKUQYUR68vkolIubunmiI2b1Z38Cqij3jWXQJWboOqfJBBLsoU
4e9wZMuJaVA6cUng/UwB+RN6MBni3zF82UUtVsxUqUg/h9cmFpLgKVa6Pxk8TAoEQH9JIx2cT3V+
+POfU1BWID2I9zoef+9I2EDACNhAFIYlQYst66Ggf5AwEo0saWXWBHzqk+hKGT2N1u2eHrglczdI
n/lS77QQXtaHof5OTZOs+Etwz+SdiqcmFrNBEgrzjjHz/HTkAe2qUVEr3m0CEG8uWkIrjogGyHL5
6ZaLODZKPNRaf1XCPFfnJ4k2Fs27iFDLTO5BzAgmDaGk2qGu7RkCXaMO/OprX47EpT2ai1A3jKOu
aizNC01uZ5on6wxaRwVC8tsZmNK3jNlh0cPOTIjRhFx2LjuXhStEXK/o9mrIxeRT5MC5GzVT6vK3
Z+pQGiXcwh8U6Ve0hmAc2BwxN7Eu1BSDKWTJbyQMglGZ3y8NbwZEiX01C2bGJXYk7VctV+aX9JnM
wqD6IED1J8I4rFcC4C0fv6NTYzOhygPbYavwm1PJMO5Wo7D5YvlayKd8zw9BtE66lcrFWKBouMXA
/HauRRo/XWhIqXSGki60982dOo6gZipXu71rMMb5ZZEJY3RYY3mMDQnENEtJ6RksQ6ags2MyXcRv
j2Ih5YR+PEiUMO55x8Ejx0ZfyUx7mb6sl/7ja630iooHaFZoMlGtUNK1ffAO4v/LDqXB8/whZyGS
GeIMIYae+bJG1Wj+Jr9c1h4CL7kGmNn+kmwwHWa9J6hliblB7WhFkaQPHRTBOm2GI3euko3dO4kw
lJdEiET1OpbuIGJwJ3AkzXQSfdf8E2F9vppmj3e8s81TUPsjU9mwGgOJPUU6CWJiPf1aLdBImccy
3WEbMRs+jaah+87OrOniNl5vvWQZQPNeRSTBuJoXKTBrAb+8XJhRF6R54oz26zY/j8IuN3yQykuo
63TApAuYfOonGdUFYTQvMttPD8N6QT1RTenKg0s7PYBX8R7KaN2u3k0O76K0oi5naDXiZrrCBFgh
a46RekTpNic4R5w6EOD77deV0lhimwEJyjcqTXu56sevPu0Bked8Qgh/VDmar35NxKaOrfABKBl3
lTIc/iUhWsFeci0DtYk4bNBchiPMOWSY82NEz58QQnQ1QKRHsMej6RHWH9ioWMJY93pwOsn1ANtZ
S4Y3LcqxtlnU9VW3OwzL+yNQvDR82Pd1ZynjEfh6NvrTTWfwJvmh/a9XQQ45e40nhH+kVi42J5JA
4z19iqfqaSWDGO6Zs25rAZVt5utweJAK0FxiPCveyNLYdPb0dgrdv2EbKPwM0pAXz6WlzATWuQjT
1UxmQ5DXndbrXj+BUg+uS0/tIfLZ0Ue2wvbb+fhrnYLGnV05tPoQCXj5ofRSj/p9Dh8sSlptPc+v
LbiWKcvlUyMnWXZRQP3ZSIryTl5X/iMiOtl1UvkykMI74Qe/S7kKV3hOCwy5bCL5j6eE0QC+QsLj
bnRlFIrlyn9gFLLL/pTvRdfCXcqw5TRrdq6oj1z4hENeoDihGJm6nVwVFLiclt9cXKUOUmMFjbPB
IaMYpc+UPoOI9vYVZL11ElzLXKBAJbmFBuZUbJ+y2N/WJhFobHMpHGRD/+z6bi6VZxSgehgK5Pxp
XCHF7dP2vxy3zQApJX+qe5zKYGQYGmPRfWq5lN52e19womuJWAWbDJMd76mWantgmEDODTnx05oQ
tos9Gm3Fs2rHMwd2PvZrItLoD7AbFQDoOiagn+9i/pMbzT/YKt6XNhX5zCyDA5PJKczWJWgLsxRz
5JkMjifuk1OXLC+nttJXpVp2mMHOAlg/KFvLAgXFNnedXLkzjpFvXbBBrHh4JY4PjOYjW8ct8lkz
pb4pBzno+pVGqZP5NpjvQcZzXNG9QOW1Sme/GBdj4z4trgh9PDiZ5T9LGhpfpnNeHai91GDD3edG
SKDU9wGhisCvi0As75uv4pmFJwBT0qJxtLjz4Y88z11LlbZUwgQBYA2V28GBLJCn0HR8meNvWpeN
Xg3IdOzDSchYWR4X2awzSnXOtbuaNDyqIhsorP2N+osacu9dEl0OAJQYY73nesnK2xSSkPaDXmp8
X/R4vJGynMKAeA3dT2heF82Z5r9A5GQD/rMclEPNnMiMDEsdPipHOJ51lnc9RTAXWwE84CqxKedA
M45f35Yyx5RwN/mt4cpzjELIKCxmLxATeYul29+OhqpyNmxRccn+Rs1ttEqnEG+OxD0d2g5tOD4E
eg7seV9NV4DAA00u0rj27FFRjBJqJRfGl2qmxalH+zlqggO30dsBUYYeUmlD+Zd9vLYvA7UHL/gr
gXD9mb81o++JMBXeSY7Uwlk+b8QY3IdPlSnMdUDGMRLzgz0h4D1cwMaK111ZSGIPuSkal8/3g0bL
ImrSiS0MFrFvs4FQuNIcRs8UGs7tDpi/6thkPmPdS63nNFdCaFDx8qvwnBQoEMYjEN+jGmaSCRZV
S7NUMsE7WDy28zj3trVejkJySNRA4b5Qv/nVx7d19Gl0lnPuDYXOmgE9nHMoTXU8XYYw5tygptC5
rLG6x8C3hZ7UUGo10ckOLkp6/osH6LgfYuN5ko/LYETN6Jen6rHAi3o2dPrIU3Bi5TpOmAKwQwj3
flbOpvI5Mzvbig2EzePShidRRNB9dcs+zej8BZ5uz8LqvmVqpkL0aTA90FdK6esdEQo4ubE25vsh
kp0QladHABlWqa9DkOwizTtGyeJVkdm24ds0ZIHGdynqqY4+0PiEgAnsQZTbl0awNNjZtHXOmE84
o9jYNYegFuuBXfO7Fr6VuWTNHjn3xaRh1LeGSkWvYdCtXbjpIBBPHxwIdOLWSgqUk0/zq4nAtqUg
oNFeC70yi4/CWXJPc/TyGsjpoO6tMIubGMy3aob2Jy8f4r7NuH8s7vP3/UO+93TlzOvNipOA1SOy
6d5QwUwzIW0+Yx98mi1fmTS9BhbsZo6DJCi0HhlnPpfSAsEHC9AUZrZPy5/5chdQpptxnMwXuaem
0YHnbQgL0RRdufKBPC8zXp4YQ82E+VjxWT6eID4wFqS+05F3B5zAr2Z2g7UatUK3nt8tiV34rsIm
HXyoBEaqZaqvDaQlG7yTXLlVUN3n09+lHwUephnIzT3dMIovORHa3Lt2ZiQajXI/iF/ou9lWuBZc
4vIx3DJJugS7F88QX9rpxjXKaeCWRJ5a6TvjnuPYzvJSn8TTc/7XTTX6eVDOS0rvyPdieGYl74YF
GVrK1vCwwqhlFzVb24k/1kn2+QSMa1TGDqSm2FtHuqMqOf+moKntxMGBI60qN8cj525SJpwGe8Fm
zSkU56HMI/G3NF+jTd7hnAdzylpzVKJeuHSO3VpHsFdV/SzatAHmk4Y5Z2DhFpwet4+K7w8WY4zz
fqwI5Hws0ZESjDdWjtNaTDgRWixb+9KIuMoPehK93L61IXUoAuvGlRrvL5w4vFYzEdSXtOfTSux+
GnW0eWZvsBzmrQfWuVyJGFBynWMbvObWEWcV+hds98b3q4XQRSiP9wzyYSv3bDd7jZcjLCENdHYf
Ga9XQZpXhqr+v18+5xLD8TXV3jTycHemiZWVqqLv/xxB2R393mVcX1z1jie/G8aA5byi3Q1cTKZq
TffOsP7ctnT+khMbFAymgk3i6VCENVTcX8Ia/ws4NAVOQD9KVyXgdcVPGLcAv6t/OQ4KcRkcwhJ8
BL3SHCfCdLBnmQPvrwktARFUvkORyrF00rMWO9gm2dv0Mmc0nMCxRTIbqfdiFf4Q9Jk9jEqWzqYs
S8lUkKNSFqeXXTJ7JBeqKo+gAoZeJEDguMr78UxpmyYt7e8H8VLKjys3kfiUetN2ngIF/Rmuihea
qzFYGuUGPR6BD+yNX+voYJW6cE576Fj0hbjCfZGFjVEexJfo7X0q23eob9yEyEBJttBKAyN94+h5
0ObmKfI3xzlxm3+8IPAwTc1OVpNxGHPd+1tvtcuMAMQ2tqOSw7DcBweNBjZ8cUYiRqvLfd6zmINH
Br76xEdHK7K/AF3gT0dim8N/I5iBuHk6mSeUZ0iGYfn7W69jsJeaGQtiRu0AUUuusAtu6TSEiUH0
bRthQjBqKmvM3bgvE83d7Bk7vpcAl5pHUKlCK/ppJS2SjznMaThbXvUZ7BVURadeRd1owouOGBUC
d/b6JeFsbvpU3AO7mGl67R0/FJqQfrkGGvL+AWgDYuYZOcqqC1NbHSbn9Scn75mL0Ot/X472+Poa
JdbTTYr5S2iAl4hJZvxGZhYICaxisSKGmDfn/C3fqVkYNCHqufv2M/EeI0U0f6xkpLtDIDdtoN+b
L3U9AVnz6dYO9fekwa9ZNJj8YymesRG5aBr5GcJ1T2aqCKG89Tm3lBSDnauWZyHKeVSI5v1UQ6px
Wa7JXr4kp8Bpbj3oYpSBX5PXniva4hK9J0oWsnEDngX6DgsS6qklC/1zdgCe3muDq5UDl7LN4zOd
M9AEvTJPmTaehq0jxvOgnxrRsjiL0dr9AdaXq6B+gcpYMAiRxSXKdY0jhHX85WSGVt+UvBvnHU3L
T8I8X9qkuTDQtXsqoDk1VPCLlHQjlpV3n1MZF/8AsZcB2C1WNSOEU9D7t4uWf6qN1dC/eDj/7aig
MhdrKGEQZuXKlwoIP7byGG3b/zclfuoBDYDstuoCmz/p8yIPxzOlsU5aSOeri50/ZuI2HnTY0pYe
RNUKDbWoIDTr/8i1+3v1Vcq4Cj1L+OJ9UnyIju16jLl5w1qnBRx69p68tDRwDbAr2h7lLVzzJF8U
6uHL2R3cu1A4kWHB3OKbq+G0RBVRvOxPfLuobjPKHHFX2/IGkVx2oyElpHKUHkf6CEHRrkNKVOFh
7w/J944YZYScmylUgLK/aMo4Tsa5Qc5LFtmksn6vkvjrXni9rIHSVwljjEavdIdyRRX4gSgx+1h4
pShuhVgrnGlWZNFXktU3Y4nENlRlNsT7dCQwIks2+OifHCGHcJ5At89CTEAXiEuKXeEVqnz7jZRu
0v0snwS2ApZlLclGRAt3pHv2DtwrBB72fC9PyJ4qoDVCMEY6cK4IDIOZAtw22ikUGcOSTQe2EsJN
gw1RY5im1n2pTqGpmmNNitz94NPlfhmAFl9bZtSt7jijdfQxojMnSF/uwA5qohmNPK8GwB0zNZot
Y1cwozL3RRr0fVrAkva2oYSCC2ZsOUrO6CebCm3o7249hThY/3qEF9OuM9orfsL1myDGjiDHYBhf
bpPYuUSHA8Pzl67A5TGHOY+oztqsoojL3wd3yMeT5lrZmLzsM9ERYN77VGONii//Ls8cDupx5QRj
up85r6PhdErZjQGwCS6pur/RdIIoqtvjnwrLv9ahbC/XjpT5x52PvPYk27vRpFeFRNbmgNIjs7/X
XEFpDbwlOQ7aptC2EBEpBwY0xjF4zkTsE5/uBcQTsc4s0pCs5tZKnB9ly1rvPhR+1M/uwNHgnRJq
0bWKUZkwA6FYOHojbJV8g46lz0q4OYsAjb4b/Kah0GIYsvFwX3sWTLCwAnc3BGxwFKKkRIeaPSAl
AL0m0sYQL2XNIob0xVdGjVX04PLvAPvdiBKsUEMy2rWPZ13AVVx4Zw0ANbxVlvIt4p0mq6Ww7Bym
3mHP35YtEzsE8ZEhdiuBIk0sV7xC8DTRHK6FEd9Ddj/4NsPzovgAkJAiDilT5LZhAfrBaf2V1pNN
Rz/mj0IMj/D5IphrgZ5bF8kh5ahZL9JWMf/7VGJ4CoFTD1G8fPFaCjer+Nv891iFpLi1GLXU/CFG
9BhForIOpvnvsb89FjW6rNdjFrdvIMWEpuPWWBuuSRnYkqOY7sWJMXxgfe9KKsFKGgO+WV8xQ/Oz
4NtVWHeAQfP1/Tz2vA1nJ8leSmv9TAdFns7+GjbN1R5FiwlrU2kvU27BLRLu5+awKhgYfHk/F7h1
FicI4jO7kOHikGOEGxyMqjD5Ib2owdEmmaYt5qA03AqRe4QVgLsvAyKaN/YopA5YL3s/VC8pf2p4
ZFOQ/C7OgUZxsLRX6xgKMA5Q60UkPc7glHnjKYgikcdF52XzTv6hx/qyHidkybD0P6BOflHQ8fnn
7VMYhP7Q+gtBEvur2t14o+CrFkTw5eo4z4h4CDBl09QIlhgtePQ/ly3eAkkkTKB14GT1b8Pw2FKO
X10g2gP4nG0AjMACZ4a9QNdUn3qTKebyB8lu+JAEse0aB7y2/9wwmX8D/66v+yWPFJxloNm641Br
3zIc8L/Z6m+QPKtvMHnAQ2FPYyY3KVP4xPulWRVgzC/TiODhZBrH3Je63VLn69XZR3e7yq0v2+cN
NJ5rdlph9KT7jAbpIsuC229CYJHJ2SKcl4S9sgJsVK0o+N48fFJwdZlwHZJbXSN54Qp850qcDirU
tHwBUeg5JbJwjBDycyCAh2eVmTKIaU4tAOXo8GhDpmcIE0EPEJlfvCY4y9jeSlWLjmFM018ugwO9
HRwv/JJyJliIfOocfztB/TM2sQVld/zMqdet/WpyjMJ0yobz4YuIn6A6Y6pSE1pZBZWAfo4nN7zq
xdxJhTHF4rW/BECgWdeUUbnxDoA9hxrZ+kxGFGReqU0sIFk0pKrU/6B4uVqi0ppug84NnImmmu3c
CdII5hJ4SeBSG54pNq6bxwOFAhZGdJfrv5kJM72MM85VY4jSt3+ylfN9u5HKG3BBmUoPjwEZhfWe
5swfTG0ZNIy6/E1LhCbomy1fLimWzAlNLKPKlIladxXkQPAro5N/CN+HFUlRsLeMHqXpRNtHbv/l
Npj2n0Mt6vVOrUW9dPMjqR9fyiyCHV6rNI6IJfbqG6lblAmaG30LZKydlpFP8Vj+xNDHPGnF4zt8
Q9K3GCC9b83yLuIeCj/trwKcZUNkQCrrqZIiMiG/HHCDvX+pUG1o6+ihamB4oOmDX9Md7M6dV45r
pET2hNzB+Jt8ICSCXRv13YoZlpImUuFG1RNLS0kL5TKMa+ZAUdx0tRhaCwqMTRWkMGnK5dEEYbMa
/FniwnBgV3PYTQ9cLfcZgHllqYPuNeW9bDBysGVfyWG6UFS3GAgSJf96qAsF4x1eGDbJvMoerVVM
QdXmdTb+Gj7fooUqnlud0J0G2DusWS87h7cp7r3wcdEmBe2oLtSiODq4F4hNREQCnUjYsjP2C9qF
UT9/gMpb4QMG58TEgvb67BVf4uQ8RO2U5l85hwP+8bqnVuV7f2UMAnr7xQbgy4iQdtL63+MlOtLs
V84U0EjzECmRhqRgeXYl52tPHP8F2lhf+cL/ZuGuewjxosmE6Tg0IR3ejzU0YKow66NN8wtKAKxK
75jjvO4mtZxWRU//M4bNTX3+FukiZ881vIbydokHUqDRA0B17ZN5w17bn8J57V3F1PJkfBkmL+AG
ltZr3EgIMH1JFXQTDc7gr1LP42HbQjKkAfKvwUshjG8pvA7PlavsUUIJWWSfc1Z1yXFeNV+KOClL
0TQekmy8KMXpyQAwVP8mgfJmUqQbOGHq64zlg2Foj+hAUo6R01QypknkBONbp3lc5B6+6IrJGmuT
p8wABp13YMNqxewgUFW0ohLKPUQusUzdomcXNmV9qbpnTGEblbatMb8Knltgw3uRzB8OjB1j9X/Q
p/5bon5Fq/yf6ewvJihCS9+nrU+F2Q/p0n0msRyp1ckr4LXAa+HpqxE/C+86KI26GApPZMFU4g7R
r523hk/Hue/MQkNMLz4sY7zNlekUQlFBWsWE7KS3ekDrYGx3kqGzUOmkCf50J9KpzaBAqC0heh+K
+u4PNffTtuPDNfb0JFJAzhrzfrRBY26L3nWH4x98VKiU8vPfEOjALqLdADUXTuLeXk8PrEBtAmaD
gUuMAsKYMHlhHJDPhxBlVUsoc3QdrVk+P2LqC0ZnktPdjXcnrYcWpgQMFDX4XcUoEhHufGqO3kuZ
MXX1fzdnMhpD5k8Ph2q81kiAncIULnyJ5qr0wiG9mrRBw8YaWM3R+4TIkB5fQxCKTRSDaApMJaHL
cPXp89VmkMWpaCQPq0OshB6gj3UE1x6Knf+S7NY5VGLlmtxox2yQ0QUz9DyDvMQM/sSr2dz2ab4Z
uCr/lGHhU5GC3oi9cC2hfrjW2zjtRusFESDYJAinisYjE4zfPM8bzS1gHepGKKYaKrbFFAkfTT/N
533JxuFDU0MOgscRMm1cXUsnOZog067rfQwA5Uau+uYg/K6UhRsb3km4XTukpj3jRtRmYU1eCmLq
IgtEwrPf934qtSW372eRJuW/LEYIuKL0jXsH0eZm4keTdkHCv9GTixAUtpGgLVn38aLMraUIQ4OK
5R1GG3+Pn9dTUufvllQkKstiUNQf5p2o1fcuHqNHMhFzUudj31VNScJtogd+ksh54OUmuCuO8PzM
mZYPRap5N4wqwiywtPNQFTbd/qPdZ8HqnJs7OJ+Wd6eU0YbbzqVUCoLxdo+lwvbISYzQT7SyBID1
iH4Lo1wodL28c8J1q6bTzzqQnaCQhBE7nwmWz+CxiyoX/kCsQVaT39mA/VoyzGgN1s+4s7yGmDKu
UNu3g9WI8LN/UxcmXw+IZU9M5Yt5cMWEEeOCOrYP+yXvuLPY12nwaIlaSqrafvlBT1PGt5qIAEWr
0tRHTvOVMVytwJyczZQMyh2W+nIUsVKf+DdRxw5TYdBbhsljN9G8TEXOOPujh9lUWgaurbCGI1eK
s2JHXmbAY+g5ozz27UTGyFdpT93e3VJsEOuUJOYOnEsjF7H9cKoArZGqGQvSL6r6IDY+TFJrZIcK
yczXP8p5s+EsnsXoBY1w/VHdDvRio1QCY2J4ABVBOwk3I20nHH70jZ2O5u+dPxRA33DWoUnepovT
tNtPJLQGBG5LuC18bDNiNt9WVYsR/c74gFCAQZnJZS0fE04m0VU1nt1M9flTrU0YM2JCJt1tu4p7
xTiolxkcNNENysOPBwAg9DDCtjelnvdlB/U0xS8FwCGJm2AB5Ycx0jllET/EoaK1vMn2phondpfd
OHhzd3hhaZFN/m/JU0QKA9l49Z7LvRkH0Y1WkQwlTvvBfixUHpl3mVi6LkzxEhKXIimKLkPmdzID
WCnze22JmB33Q+4tYb/DB/Xko9aqDdpJFUloQO/WohUSg3iTGdILNfrOm0MhlwKuQZKFpwOLbSD5
ELy2600ULkUUeSf2KVJRZNXZaJ/P1roN2CyNGaa40ouT5tr1bI1N9XXH591Pf1XiWYGSn5gdakpt
8fFmN/GM4Q0lSD53KyLi++jN/+ZJrcjLxCNcuyldVmycrEVL0c3nnpxSI0UCv1FrqtRvoTLXshOd
kX7NTcE8ZdtdxHsKM3MTg9vdusZ0xvC1o567aEv5HTqkCmXueCgHkYYTL40g4wFcRPBrxjbp0CTZ
CR1fml9CvGNFealROia1eSYvr7hd6v4w3gwYDv2I5RnyVzuCVyDlHRr6X0oU5f5pyGZaemgsREjD
gn5TWhNyjsz0AeLTvrMzrxPE5qpfuSAd9hpgnsyCGz99GL1LYhxjA2gbg2C3ZieAgn9tDZgmL6F1
TYElyVpGnGgHrHvwQw3M6uK/KB5g1kem98vK6NkMh8VpVvG/OrFUalxnBPxKwda1rB41feI/nyck
j65A1RZ216bw7R5T5raXZxraUImDFyEupTxviHJc78uERz/ZAqJo/ONuL/OuTf7Rsx5/1sDHrrlW
XimRheJ5jAtrRXsR4xfpkyDKrkAuXJHFhIjsBxOTSsSkESrDZOnrxh2XMgrLFvBqX7w0mEjaYBt+
SJb/Y4FlSwOaa/kIVeFrjGnFTvWYIYU0YWXCCXHpRN4GKlaLC1qa5JokGwxbCJyRPRDgAmBZOo6j
lkCHqHhojyJgts1bKKbmO5HxQmPViqK8L50LUf6r/F91ixfjKbPF8kJl6yxumrXrzb79nq/t7TLl
P76GuGWx0+MTSlGLQgoG1EVLcYvnHzpl5h1hgL4IAHld5CiHRp3cswyTTHQ9HEA1LJFMmlFjMYyd
SI1PvF0OPY3uUqZH3tFt0+oOpLRqrMxq1PCZSYj5clcEaPTEDJDc74hW8YGfYT4LsogJWQewxKv9
9RosFkx/oNR3wJw20JiyD7G5IdwKe1k0+Tbvj8/NEcdE8iImzl6zsE/egF8tZ2eyyhfz+RkRyQS5
DCRc4zeskryJxvAOPYS4DyYjJei4bvOICsNhamLa1Bb6Jb9UvgMqdWtqaU1bj1nlYDmoMfO3w5kc
dZnG4LpGnNzV0M5JVscAXe5EPipADxUsjUM313Diow7J7zgcjPj6HqifE9TbtAkEH+6E2b2hZXhg
jn99fke/AwICrqnudF1gDtW4QXjzXOrmL6LUpTnNzOONtmlD24UzWnXGB/yR5gvEin0AK/y31ek6
fnTMXZWJFHBMJgtvcHuygKPorpAnwQMz25qpj9/rPGHmrB0kJfb43lcTvlO7b1uhM+PjhPDkWL7R
4RwER3+/Fb7f0PxxsPdGsPA/aGoVsXAxknGNt13K8kG7WfalTL/+NasRs/SM5izAhaqG9npkcl9E
j5fizhLgteLWnOlPNbJfz+MsEv/4MyFc12G6kbo44JA+TeEkhPz8t2umYF8u8er4N7n28axTOzdf
knwpMGBa4micUX5kXSSWFy0BgsBUoaYZgLr4bVeF6/gFai0xPuxrtqPiEsVCXrxlJTbpy8Nrr3r/
K9xgQVvrIYqgBfYvpDmtorv0V+V4M3VOs6uwIQYW7ITYr6J/MVz7AQoMr1tKxQpxPbYWYNgFdbIy
OYEzXq4RQJrMIHyy4pzgx1Y3IuJf+NtoRlptKQ0LxYjuG/+a/mUakIbue9XcftEgBjbnArcnpXAB
Sa2a2xoTlNJRADCIDpMbvvoKVpfoPJOtdelN7QDDSjqwZFVDAcWAODHpW1VV3je/M81609jPsil1
EpN5ELE/Iu9ODqjehJW3ojz5H55beDonPjypYpWCx/M+laa20E0Sa2M0mNXUUpMIeAT63Sy/BRF7
qtYk8pQFu5ol7c1pusnNCewqNvKz46g1rkrodsUkOCiBMw4Ua7m2Vj1mlMlvM6/tMOU+OM0VDmCV
gzkb037TzGEPQiaZFyu0BY/Hno3yfbQmtpcdfijDIuWuANPdTeHyih6gL4k6PIFLVuTMGd5EDjUO
wL5A93+ECSZQfLiiQIzrtGnwrRbgRzg54B2ScmNlcdiZVzUhQL293nnrUjGbdXyJ12nYmXFvi9Cq
3hJSF//DC0cLLtYx+rPk5ICslhZuwheVl53P8NhNhVPow62XOOLlG4UGeSF9J8J0jaWSzLJyxqc4
tU34fAG0+M19ktg3TEZry0Uq/oWpjRal1J9oR7Zu29mWNxeyLd5sZ/7hrIazxAiHQuC8v78+pvLB
2KJlFChDAPga3nYJL7K5E8OlqHgCotVL2MN49omPbSPSO31DzaFWRcrePM8FS9vjI7lT3K08KN5X
VifpnGSWAiSkyGQeHet5sswh9TzyJreZBtb7PAIKczE4S1N/hHGthW1ufOLAtiqcFGLubmBlDHKa
ZbVSYcsbUhuS0IfUb+kdMyJkenw4PGPrtJRFI5+KGq8J32cm389Ui1Pk3UH+lKaiCgFOA6L+lbs+
LmsP+CXkMTlHKOkkffLvCH7j35Xdj439GUi68VtLiHnW/xBusV6oybDD6vjqCT7EazgLsD5P/9s/
LzdUu8oZHNKB/9LJcSlGZBErb5IoGNg+WSkForzoJIoHWK4IsHVsRPLdnN8jGuqlqLLwmnMQMXt+
de06fw2clRcSWwngnrpykmUzfLjIr6hUCa8Z0HCGe3JPmsYu+SQ7Qd2I+LxZLSOx5HLw2On2mEZs
9KVLhuLRh0J/m0UCcs/MmIi93ZdVHeLeyyFuFzRkmgZP6T2UZm63fneHProV+LkgTCAjrUUVBCPD
IG4h5xszESbUesPpiuTb6gnKBurNBv8jZNK25Bp8dL8NWjnkOJ5Isl5KHOtPxAsq8JaXne415O3/
PqcKXmC39nVP0XKwihQyAqAke49D5/1+9YmS0MybTr/ZLLgahLChUwN0/OEDqjXViQMaT/O9QPKx
pZphx8Ae/JkeEZAbmjZTjHsAIycebMPPcnSuijSNHFRIF/gPvZpUzVK18Y0H4PyPjVSVHj+TKZKI
WBmhALy8XcFl0mPY+RCupyw6/nph6xZViR3RhjVidU0HsxRr9CSVNXzSsyLTlEUTaD9jqD3ysCw1
KvmmLJSn9a7O5WU/85EFP6V9fV5O2MZdIC4LLTWxzxxqM72AeIHu2RFQ5Pe8Yf+zCS73OfPxDpAA
g0+fNsdyVeWwLA0qWfyCFuQUvPMuZgBXr6yWt+5FQR7rSbdxm04/UVu0J+nfm95rrEkRQoNj/l8m
pc/ehpq2K3Myd510YPFpoOoz+w9g9aFXk1rfFHTLRa+TDm7/h6756U2lEcT8EbCfmnV19cj3VaZI
63xy4SBc051NLUpbEKVQiLbnO9UaJFm/tWYsjuyj2BXKn8fCVJKPtYuBxvMDXT+Q4pvLniRbNQvt
tWCTrh5oJuCtSysM4EshWLU0V18j+AIuZkZ3TR0QDF4edobM8yi2Yw4SGILZhiEdmXfPKxv6Ytyw
2lkUrQGeWTWtfzr8KckElRc8r+ADWBq4T64BiisgjtMB0nFrTbzhGyAbzKAsY/ahH2KnVBKYTxBj
WQ/gJexF7YyIW0QYy3lFsEuXZNp2tZ1AkFiXVNzQhqyfoNSutLNnXofsuXMqiQHjQ0xwomdw9fZK
VPby+XG2T7CV7hckzmlYZeQx/HPgvstM8C0Jexusg4OPTNy1yFjg8O2S25CEqyhUxD9XTUGtmBGV
UIaeLJ7lmS+uT7C8nbnNQPWPa5zBEBMe37Yl/gt9seXMhNp7JhfgY4qEQRj2eaaU5PLspUPRaQT4
mlHoWrXY/kcwba+ChMfeRno/7bZ6Tm+7BjFVjaYFZM2m5WefGfW6bQFmalSbGIEJAfU1wknPAc1A
lQPmMO3LlKeyLA64IjzsRCxp/1X9ao20G8UApXUVwjseBUL18IPsjQsk34g8FA4rhTkkt7WJ8fJo
u9Dm+4hAmU8aTauF9kgjMDy8bqxnx8+0aTWld9VUWxQm7cIzFpyY5NhQn/c7Fk8tz9tRZRIF7AtB
saqeapj0CII/ySo6fuLN/2JmYeqmIX51Ydqus2+yoqsX5vX0B07mkWMiWxuEfggu31fN9ADDoY2x
5C/QcmE9OL/eo6hTbqYA3w7puaBnQzaXZvZ20fV3EOV4JLO/eqyB1yehjIf/Pd4PJbJ9fqIvjIsG
14CNhdQJlDAWmnGoE0p91DdkmFQHNY6JC9B1+AicFhEInJvNtqTQ+5TH04VADAztkNX0KKtGegdQ
0X3gB1Zv9q0Zk7+GeCcqdwrgSTVuQY8hGsW0L2jRYBmVpzwlb+VT9LRcvxtwrKtjTAofv2YHCNXC
ZESmvNXgRFtbbIXWuqmCPUiyQkY3m+PUp2otuFZUopsKMOICLOgIZzjutFynlklJAUUhfaH5jofZ
MKTH8DvnTG4WvPE91rtbltPZL0YH5/O3yMVfFpgNKlkz6fOAJV9ExUFAiQHhVc5NPmo58MuUTLTc
fqiTeYGMcq139MnqVua2B+z8mhcIQPhZpNmZpOgcZuo3MObk/YJBO6U1kX7dkVvjpMAjrUbDFbS+
8ZmwJpwN3faz8HzSL/EA7omxGda/JnibwfOZaMA+q7KiwX3Ys3uk9pHeS495BiIHFIOJSgHM8axK
iRmeDXSnQ7u1xzfhOnAYZx4KVc0Mw8RZaHnMJvgXYok8+y182r+CjrV1F/Z6HSpW4pBPi1kRxM8E
PWVgbltikGc7iTUoxdnwfEWtOS0rkD4mMvB0mBDjwHuL8/3O87Jr3chl2Uxh4o4/hwvzbrHxMB8P
O71Rgrraqa5pfSSXgAIe5FkNl0NyD/0et6uepR0dGhIBTuJbe8nQ0BkTAQKfYyruIOEhp2sEm4jN
n6say2j8UBw2v4bN6hG/+DGyLbVWym2ybfYXzVVbfLpzOV85P/v1ZP5nM6XBwmkF4//CW4yPb3S/
Hh4j/zvskbPQvuZD44HjILe0U3qfQi9kkr9kIrAzWSyBsI0sHXUhYSJrfgq2ciqU43hjNay0Z34D
gUhjnXfxqCwziu/PVa/x1SkNjG93119SqIebtf99elj8xjNxUpfQiPA9ATj9r2Hq0fOP363hX4VA
VnNoTunH9Ko7Ag4AQa+8FnCrf5oiTLfm1Kt6EelIRIeS8q0Y7Tvn9EmD/YgHTvj2DYlrfhaAtubt
gx1UXoMKmWRN36fWl+5SJPirNlZmagqGw5H1pwLZrIIUXzjk6FjBcr5TZsXBIK9c13+XOI9kFuh4
bpXQyxAhCwEYsCCwlHDogIPhZp2rZfWeK0asyl9ACBeMoX175vpVuq1AcupKaiVvquhIkO5NIAGe
XJkh/InTx4jwC0Pl4yse2ZlfSppLYcfPp+lE25EfhskiwBxhYjrTPajVM+7uWx0I1PJI/YMl7Sx7
93VnjV5TY/d4lfOlJjzfaMN+2fvlOVxUYqQoDYOPVaHAEV6HSmfRWlAAKn9EtnEISrdgNZFgjzJb
JOPxZNGLM57MipqWgot1+rFmV1bwCkWc4ksdAFxxQ/0y0zQl/7zypd8ScrPsxjw8Pk9AEs3jLaHI
TTGq/tXfCC76vR54ndZ/Tyv3IbrHGB1/yJRrWK/Cmf8bZ2YBIpdsybpXrBf+6mMihidLiFG4gLnt
cIFLa+0nm7X9or5qPo2sqVlD6CMS3/MUGDkI9DFZ3sTl1sGRhKWirF7HOZfsBWuTRAj5bpgHClV3
GU7dQqVOdrokE8CVEQK3hmrvRvPeybYQcj0MuLOxcSGYKJskCcYTvFQVrMENoJT8V87n1FZptyTD
27ij/Z2+3GeNZnP7X6KzTliQK+rJpDc3ovCy1BHm6/TDUFEXiwfyWyp14nnsUWOXpyHZWYgOc9lJ
stEWKHpqDtrA8/Xab/NSbpHZ1WDIK2rarymveS4TsSUw2dHiMmO1SzaKjUlqdqsQRsCNgYAEdzeb
nzEUQV+8Cp37mqHQ4/dPRdjUGaC4kxsJJwM9F6RJKAlmuuBbAgnEThvr/B//bVHOXuply2WnxUJl
WH9l499EYMoXjhFqzl5e+EGc4UWPfKXc7VdM73yBlDZcJ1MER96mffS9egwiib4OcWXtTC51TIlh
dMg6G+fcRGzZop0UsQwC8+b9Cg29p2bzYHFqBoImCA==
`protect end_protected
