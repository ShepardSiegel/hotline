`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
noE7X8Y5XTchLki9yi0reMUrdEE/d7vmP/0KMNQoH24wsEJJUGx9X3VVb6rTJRPZlexfpPiO3QOg
0geS0Xrbdg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A4u3ecZMnKABp/TMiN/zSN9D+JbJbW9VAcp4FdP/eHPF4IzZ6mvHaGOMrrg+Mzt3MBuRBnB60tzw
EYPcE9eBAnvkV8t++QQvOQqnTqNoUnoHtYWxAAu21o+GT9lPMcEkqPjP/oa7CxKyR8/uZVlBhbtt
z4P2u2LCaQR0qMHGJLM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ccOqie00RzEoufOPEVpRV4X/iAK5NvCMRi/05fKmHAl3l2ESHXpUTLiq7ybYgXNTtAcTojMMRbzP
txhxkAdDFCVdI4aLyrYPeQD5lvSqqUnOmqoKzbjJtN5wBH/v/n7kIlY9ZXXIXYVfV+fYj583eKVS
Sm54UexCcEJt2uCKry8hipiAyqLNo/1NBVvKT92XHXPMdLKDwfGbb9MGDXs8xtFo0qfTp1K6ZPPM
DON2F5tjyWFQUZ3GQvoQPN9qQ51qgtUyad6Y4fGLJ71NUPaV7u744u9oj9W6HZhcbDL3ZhYXSJhg
8vQz/sz+KlMPm7Gd8Q3k/OTHh1qJHHnO/2kt0w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sB0LZhwYzB/KitfkiJGXsixK3Ndxnvdo7jlVxVUKdjCu47gTlnedKjBhkPcsTHt23xiIDXCryzhw
VuPkPZTGgobLluD27mXkWhd+C/lzP1brjRvhW2OzHgH38DUCUjOWCPKdqx9tV2+0ndiejSdMHvbl
54wrGzLiridy67UaLCk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YZGEEeGJgrAeSIEgzT200zHz9/Im0Le5w83UJxkpAGlR6GUk5fh7+jDFtyhlEAPnQ17k64U3JMM7
rwJuM6ABCakXvgQk+dgShT7uwafR2ZVlf1Blf0J1bwzJLw7FzWZKlOSd5j1G+UDlJMXGSeyOUXQm
146P9ZK3Vb7QOGbefh14hfC03GqeqbzG9aItgwFnp8sO/XvDvm/2bV4KEKCacyU5SDf9LCh8efwt
xtZTkxV9yEBjaoriwr6OFNadXkwebznGPK4XogyufSYOtl11xnk8f5qksBlFN1tHzf7BQivjLb5T
54qZH4VTXodK7iq6mVg315Hb8+qdyvW2POrydg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30608)
`protect data_block
EXWVyyGAZiIuCQZw0piEjPT5TQU2cqm/c2MFRz17JQm23KYZOMBrwSuynYgRF0X2AzUVdyboLjXO
q+0WUTN+mpyhdwCW5f+bfPv2vvTf1RaC7dHi7lqcR6xVjXovdJUJWe8ff/4ea30YjDdR12lOpjwg
L6nhbxI54QIHsI3Na507yTw256HGUBz9SuIF0han83K0nSn97g7N/CiZzmaZxujx5a/xR1hXfZlM
X4wrKK/mpIMl4/zFV1tC4Eyknd0toru0v3Vg7u7ZfDP6zp0PWhousSPQ2iLJlBkm7Oqva7L+VKES
0L/b/cjmRxiyiLWx9zel0NhNSZP6TmIe9MQKris2ZHzq1uB4AC13uUYKJj5U3uabMN4nLs/MZECL
zOYDNR6jBt5YK/QYvALvAYxKw+SMaQW1brCW70Ygh3PqYP3SgrCB5IcoqHUB7qsCvKAUUmpfVtnn
8UmVwHhfGVi+YzA/wDBxIMugQ2D5fr0KS0gjxyFMeU3DnmmRhRsRKDovkkI0od7nhViwbfwSdffN
+ccFAmJoneTJ2nyQQQQLpaoaCZiH1cC2xiZa/s0UOubYIULVdRO0fGC1jglReqhpcOVw1k7ymH25
lgsZkdz7wms7TUP9OPEoHix5vxGqK6s0eeMl7VMDKUZT1S6xdlg/eJM25LvHw0Zkb418e05Tr3+E
cp7DU7uTpfx9lGXbp5onlJ5GmNjTGUPjgdGbzA3si8a3fMw9WQXnFvARkVSYJ4TJYTFPP1iByiup
5TOj5BsB+aWrdd1LO5rttne4lxMu5fdXFV82kDeATl84ckL4vqgi2va1cX8V0CBbbQ+pePnNv+pf
gTwLs4MwdGIXM6HKYrtGCdDRnjMC3OQERLy8ddrBZNyxrTvOu0dfDA4bIkkTFPKg88p/ET4rAOjE
b2ypeqvl3mJckiDzRLzMdxXeBa3YXUDy5s9GMVHBK39uQuC5v0fcK5lC+ONYyThSCAeJZSMfkXTF
sAGTXFbCKIMfTLOvPkiOs/NPLZo4mh1BUFuuzR+XBFg0TKDWbuFwa2gJQEZGJfKQ2jecihx3UYlK
GdCnYO14R4LdqngUl5fBRG9WD0dTQ2F6VAcayl8vNPYBohEYNOSto4+7Z13UPJt7j98JTzBnKF1B
LT8UMnrDHDUu89v/6Fo6/UjqOeVNZbRyrWXBZeK0CLk/yiFu/8oFv/nQYwKx4JPtXXMx5UMKgHmm
8JbQWXDm26ZQ3dnwCkdcsha+qzeT3HKKyRaO6wyoPSktSfloFTAbZSrTHyT6IMUTxj6wjx3zvmHG
R055CwF9YaXlLKGB+XEZG83+Xd7+rlTQJZ9C/1aCRbM452VWG8b6XytXimRI26CZrebMg075mwDT
fRsmN1lozhp3abedbVcRaIrjrINkb5AB9bcZAUwQ0/U9BsVLt5F2cqG1XvH/FDMeTeGUfBVcPZe4
EEjhEV/vi1LP/kgASihoxkEuP5XG7L1sr4NNi1tl2Yj0E9FiO8GJIO84Wv+7uqDsbIvY+SkQ8tzo
6XzmtR4VqYg5tmm1pWwm6qdGzgSRyfW22Dlh0AdR9eMP1WJ3XiJntUOg4vKy/mEFNsAWlsJfKkR4
OJsg11AEFvHN76FADJg9jyAe7+byVDQEePzAh7uqXZ3kqI8HpB7KYyJdRtCGGe05um/mLE2HA4NV
nLu0yebvkNQzDLTaqeIBfVAP/pUwThdaG0mBQFSou7mVKAEpoY85Pe3hujyJfXT+3KhKj0pjcZFc
fK0QHgIavCo1IkgEa7FlTMSlWwqQsFf8qy5rNbh75XYClfeUVlmxM8ELAk//hHcyW7SXmDcPC9u/
6JYjG3/heY9d34ym0X5vSf5RMTkpRC2yWwFVd7cEmGMdD+lpByrBgUb5s5Jh9aoiSzEtq6oXu4ip
wRpcWC0hJLbW25D8QEp/4s3eIgQfaN4zTxNeTtDGQV6DMubKI2tPgOD9s5tirvfkuH8sbuC7cz7E
KzwuNHuO55MyCzlST6lohHzxiViXY1r/sZQtyzTCJj6ZtgEgmiF5+5NceS+v9lSYZYra69yBUsCw
hHcgSOpHOx6O04mNH0VlEK7ZILAhhdOBq/X8Y7HLel1Gs69FSzmV1OnXkiQNV7AS+qtj/3WDdHCP
FDk+q+qE8qlODb/+1TFofNIiKSPCiGmVhTYrTkX8M1qg08c3aNXX3zCD7p4pSDYCwgpQGSvikPzy
ybGI2X8n9Im5Bn2we1O/BahjQVYvjo750aIoDwuisp1eabRu1TK+GXCR8jwFRbF2EdfpD9hFgbNk
A5d2CWUDmycVMMCmJLwS7tEIDfJo5DppjqfgMYqjNP5T9pRX0HngrMnWeikG/MkUNbpVOwx0KYUP
rb4uKFkQy7XczQi1VaqvXYTweosLNECw22sl6VUWLhQDVwuSA4bcOW2u5C+dvajduDkZcHI+HgMk
3annQ4uI7WyOgtaEBHNFKUoH9gE64lNXH0/rv9A/2+POhFMXlA6DGilS1JpxWZpsaJ9mjZ6TZlIj
3Xh+YuHZQzeHp9yBf2svp1DiR6cPj89p1a35TEAKKZUjHbp2lx2H+1ZmqzBJemVz8DPyNgeTrFBG
C2pA1YnH4eiix1ZBP3lY8+rn8Ra3lWz/qCLXbH8fF5h/OlaLGZrAUhOd7uC7c8VgNKsx2WbI7Myh
auwQTei9/D+KrkZjAblKvSj/SMaLwjoDwUMR7TBEq8b3DObjvPwpeftjjJBazM+np80X56AsnzRd
G+kZU3zr4tVYX1RfIDSAYaOfp9bT887uC6PHasSdoNXlpBT4cXDeI69CfMsOD4CvUH9GGzgTbW1k
XcZn5uji30+IqPaeQQ9amwEQjvARzauHiZAkYn6uIp3myWSxCrCLtu1MeB2Xii3l7frfOZKvklgG
Foz9Qkep+TMa4tLImz1aANshWShGs0TG41HyjZq4puWjvc36PCIrv1+fGC4rFBTvzi6HkTht2OoE
5wAlk9m1PWt3nlyjjltyxhWXg4qoU/hcurEtkMdCu79BdHotF3aJ2frdwZAElbUw31LwL71hLmQL
m7lv6PG7jSr0S0VYxSc8DCnDS39Fj0nr+n4VaWN7GmswNi0UE7wR0fH9fPU12ywWfxSv0ym4bPJx
IOc6fcrNL7Z0jm9ZPPiXkrXdfimSZYnDdbmFZo+FFpqGpaFKh0LOnRd6SNpbaR+cW++QCtjAHJku
x/zS4Cc1IohUL5pAY/LpiNj65QH2KbxZjSOpfKcKYQ/Kx3OnzFV+71zR1gjtI1oKdcgYHj6OZAPH
h/dpMhdZXYNo/N1Nk+GfQj9/Eh0sCy5deZJwzPFzovvOO0ToiwLLQL9eVbjob8aQ4bg4XskBfZQN
hyt47RvJu2P162QCxduPxh0+IzRO4j4SAjkzdSZlMUFRY6T+UgGAxZysuAZfRJ53mbIfBufkfbDp
jVPdr2Co9VexcHxRY+wA90sfycLjtUgdmCsH8ZN9FHlXZWVvM3OFiBcyM7AMsJIshHE/K97n9nLl
KDOZ2oMG3Y32oaki0GY9PZ4+6Sgsm3rImLXQiyoeYrB1QKfpvmUTQ6pFwajxc5MLHonT6HMBjwRw
OCaxBDqZUkx37FNDieVv2LKej1vMeTgLFbHBz0AP/WjTELFsz5j8m7jhvhljxk881+GUeCgLworH
LaUfbYYpmQXw1ke10bqlqHwH0Ts7sWVNzsSdsWkndofeaHxdRxZOxXTd7uazW+fzI+mzRCpM6wMh
S1tDKMJ023TfKHhg/0Spvp15DBwCpDfSB4uBcACyoYD0Jr8HUU2hUtus6uSfWg1sC4ejzC9VTFpb
+p5oC8INJmOI3SZP+LGD5eU78Y6L6Q1pB13Vu17KpqKQGzVpSL7ZvtpmUFcdXDwnyomxgphcXR4A
p9T4tjFnEP11Tm3IE74IuRgYobEb2rWIDVfeMW1+wVe6EYbkxifsVV1eeNjn6P9NzADxn/CTC2K0
4BtkSsVuXXn+fdVrdthoe//H/jWZEX2LKTRa/QmiKQSGXWIrYnU6o070H07b0zcMh2vBDOO5t7Tb
VDyhHcSxCY6hYPGwmVbVQYeW8GPws+U5vDriIlJqUqXFBII3x2Wh6zyb5Ysi+gIuX5yvUTKrxLqe
42r8FP9XjBsdQKhj4/WDMxPRuRF0lUpVYPgRZ8vDMQhYa4oThYfXE7j84nuiPeea9YcZhDykHu9S
0J1j6x1IRAlkE05CLlCvHJfEA9Tk8ZWGD5ax1uKKNkzgP+JleY7EoZSWbFogyD72555SQU2d5wdT
A1bLIBLkxP6WODmBRjOyjtflELL3BJarOL9w/jMFKk/SpiUMtNxkXt2QvWI/DfOopC7LIeq6Yq3k
0XwXRHam88v1MDJ6PDf6FWh00u5CN5av7qezO/HbVKWU+N+u8hRYRKD6BU0FOkcyrFMtfjC9yuSh
Ca4TyiWY1EWYL3XfnqMvBJQQNU4ZPsw0vGq5FA4p+4UuYl1tt2k/HAdPtAPIZ12uV+3eORG3aCYg
ioOuB0hyp6Ctz+QEsYT1HJEWbUmSd2a31dri8lCaRb8g61Z9QfUgvYGgG/n0CzcjdEuFk2j4haGH
fBVZ4rBRom+j1ngsf//gGab6ekpy1CnSThm/owusIxTXzEe6PWJsRwQZfiilUdsrocDe7TtZpE1v
n6frPRffY0BfocIzXqQ2n9t45DyDpr+wCf2ge3PyzwSvaIJV5rH5vZf4ZHl/a1EUnkerEvDfA6q0
TVd5yiDZS7S/TFA6Cik02q1t7IM5hdnsHcD3SEarjf1DKF2rYPnZdwpxv0d1ohXFcnkal+UrLroh
+XTJBDt6FsqxyWQsbwjBS2MWN36L7sYxJclnrOwIdKdiSlqBwNEe1/L20FK4D3mD87mXKTA8mKVr
22mF3hBLfQeKhJ65YV8XlkFWNXj568r9khy3MffWYBweDhF8rJKmvcpDZ6IJ2F9/BH5s2+BfKMUF
gkHbZ3VFgQjLSE7Wz4b2QPzoqkzKMWrRRgb3H/xAys4+WWOVM9MCE5URROmt2wlGxR3EbwwV/t36
sefpNED3ied1H4ZU43ATGZU993J9bXLaGnGgpQOYJVF7WYxg5/kdyBT76xFHhcTRfG7ya1Oe8Hfp
fbSoG+ukfSeEgsfLXTYEscHIWNN9vTIBrj8+sq6MQ+5g2gQh6gNfbcUFvZpzzakhiHjDZlWgLQxk
tgRKn2a2l0QToOOMr3gvnJr3W24X3Kf2r+Pf+CzR0BTJ23yxi8XIE6GoZ20PIHZmXdRccmDoDFaT
lb8FgC0QdrOBQ8o7GHeAHlwuKYZzxMiva1Auc1tW4BfIfTaSfvrue80UhF8Sk1G2Ev34rEmrsYyV
764MJaf4LOo9ZrEVsxLiIVW+14sTJucowUjePCyA1sP90zvesBLHue18wXOlO4LBiB/o40H9LJbX
XkQd8W26Kjg6T8Ye9SvmaiI1zH5KdLUyIXqeOgkyhJw9TmA3J2V1EXUc1wHKEM2ivLDff1xy+9Bf
+jpOWEbuXj1sZosWR57s2ecnVEM2GafBr16JW3ABjOgBozxlvJaim4/F/Hnli5CXgyKoDkuGfovm
vwMdftxou9gJnlM+2kw1xBjOnJGAVIesuAWnQ0dZxypseK2hz+lpIaLNC+0q70OkPkzwGcaA89Wj
v4IPbZBWP3ksUbjbaGrmDidvgZFNNrCQ2YnTf8e4nPPLbITE9og40OT5sZV33R625UEu55bQJgpe
LpThoWMrQuxeWPmUYCuoGca1+UpqVU7bYDLxhKR0DYofKMSqSv0GqG/5zsr16kMqlk2ZrIDBOgrv
juJ/O8TFc3LVYw+6TKAUg5G4iUDz/7kH4RRkcScecIXHug8qK6++wB12Y5Z/iCHHJZ0oW5EH9nK+
sDrJbKrJXPWrC9P27KQgANE1dOYfXf1GpFEesAhrD90S1Q0s0V4O1N78Jb0ItQ72A+/dUgrY3z9U
ho/eJ96nbVkqxUvQj7wFiy4s40wehH/2Zzj9/k1BOrq/7qYi+1cLRNF0hnMRwKBOshTyCrlDkpEg
Kt4rOHRYjbcLqrj8tTpHIC1Z1z9FXePISgDVutDmgMYxDN4eeo4TWRbZfFwPyJ+FxKkQrXHtCWI6
9ihYcC3QX8jsAyyl9GYem88GqZOr83EnyiP2R49CYEPC2pxX2h/iTwVDXORVcG/L324JCthVYenb
yigmM26xUtYat24yipPcFBMBhcYjEpMCh/AysnnLXYcTPt4BhS9ZJQpUzUNWGHPHX3CmCrsmMUT4
RGqt4HFTql2y2x+LQD0wqeEu5XUwk2nTMKM9GJLroglmRF6nMykABL9vvUXU8hB2COzo6VhA+9Al
bR9tGwRSCtyQ4uWzmyBimR1XjEe/eQ738vMQ23zcQF5Wudb0ue5g+yHrNQQvJptu9Pmlg8kadksM
Kf6c4n6g8PmHuZhAVeT0qNRtE1iOhtAg8DguWQ29/njyFsE0M79DHYirFp+luWJMlqEqlc2hBYNo
yZ8AfFUq7MepHyNcQQyNO+q2f6GxHFT09X7WtLwKrg3ddrLXfjvPU+r2OWAFTDZ0RsERSCXKdVRk
MvqiAKDYS+rhRhbLf6jeGxjvGhI/5rHr/IR4XwW0KJHiYajCzckVkql6BIQ8Hnln+P9EjPOEtALy
2ub6XbPHyWendhQCWwS41vj/H5jyyq3eUJ/V0UTwt9Spgjo8NOBRUWQ2YZbwAbVbWopG/PCLEtB5
WQsDN8fw0BVuA9CWlQDtptTwqT6jCV48N1JZH7XunZ7M22ojcbFgFIeKS6HlFlJ2wjs0sTWPagZr
kSRCrplN4Yj8WgQ5rNkLdYkyZ6u71upQyFxTDj7G4fhNUQEtZP5fmva66fVuRGgW/y/Ul6x3KPxa
YJ/jd1GFFiWJ2YGqv/EqhG7DsksOaUxy4lDMetlhL8MB5w6dSqGpFcGT0i8deZmMjKYcsAABJaGH
Zv+cHTRq7E5+LXqUmD6hneXtPSxwdNFA+pu00rj+bJWb5GQhCE2hqFg011B3yYI9tygZANlt3lZ5
P0rOF+hO/LwbOxXhWdgxVTqsRaBO43wd1Fn/u1QtZtVEcFjtUqt8xqyoagh9dh2HLDGGXVY3hf5n
YT9V9dMmT2ROzNRqWqOpeE6lR64RtmH+08ikni68azvPGePACANTQUBm8smf9xTK1rrN2sNIEmu9
32NcZB/OC+4lB8Y85F9umsZ7ngJYLoqBiL11Tk3jKcuNlzZkNKLGKfMNAVv9W50sjuyfDsuP+B8P
EbjEWczSqmv8ECuype4QEPILn5KePnsMt7i4ynkucUSb+9DKg1Pla+rp/KVaCGfO/uk9hhzsaqwm
MRMERuueTYf3Llj74b/+73/blSQb2T78/dgEr/XOZM+A7EBvsCahmNUvQVMxD5dF5moVEItkE6Mi
K2OP4cUarDZC5niCVHVt2a0pVT9Jeu5sd8t2pPVpX0UjINctBgOR+7uRARBxLCb0LzBmbJCrKSUl
nzg/EbrNgRvIfuNSbPklEwmlBV1mayWVeoWtaHsMPoEW7Ea+LRkfL7CSXNkvlYu3YMcunyqV9Xln
66wzMQ0qrEfGh3gbgFHZc9LFVIAglRin8L5shcWSHpSMQP/XM6vUAO8T13ZJeU/WxQVYx/k710+i
54iXEIIrt2QNo6u4f5YhwVX+GxvABvcaNCp2a6hES+0sqnU3rQ5dQdn1jUTG/KdqWlywOyBY/ktH
KJveiVSTIY6YSf+QdoWV2PufLstYyfuID7OUtbDaMTNpHhJIEH8TdhIduk5yOtyokCJzG+1L4opR
DrMLjxTRZOY9IZudttZwdwzH+wMV/d0BYtTLtBGeM+4zcdL1yq82aHGnJYfgcUVBi15Y34rDXKxN
bpt0TMxoCL2WcsY0MQSsm8U9j3tzaYwerm7PityuHC6RReyo+PoKpCnMczWOLs+fd8mpOEcxAUqg
2fis3nmGod6vWI7BECNkd14I9Von8hNIwvkheLT5msYB+q6Pe+eFAqbnKqGI0Zp1XYVT+oVthNG5
J6/j5LyYTVawEz8ILujRcy0cxQRfMzoRRBxNfa6VhPIDO3Y8BBjPsfE+uH8LeNkVO6VKHz2gXzro
qTfH/UDq9YtR8k4O/6rd4iBe6J4t71WnffQVQ1WLMU1ZSe8h9fqlvT7Yddg9EBhybH3olqq2bd9y
LZsuzCCLscA58Wk6JNBKYD8n5UeOXz1s4YZmrlhVT+3Kr03cxfGIbYDxYOk8PG4RDY5cSeVSw6ra
AaDstze7pHymabYOymjM4hzXWWadh4jcplLVfDkoWudpf+H7SEAUKeTHRMrNYwHhkp+bz1L1vIz2
qLYZpLBbvDeb1Gj2h8WfXpGxufJKTk011WZn+Xixb5PIC3RahoIfvK1N80OFChn4ax8r4qoWMbX2
rT8qCx6hRLkU6Oy9Qx1EY2l0X6WW9Jl72eStk0wjhuobeLyNgNs8StCuUK7Ca4TAZd9/ls327wKf
ALtaLq/ojld3y1bk3eEh8RuA+kby6XNQW1j5Yf5rgMkxuJJNHTqmD7Y3CH7zdPO29LjlssJWT9qh
xciBqpnguLGsCmKEu4h/vvHmZSza7PBQ3J/pgxCo0E78D6esVP9tHq5+kzujU8XYBzLO39+74PYm
k8Q61XNd/aOmIsiqtxZpZWyg/wnd1eJtrisEmdyFvas/0mc/8Mm2X52ujTqnMN6JaYbyNOl8UIE/
SGmfH5AdqaSR9V3kpMqpXA7ZX/GmLTpNI23hUqymXKxylA4tgRnzDtQA3wWOHmqsHIaJ3h5ubho/
6j0jEporCQAT41yO+ecyo3cH2/H7mG+R2ZVxtiSx0Ek6adgrVSnpEsE8kjp13uxZsAkuEQCaJpR/
BWimiwn2OqTSJjn49IuiDYr/3h11CLTUeeLb6kdHKL1fNnNAURBfCLJCGD9gqskh0bHe2Bj50k96
2tt7H/Y0756QFjo3JReiTF9YlIS8RGSN9H6xt7Nj6YFv1j147O+i4Ez4GjPhEhAwAmr9IZBG9bFe
k8APOIl2H6jDW9lNE78uBCNj6Mrl8H+Ri2z6tfTR1I67FN2AqDRHGhpkd+nk8KMIvLTiZBmavQ/h
bn60g3IIZVTicMhdulxiOOV5HRVdtpwtljBqtsE6WmSg7DLXPWrUQmpcb/D9daU0+TLnMnc35uGZ
93revzJ2esjIcqrwj5lsPeA58Qpqz9JuwbflQESVhxFm4xsvSAK27dCz3R9b866lBFju1V/vkMLm
8iFqajZ3jajrD6HmwzDpRLas/ZGCqGMkw5gEl1Hr9z0IGsaQKaaxYcUJ2B7esMhG6VcNT7dG7mOx
hxeUovUhNyrC1UhDvN+ydN2e/Z22CiUA8e5EV3TGlNfM4RAkBCdIuuAXEkuonbwFkfnHpnJIqYWH
iIZi2U2qRVy/7uwWGWGXwxsiMihQjoBIDA9MFWdD1JkonW1oUY7tXrc+n9E0z+fBdg6OKA85EFEL
Ob1LpZvy2rHIcTOkfdd1/ix3odiwyE4He5Egs28kS4ZvwWbQzMLZAEPL/e+fA4LieHgcQQLA1CMp
Wki+RWthNqJTpV77GFiinlyHvisktZvo5+bw8R3FI7K4eirYmrZndFFk7EsFBSHk8XUOGzKvTSrJ
rBTJ/0+8pUjuMZhMDnlCWUTfpvixyIRJod+fzQoeV2CW7ii/sgKidquqqJJqNcPzQZPHZje8Xhpr
JIKisfEFNvRlZluE9TDKe8CROXaJNLYhT8ZQc4mqBMp26RiTkNi/yMshpkyYUM4oWPLYB284pnOp
nGnW7u6k4zkFs8wZGPNnAeqlMMYmbcMfLAi77Y9qCNh9eZUFCCHiF3aWfEuTelswJoSUPTnbTJad
13X20lg65q74PHVQ6UFk/Kl6S0Pvwp0NvpkgufftC7pPPRtU+bifVMDpTTTPbYjkpFm7kkw7L9Sl
SCjO8VWEDuhaBKx0iaC9ocqufCfoIQqNpG4luQLYW0RdZc0e7m0AdyGn5+bUPF3/aiV8WEala6+7
k+CS51w62a4Yud8k3SLNJPJJEasAtW7N6y3oD/MT5C4oE/+DIq32ce97VhbhpJRPALP0paLFhRtX
OyRGpb2HN1jWLzk+xISbO6grJR4SilWt6KPkuK/mKuIxLD26qUeRaTZ+wng9NRc1nVaKxjVh5Th7
RA2FChFdNilfXUzHdB2swUJNGzNUDSdOd/vqzCbDpyiafYwDCg58Act+9FxS+aMYE9j+MscPMAy/
3hGtazmR/1r0hBk7vhY1k4uA+clCTAmmthwlVmCf5jhB7IpVqHbMChFDCZr9A2TyaI+SHKRq0rac
TMhf9U5ydH28MIvzBpnokbTlG/9KAlMQ9ZrM8H0sk/VBLFRnjbIzWsSwPsX8ZbIACeoRmakTlrC/
ZlWJiNfgvv9VnFjxgcbo7/uMpVV89jM4g2pZTwl3W5t7iNvNzEouXRu+e2f/hvuNZlBtIAqFpHAh
bkVUA54aS/CYEh0swcff5/iqL3VqfND34ut0CZfc4YRK/YVOtrwWtcPBh+vFRb7YCwTbkJHRwm3Y
aFmZp5iDLnuprhXVnNoJUZnwO/Jr7XubnOBm4Wjuwbov9IFD3V7SFQiBCWF4nziqFc/81iY05qOl
nuRnaJ+JjPvDME7Ba/r+NZSjGcHNgtuyOzEByDrxfY37WCndcQV0EHCLOG0q/RylUI2PlyusnRUL
dGNc46MxyY9/9Cg8IC1VYrscgWTzyNBIQCVbW/B7y0KViVVfWqD+tBVdDeEq4qH2i5/lOhoGaoA6
hAHfi75ahzh76PEF/dVUcHoFI7h8fyqqtIprmuVIMthxVUt6ZYHfvWG2ozdhZEEmXNHE7yiU3o6W
JwnDETVrJeNM4K26/eI5P8KGyxs/CJoyDjhwCSYz030K/wu5NLoEL/zeTzTqiiW/3bCDHNEsmAY9
2wOuJZLXFtrc6APEiANPKwLQ6pIrA+4p0SBDIV3gZkyaNbV4dwipHvcy6mQytwyNYQ7TzXmbvjHP
+Ael2vDv1DgUhil6MylPATVZ356Ale+6wHKGEaGT5q+whGxL4oVYg0zgbH8TVhe/MV9lCSEsgCWX
qPCMVlxZMmwJY2+KgzBliMVhHnGeKxYURVG4jOfubMVEwRm/OQHz6FQZIuCJiH1YfcdnVbOnUKh5
QOywzfI2QNHSaN7gDfRS73e49jDW7xgmL3M1ZGo5Y8V9aJLA8qaUUt4N1UZbDwcnWaQ9tlD+94f5
6Awy+taQR+lQwdbXXTIh3wNMYb8S0mu9fCdbAxlBYN95WnGL6PTBpluRkZOUF3ZmboDWBbfkO7fj
kzEALwnkdDumsjJf77BRuguRa+txcicTk4SA6AX2Oc7pM25dVQchxbwPHnThYwPCQB2AJl6Ime0Y
nj5K5LQQC9jNx9N/rmRWpUtgRNQYQ0hIj86aVhf3vJYAnb20Vm96gOdgovsyDGMixwBcgmIdhH3y
tyXUempu6kki/LfOCTwkm54EmH8yiJVkMtqntM9wPZ7eD47EGBL4WNMfhZFou9TXdV4Q3+D0xZGp
V48KsYHQIPHwsqov3zHmiQAoHUC+aUVGSy5by2RfRSB/SaBJeSF9YSTghdR5vRsFCzVwRDN1+IEn
rK5Kbsom0eIjcbXyvJMQB6d27dE8vAn6kMfOXW3dYMBmZTDp0Kienhmn2lPM5Bu2ahXP7V25uqAt
oqonjRJ11Zop5nW6dESY/CeGk08XknEIxzQ250mCVNAKkmaAKtMbCMwZNp//elxcYeBlEOObCiX6
Ei8w1Ed/njIOuWHp6Am6ddqCbVIWRzowO7Z70Iq3RwzYJQ+STczNot39pVtGdo0gHs556PDufPR4
lyWASvBP5fqs31aGVCXUM6kseqo+95sqEutv2oVEz7UgKDOm9le5r3mNOpd2o+OHnrzMQJNBtQC0
aDEe5gvgtpbeTuFWXhD3wd6ozIqUEQw/YH4cnml0JYkYWi7LC81ypCQ26f9h25urzxdQMdtiFQk6
vxuX5UEWgGKQUuir1szN/ntPYjCwcjDxMYrDkzDWa7XbNKyYFH3aWZuyzLVLPVjHYAboRVfZGe1z
J8NTJggsBvDJn0WbO9Ztu5/B6ITkws4Uqf9X4GzEnxUuJcpbCIFkPsBXErIIMy+Us/EyeBgn/g1d
c3ZiMZbYrQWvQ4dgkKi3wMkWGG5pPFv5Ks9JkDVDtCCdQoKxsRgwpE2os07VcYwjiFLyHttOThVt
E8A97fwexCS9HxTKM/M0lck3zMZRNpWNyMGJ2gdvpLzKFEovJGyK2cUDrvOK6Dc7ye8LT4q4n5Pw
gguJIfleSFPC93RRGX8Qh4xaDNCr05Rpn07F6cuxKtMXpmkvP04Mkt2FyACg/vENDyOAIpxWReUW
m8gT6z44QYpZizJmXlN17ZrLn8sCYH7wqn+0tgRcQtVudj14WvDFy8EB9Srg1e+W2xTiwFMuAGls
/TdRD0CfK1gx8146/7C8cfCXZH75lwh+9yAqdy5wdZWmVCMvucVMqqm52/2muPNTNuILQxokkTwN
sXEgzV/1Ssc2z5FnjV8jIPl1F1h9/B2Dw9QS1OnK2o2c9KUIVLPCICOneW7jlrVTodm2YoezVliu
yJQA1jz4KaSpGZN1PzdvFZio1p1WQPUqH+0mV6CjoY/jLUhVpsA/xj7d7d+mp6y4dzeomxaouw+M
Ktk62ZfZK9hJ0Vi2r21GeZ5LHniGy/VlAwN4QvyN8BAg7x70hC6krcrIWYy9hLBZFNrY9HGTKsTn
G/0oGhKoG4Xuo86git9fHfHhs3HSEofivIHTTxD2ATur+fQ+UgULIcx/8mxvpjuj4Va1ypAwvk6U
kqQFjWGTvMjEzLUPvoWgE1B3SOu2uhisk7jsTOiMGBODMf6VLI8eZv/lmRF9DgYOATquhfnkallB
10KPJWEzRKPZ/MuDCXedrLU/pecl7QxPrwLaOPyE/pGh9egdBBinggyPg3ZqJgCHd37AVLCvH18z
5KLNltS9OjvGOzRviMv7MrwZEVPErvcaN/XG5jjRa7HWptRjgIOL0xy8OUKL9jDgdaCnzMHL1caA
fj9BfC6X4b9nMY1osVfau6wZrE7o2f2au9YkF+rpg1Gt5Aksl/JF+kmFGcN09ekFRcQqoVBs7xkY
3NPDeynawJE1xk43/bdGC6fst4aHjw6PxuR35b1o74akmUkiSmo/LEQEY2V9N6H4Y5gesalG5hJk
8sADOe563Eco4znFv1sjbuCmFwGopr+rnj79W+mAUrgh4IhfB+HE3cGwXWYYFShvtQzuICdAF5bQ
TNinUyK24UH8HIsT5UBRRDCC+GY+7OqBEYq/gMOwavir47I/ellkQutcacnnT0/LZMGAjIXwrOcj
wr1bz6jo1497Rn67tO95ZFnrLu2ImOWWpmWA0HdZzjJYCHmVCgve6AT3QZ0E8h8CzgAtlqf7GJYo
RXIHUrLbp+9iq4xHN0aqSFN6Mn7OYOaaam16OJ3AX6yO2fHhvUfHoNPwcrEfgU3PXQVdtEO9nORQ
NCtGYk6qE5Tj2gbqTqFuuvk5fCsvsmuhm7CsHoINiC2tdrFaPTBpLPyDmMBwR+s6bX4xtKOqqC7f
VsYnwM7ABVd7S2rwg/AknPc8QxJupdrcMmOvF0YB4C8tA6GVL5FB88fbWmU64TqOWiRYrDSIhw47
vLKhFZtyAQ/TC2fd+GUMzOcWTa6Vh+INsX8IK+liGVmTkC0gaCMqq/LWBa+2/ga2uUdIH3u5eVYw
Q83B90cyqtWA0JLViZoYPZRkFbUtEw3CQuoli8ZBifVYdujXpQzH/tKzqk46k+9VZ2p4yLtdO3GA
bA/AmLmjKS009FbYVbczoC0F2qb2E6Z2s3g2z5AeXWulC3JM+ryt2ZHmiKy3kDgyba7oEmR3Dbsd
S7iWXKpdVjtA35gk30yHxkcT5ogMN6HZW4SXHfPr96LAdZaeBObxIeKN7TdV9ObAaUBFswtzYGzf
bURfgWdD2unjd+WoDvv9kaVg+J9+LREYc/2G9i5z3HD2eg9WPTUxGtSaD76bDjRpH8pjnYWnbiDn
iUvo+qM8Lwl2Oj9I5mop8qbaVPIwhhnWvLspa2iizsG5Rf+WcCHNdgusPiMto3+MeMvbN7NiJ313
3nQCI5Jass3ujS8M3W//YOVkwJ1etPDBymWj8VJVib4MeuS1PC5YlCwAG3dFfz0g/Nb/ATGXIGDf
9mlp1ebJNiRMLzZggyAyJXtBimptvWzSYCgt9vBk1Vzp1oy69fF1UgigrYcNJ1zTBOVzhWbWEZwB
92uy1Aj8+LqTx79AFSlTDE8GTjDgMK9NROGHHJZMGfAcEz3MuE3/5e4EOlFA6hpndFA+WpuKH1HE
e39UWEspuqIN4mTa2zqE//pBNXEOxutPGAXhSMDHpEpTlqdxk0ub74z9F3JTiixjgwQvhcOeSm9h
A91OrtEwGbKKGVyQo2x+6wasVLuojkgqauSBI8Iyewz8fNddhBVLJqxb3yqs48mQHSX5gS5niznR
Le6dAl8/1zHvsCxf5uzy8PE58xTxKD6iEulv/D+99yXfK55Rtz0zlN1N90tRp8BoywF/vPiXm7+e
JoNZfP5ABBPO9syzLswv5aQ2mG3ohw2Q/SFnc6aZHN3eZo9Aqf2uZMd7yhzVSPksUqf3jqWe4APB
6ldoIQKt6WQJGPfTfpQtzUcu4jc7biNvLeprjI6clROrRp6aEhor0a3ofXn9lyVFNrsa1sk1HyT0
07vrGqQy7ux4QdkiRQb/fCsG7TlyP6KmMTtV9F5MqTyR99HUoRMnuVYXqLfZn0RRJGSRmSMKcIiC
p45s2g8XUyQVuvXRUKncexS2zKMxw8hHbUx0AL4gBt0V4e02JAXN+pa9vyvb8gB81peFDFVQ+xqp
jaVpALOaiwTJGJ0XR+Ez/H5dj4g4Hx8uJ/h0ZBkjKYmfQiifQC3pFoTAu/TBbxtns4C6tkTIKT77
itlL3sye+WUcGwomxYgc/VmuZTkB0HsH3GvirHSvmCX6y5NBHAUEMrQa27EXSF4KZqaq8tZri97F
Rbgnyof6K7CxokLVUeKPMeyTf7nvlrs9TaIWA+2ZZqaW4wMsfEECjXHI79KpA5ehQnl4dZqyZ6mR
PTipijcDbWVfVVy2YL9BbWXFn0PVh6vE92/PLn4uajIxcpYRYVLVJpnBBUrcscGxcrN+mM3Rk/Tq
Wk+1zEFcQwRJWdIqs3u4Qmp8WJdlip0Z89RU1qHQgr0Hw0KbQuABqL755SWXbmBMN2ddvELCvMYn
8PywxE5t/ZQLYrjlOTsXK1Pn05AQSrap/QdCCwcy4waJoaVEp+67xMCLu0ni3XpBLIaZ9TwLNqh6
LYCTiV4vVWrStn2+l1wv4LIAsjkYkX/Z+0LwKZBuEA9b4SlLcOEI1PXv/et8NJyvo9qvA0qcoNP1
lilRAt5WCBvyqvjPl8rKmxR7xjFRZf0Ee54dpUllCYWnhSLjS4rsCOhmotUNuzCY1GHEwQ3r0cm+
n2VOaVVBlhKTlSGngWjA2Qj/UY1u6LK4YkAcgzTEL6Km5Cuvn6h6KpAf5bUXhvlQHTSIQAG4m8sW
vumPntLlXPNlJfZ3/TYoxzWVEsg5uJvhH47/H4a33ZhvlttyLkFPkSS06rKaSjKxECFBjJSWB00a
YfVCC6bcvFVLdbC607387HGO/UXRWvBbiMHsApgLDrVjUuuHtx+ZmIrPuqvIw6moDz3WfyKPrrJf
E4BzOTkjrczUiKNaCiNr/eXzHj7OYmarEmZieeo+4eKoWlpxuDt3yumLF17lkxAwYPtPvOf9uR36
AjS6GodlV12p+ABToa29zSa+8wWcTNB6gz75IwIWzmxtXGf+WjfehoMorDrfg5W4n+On4cMCkKE3
QJ0ePpTUBvE9ycDpZI+rHDv9xN7MOHxqAVFXptIKo8EK5VTOYXCdE91Aj2hMtJSoTfJstY6Gzkxy
glkYvTZ38tRSKES8inhqYbU2kurace8EOxzYs5UNk9mPWJeUZaBBMidp1IYHWJRfMdf0To6tKJol
HNPEOyX0KJUCa5wtZQLCZHRtiEgeJ/cdT+YbQjRwhy1SKl41NtOddiRjvAufJ3Zk8pbA7KSyfHeT
222UjiKqX7HrAwkv0APj+vQR57fhco+JBpi0fJyCEkvSOTI1KpM1iBtvRvFAM/gHTzHDxWO2rZh+
917S2dCY4WjObIwcd2yTU0+Nbr7/B1gllGftDdFDMSUc4j0yOyM3RgDnpY4yNMDqo8u9ODs1HCvm
LRja8dMFbZEJqJ+f7fXdqrAWawRNt2wYgzigwwlKcwzH5MpNu0nuneUOQucMcAkMiu7X43oHCNPC
TFy0XKLhHhKssApqVBRdoz8dARPPlRre/N2k1IbZy6BSS1cAU2fWjxn8OeNnQYBtBrKv3Dn6uLCT
kRbuHFIdGN2guRkNAJ//yeRz7F5Sh4VzqLPDZRDKqUZ8dwepNvDTO830Ei50Ff4pPYsZYI6EqRED
TJh+mgukjqOXG/mpwH7PVDemnqs5//ZXHQjiwFfhFVxYi3vssDdExuW8ndnJ0DLrlBsAfL024CGT
O2FxbTPJrZelgNsRMSM1Y0PF/s1xrOz9lYhZ0Ei723keErozb1m9/MqqJmH/jyrmQhlHEP5XGBiX
fq3y0z/IiZ+eTCkC7pg0Aicm6+fDrWsCgQDAyKrzbenKCHUvY3Ah2+2mpPH7Ue+11XXDG7vEyzVv
OAX0d0sG8PhpE5pf0RqryI8qaISag0f8AlbpS+KtQB2qhKWKF4IDkKfYDFmBguQn+rfIJaZP9lJp
0JwVwfk1sSjkBMSawzNcyUiA9awuhLjWShGbJfte9WXkfHg12216pFpBI0GrtHSFc7D8qtTVhu0V
CO/ECZJVrRCC3hu5WnlpZU9G8kOQdXPP+CGJZNCQkhk41jhxVh2JUo3JByHie2YXoqPP+W5xk9kQ
xIHKwzbjFNAYkVjcGpgfDrMVyfaAUoAuK0dXgln+b0foTJsAvZCzgErav+bmwHogWL+M4nYnoplK
S4ZPo6I49JpeyfnRuaAemZc6z7saKcFSdpPueAUwdilh6PGnCAZHASpzk8+c27aWmbz5/rQMHus3
soRLLDZSCo5tAvzcTU8XP4oTedp+VkvJ2d1/UoKQQUgUJn+BDMvhbLHtbEJR7gAB/FBrPZIUs6S8
sUyZbZhXb9WB2M4eAaYt7upCCu6WlCPS1u11SLw8vJCSSVWG39CFyWvwqjqV/EVYGaVuMNRzW9bg
Bb7qeSfe7Qz9/i4H2OITzNAG0mOx3b/SCxrGI481Vnu4rY8UvXUkMAJcpadl9GOeALV6NJovrfqO
gTriCnIKTesCaEh7IwaTLcqjVVH5jrhoJ/ZQ8X0THjDb5lOl0E1J4Y8WV6HRQso815+vB0E+Hfka
IFbR83hdC0/ATmi3d3X0v1Ya38BMYLmuB/FwoPg4touNyu83Q5aybvMwwRVNHuShJYoWKRuIz8Yq
DirsRHyB7akJJ73gqcz28wbxMpaLuhmSmJmHsCq1J1KpTAJ8rlvgwTl67YrG+ZnYGlYIZsyt06Dl
OpC5c4z+NQRLVFvBBVng1g41qNSPoM8AtU/Y3eg7/NN7x9b6WIrd2qFqTyZPE6WWWnWqatj1O9v5
LbaTOQgXGP/fSQhF9mc//9fAq5RAnRqBHQq45OlL8dmNI5QXp2ekRoe/xQ3Z/t1ywdedwpclw7P2
3CQQTy/IswyEopgZj194V2B0WU+XdHnsuO+VfuezMdA6DG1K1zmb5KJ5SL67faBiFxv3o7ev1xG7
DTxDqEjYlpG3WQGLvAeN0czmVq3W+9BdQckakLaVPRs2dKinVoQ31C6vBqV31ICj6SHG9K+d6Q5k
WO2aSnQKJmIN9pQkXycM41U81ZPPwV+XIvvYlYDzKsqmgyFU8+aE0evF6N1+vG7Y0OFRT5KEo9bX
wWxqZnQ9BePq63zxkzFgE0GkTNxq21ZaBJQ+78xqCVAVhdVTPG0CwnbvQYshshFn/cgGZE3qFYq+
HI8fFOcuFgAOWE42W0Cs9SzG9LpANCQz/zWRYq7WOPZATSpyE6karbF06I2Lf3mNUj9GThGvj7q+
THilk/VTxqlSpX0ipsIaWsVIpCA8uPXbeSdGCf6LPAkorwtqQDFZ5W4JnkcSY4VTKT0d7vyx8c9w
QY5dMooaPqNlOujGRYEkdNltDNkSWTU5qcGesEYatZoncT5gnJvyzOTZk5ws+qLDqyCaSoJ0DO5k
7gGUkExazyUW4WM7IbFFRDgQPxeSW6TxUtdZel7rzQhhkbqyi8jaL9Y4VBdBo3rFAtxGngW75CC2
+l2xtanauQ1vDE1LCZhugTyYajOn0OJB/L3JIxwBz5IjJ+Shw1Vw9DuxdkGEcB6SutqawzJQwnyI
qV5Ja0hashwRcpnXQjMiJ/uPVswbGrZkVwrElkT4hQ2OJz2jOXtUV6lejYSYHA6V1RKDKx9NW7jF
sh6Qqa/xNo423x8WbdfnqqTquw3nj+c7bDm3GPpLi6qNTC+v725KRxnExt6KFpPXte8x4FWA0V2D
XhaOZs3F+VTgpb8O62Ts1u4IXZe2bGZNPN+fLxB9whmXQiOw8dbeb+NSLpx/C8i4m2s9KygVuXUj
S5ujTXbNXD8Zm5mDDv6zUbBDPP0La0edZTOhlkUHuG0z54jiskBZvgJBHsWQb7Z/CaUZCBmXx5st
sBEVk55P0mKRI9TdQBkHglAmR4+z3D6w8spUadUMaa+6l6Zg9u6jr4Ys0GRPr+bYIv+R+vt6ZqN6
k1PVyKDfP/9W8pkut+Zh1QhskWhBrInDmJyjgqNi74LOlKXQOBdtp4lLkN1APLq53sSHOQZ152Zz
2HRLK4lCeCjqBq7AQneMLChDW+TjFwsLorZo+RK86e0N/qUNPkW8gEE0O+ci847gV65pcb8G4xGc
x27pJJFo+YT9PD6S4Bsv8xBuxjOR02HiOXbQE+mX64EGV1YU1ST6kcVLQFMLFns1143yU8R2TWin
7O0IV2DjHb+TLl3QsikznTZ1UYhVTpom12yfGb0gFhDW8LaytWR6iFfsLQ44yT7BqAbRtv/R95GJ
+52ailmPkO2i1hmLcRcOggF1275PGeun2sgWU5sBqvIVe6UkKs3YPVyVMiadF1fP7TRngccrNarK
DL/tjtmHK5bJSGOCAYz9TlXElHqfZYBXMDuqeyk4lOCA23JABV5j5QH4ZCwWBZXwDu3yeW8/jG/n
w0NuXtCaY/A0BAmGl5wKbBK3c+rSQ5o8RLPfnFvR3ZrRjvr1oKkJreF6xkMtv7bJyeG6FIiY42Ex
WAxMtZcO0N9S+L8WoMfpeBJTKwp9n0cBYXaY/EIqLQiPbVmXdDv8SnKvWvXMEq0s6+n4TkXBXye2
qs3wAcE4Kz5QYgh7H6wTp7xRocmsAFeR6phJb5oxmUPh9XOBtTeu2o0XmblacVR9ZLS8OTHRSDlM
ygE5I7ru25iAHK2nN8tDQ1zhaJXqcNv4hDtgvPMXt6Zw4V5tWN7MVBGVF7qgdZSExia6tbTBFcY+
VUCWdK/bySn+3ng8rbvexyKhM6DJVEBoFL8KmFt2WBT5wgyxzXkoQKP6lV2fvydRedCH7PEQr2uZ
aE5v2jQ+5A1Ly+8WfGMjdBPzGkbb8kZDpakTGRhAOrF4ibTErrgBhFXZiSnCxynHvDDvJGGh6q+R
gTL0HCWniPJKdbGzBClnz3sVrhafkYCGyAYjsNh2IJq83jrfjmfV4eUWux7B/9M5nbQqSXYZDmiN
VMSeFrBHB7dVGvtlMDHZ4WewDnqObNj3bqJuTvIqv6SiqliTv1Mr4UAa9z92Ev6qvbg0M1V6GMxl
r7y0h71hAPreeSdAk/grFQ7Va4WCpFHgSxc7IqCZPnEj52a6agElv7G+HCII+XDt0vtVXAi4mc3u
FLrZj1MNLtPCNmxD4oyJmitM/Ay1G+Vvkb5nP1hsjZkmJqags7UhisSNKzTFWEBMtcJSuJhV7QBe
wCg7LA0ra2ZbxP8ywufPPb+B8nu5S0gTg2xS1gtMkkdMsQzjtvI1Ja7pYPNoKTFoTjgJge9irWeA
UbJ+HKQ3+mSW4cr/QdRkxPG7cQI7pHrhEUsii4iyuYlu9R/JPtgYEJiCn20p/KDsCt8q/nSfulTW
PxHvyZaFDkM8qLb9n99WnF2lwi4MWR4vK6YZFQknplJpJ5PH9ZZIY6L4E9QeFZBJYIn/yBTLpV2w
3ET5nflyv28u4GBnyct3EIVEska0TsoWbNj6pPh57+IzBnlmitLunDqp2vabL3z2O/tuEqOu1OQ1
xvpJoL3MKVAB87FyB4RNH4WzclZBeg/VAGglCraJMU0oIkkmocRfwolmBspfaAIFFvPbV2Wc5HXY
D5I3gHvlbb4aE11dSz/iSNEkmnIyvwQAlf7osXWAy0/a1oR8n0sIjKPWSmwKn0XFG42IPqSxs4Pp
PHgqdvxIYWnFNv28/k6MxZ0hFh0maUfNrd/YepnGKDOnXtOyyGKNC827mF4M/vK20QKn+OFfE0L7
Ue9AkpUMjQzGfr3xWOXVsy6+dWs1w710DGXQXNvt+XFqmA5JXh6s60vbXQBWgUq0YIq45kM5naJV
PuJvkAwQ9iH45ixtK43LpZ0JPm0h0OcBY9PLmWDEbdhy3SgRHPNt2MtpmR5wR86QYGqQxTRIWXpk
rIfiNcflYk2y7Py+Ma0vNopQmCzgiB4uc/2XU9t/WfgiQJg3DgjGM8Ui+1Zx6TzzrL2QLwLt/P7p
qXhONfeLmJ/kgKUOokTPx3qhEoIjre0mm0zAbosb06TCtNhAhD/edyFa7EdjAotk3suMYGEgZa+R
TmHZ3rrVDJnvddm2s3vifMm9AbNVdGt3Zw4ZO6jhLCFjG7dT2QMT1cvhCroa+LifZNX2ewbXrrUW
OThISy7qh6YLhg2UrpyHwkPdHxY3FaKR2uVmYlQSp3gbNJUMZ7aj8GuOQjcH6DiIOSrALFl+YpZ2
t4n5HNyBsNtVXAYFDJNPMOWU/0lAfzQjyfj3dkA3BBnvj11XDThsnqA4D77sIKx4YaSdITlCp89g
ckRxoiLMBdlToqOV8k/uXVp5e0UWYQM5QxQFLUSIngIkZ1wxiCGTQewwRuYuXC3YZybgeI5jhYzY
/p9qaaZ/HMawa3GjxP7sTR3pihD2I+NxM8pX1Oj7n0mLkMIZtD1ZOmjtATAgbv3Hh+A7JQl7DoK7
9yblUGXwDphICfFH3ViPrUPTjBKxrK+NnQ6P3NBBeyOpDtPjNX0/k5lPxeAgVWr0GG/QnNi3rZEw
U5lnBEITARz3A1DxkN8TOnA4XARiUtb0SnC4toxLyYQjbCzBNgBgSheN1o6HJEaNjz0X7pNbN/cM
SgYsQqFZdJF7CmoTlaaPX5hf+uXB4O9eNTDEm/z2cuMVpsHQ498uyMiFy2x60cMyjH0zAdE5Nhs+
8c8xZ0gOYWO2xVfiKFZSUa16f6+MQ5t8qM3rxx92QwuJ4WgBIUG4B3/KsS01KljWK8PnIp8QW3yN
Qs4FJ0ZzzxpeojWZLqLTSSRrgKR0qqZZC/XkbFWtE2G4sOFuozZQ0IQcbgu9HywxYoPZFZ9X5JuE
40cYoxjRpm7U0/WvX5Au6WG8OBpL1AnBMWNUE0KXna5MPSgmNNu97Vet36WhGXrdWFCf+O1v8oen
UcsF037deDWP8OaiDGMJCkStKygjNGR3H972Dd2Da/WCn0ZENx0pHrx3QUiXb3CR/s5wLxK8D6zF
5I8/1+8wjnMDmlxGq2D7a/P/oXGGhqJ6FqSm95qmd4aoDYIU2glUO7vJp0rfnfuImM4bWnujhzRi
mo3F+yIICGUfrGakgTqMGvRn9dmUBwzoFKS8RHZNx2I0F4QcWdPnWufK6PaqmIBTH+QnJa+wdZZD
ngFTOHGWWAc3k6DLsuvr8hoKsz+NWbL6ve7undupgecIwKrLLecZdCccHYd1CrpuyfG0eCAKjcW0
x1IKHjanQT9FGCNJLU7CPyQxSIGoywNkUlSooHhktOlRMhfJPiV3AK99fb0YksukgGJZx5Layr01
puJuxWCBUymwosDmaPMv0UhhbyhEn6jIQ7Jnu2xBJfcukhLoHnfyoxSygfjMsb18fCDikPALiGuK
ZoAJpI1Tqhwf4YNgImHvnUhNRBi2Gw48Igd6+/0ilqpG9ODABejKYpT7VLelRk8OhUMA2L54HLXy
5U7tsDXVf7WeAWDnneXehYlaLieZKh2sOPYvCKjTZ2DWYPq63/ueQlsjQ2B9HnBYtYk9aliG2zUK
Q29bftnTAJb/P9tYfOVSpzvEQrqJYRSpJ9yU1fKEn2FFEV1eoU6P+qwsaSFraXGzt4JiESycwFNh
lfladYAAPZ3WmBkp13TXcJ6OKOtcs81JAWyVZgmyqaP0yn8TyTJgDk55UYHbxxrHDDzBMA/BfZuv
TZjDKPDOO2LtXgW9SHcMZnbR2OpAuzP9kcomtg1iwUsmfarBjKrR8x4p2Bad/mcd8VDdQ/S80eeC
Rbgad8vd6AWstJ5dGl64AYYVwlyHDwNZlncU1+Y7b9jwwBxMrZu7rt5W9GyGhtbNFTSo/hmXPgIo
uAR+xY7az2bUn7VFZ/L719febuREH81hji3mTJxTLGxcR/noT6gCVSPsotITWj8q4/6fBa5ZmJMI
2sSB+ko9tv6CjWISAShEUmRLJf4Oo/dZISBkomOtI7JS3vf//cOePucqYVhkE3n43hv9VorgdD7V
wALRPKPL6ASVDpP28NfWZ6curUfiGHp8TcST3C1SjrsMIePxZMRf4Zm2/g+5Ay3T3kVKEMHVFVNI
54xJXdnzsFpIEdbMbuiKwzy5SLXhwHGJEy9AJNlPEywCtP0JBae10Kq88dza8XuxnTMTKNd4+j69
WIXyDhiMgYeu5065NsC8tK8icHxhMgSnlRnWNW89eprs/OAuw1b/ivPJyK2TEMxtAkTVdMLdP/2N
Ms3DfluPQkmJ4B7a5PSby6uCLqEjCjMmcwEC/fjkMfXlhPnK8d7EvNuM+zfricSbT/bVLKboLmjO
Jnf1rLuSvkNduGLKEx2/E8gE6VbbTpp9Vb1XUfR7Aij1uLKESq3nV/PW7xqlx8NPPecNVzGD/mtL
ETog05t3SBKAn++5MGRF0/GqInOS8PNFojs6//E26zEeZ8kxyUHkx2xkWBIkaH/8xutltnSuQwR1
TF0Rau/7L0zN2U8Atuyn5pdvMdt+h77DO3cVXQ9s59XFk3d645OhXqyke9FdwIBmaj8UbMyz7sla
KYy1E/T1hhLKJC8LHV67A+e7gQBFJ5KNnx8uy9dchNy6/kcqlQ6aPHMiU1iZ+V40dlXRwnI0szHe
kVlLHAWonMWHPHIK892Tbl7K4QjawUZYwZVUuxn0kzqW9vzbNJ7mcNI49SpAMD+mR2KB1Ie5nX+N
0Xg7LaA5X0D52dZ2hOZEmpZbikRN5wgMevCyyiwMUSju+DNt/gAx/64oO6dsi/BrKRr2fGlPFzMe
HkaTljUGy8tdpY06FqiarJYoPSDaCHVGY+Q2pKZlOMOCauV0LFkKPv9wi/9za4i4OuAnjccdlF2f
hVCZ96F0qFZ56Q7ghp6WuWbDl2GgplJ1JHStJtkZB5SQbccWJafpTiozoDkCO2re1mbN9waQ4p01
lT/ghpP49t0cA7pLK9fzFiB8P9fDrdBCyLwzWcNI+d0orHDGhtv89iS8Ns9nY++MipfIi8U/HBrE
zgUlYpnhNwcCE8qVI1mcsXyaaUOVdWGvBUu3RN5dDyYjWmGaGkaJRTqolbyRQKNZLVq7nwS30m1b
fE8WdknVFp/UVga3LW12AWdOFyK2Tnz5l21RgCBWGFauXQI/pUCGna4zCmf3g3RSSn6PJiaOK3Qs
91jtCpTFe5oPADwrGRyLVHRfshGtLuqDH10afOqKJIEXtYF5uqVm++gv7iharcGDD7RAQMjY2mtv
hEO/c1QN6oQWf22cL8qCG/3WUgCSzlVzsmLJBZmN5YjwVcaibmCqn1Wzg0UP5xeIEXrvomIRqXSx
9DT9+kISbs+9o3s41SI/fhMcAxTWw4ZJiYMKJX9jwwpnjpMlTtxCbi+VtfLK8j29+RB4cxkwOOPo
6rqjBo6Gql3TCtOMfu0lHO0gV7iqW8ehoQAnNChhTnV6cKaQGBPqUFo2v8f37RCp+/0mydQRWlZv
04LXX9nhbcIDsRALFO+uvhaCIRWlZnHemXVRf1KnrRKVJtRSCrL1XLQLkIY5eYjUROyE3MnOQ9ci
y+f+FNpxhS0DMGfLU6QkLzROKDe10JexxCiUyu+f6E+F8V7CyaoQeV/+wCXcxC0BGfnLjFoYv0iH
++wyFERrXbJPU8BRsCB8WZpoMf+Fv1Utc536i3m968vM6owslurcXrfQV5hMIT+3062yUZJdqCJ4
2ovL/gq7T1evInYifMQiyvIQy3PETev9c85Oe30AwiNACmF4VKS+nNqJ7bWDtCNIy5suOtste6qM
wyF44ejs10HQYwZF29DZKAXq7ydnex1YLPmvVg1jO0044u/GM2x/uCzbR1pfIvhfykacN7PTx7/J
OEdxfltv7sAVHNgm2cHqGYCETVbGa6phssOqrVZsZw7G6C8aYqpyFMTl0bj9tj7YBL9LHOJA5rFS
L/i3IzBKVLpFx8IVvdO6u6C5hwaJqnn+PNJYi6AR//Q59qjAAjnUxyM83gdWnPq4zvtccj2QhT7N
h5d0gMYg9f1uQZX5agOWNHyk/C5Q2ckyhi0Dws1xJXCY5Kcu1c/u/ae5PxP5C310o+QVYW9O3k07
z8bg+QbKVhBA2p76dyLdNcUege9J5fANCLvQLcSdg4vSrbbevOc2WUJSaJ93Yg00vlg1CEauUWlc
3DKsAXzbn6WTiFF+huJtjFXAuQ0Sd5XPxagpPxptWU0V35xPHxO7+dR5+LA+ErQKPXmg0SsDfrUn
T2vBLGc66hbvjODdlN65t5JgQh2PJj5gkFxNE67hiQzHVwhQC/yPVXSCxMORkBDZvm/SZEWcFdUt
TQY1pqDQZ0CxE3qZgRO6AsOl99KqEmRAJnqV9KtE2hVIoptNvTWrquk1hCzZz2vy9KhAfUSUvVDz
f8Sou8zk+4nI7QQHNFr0BdF4mBsFZ+S8M7NSVn9ebUy2ma3u8YGfRA9Zg7UYq0FnR8d9TciSFJSR
kAtuYNUkNP9BxGrpHsi3rVwS3QYXe8e5v4HfhtvghwKz72f5UlFGLwMh31+7q4cu8ZXVUNdE1l/d
7nlRRWJQpvCPD5FbKxCdN14BEE1z6kjDO0MCiAPBr9RmYS1slVyA3fE+Z/Wcelo2MYnocoAo66n1
1nZspY4IobOqW+GQuRm+QYoi+BxUiOOcGNaN+ZxIyQQ6MAf/KbH0yCra9ImXfXogxfWJFQx0/k5L
qCVa9fl7ahgSeZSy2Jp9usOvx6xtIBe3YFLnszUnRcHouynM3+hItEoiHsQMyymERj8zTg5t6LXH
U4WhX+CvPpMXma5Oe7M8Cc5/AFMm8sj4emAIbvWCva2jWxUrAFISMV+X0nBQ0H5U6irTbkdVMKtm
Bnkw2aEHvqupwqfpiuJg7nDLIjugr4Wry+s3Be3G2NChSTop6CTtc3FGfft/EvZRqRBz4gIOLXZR
4Nl4EiB1eg1wZ2gOfmfQbHqGDVFqVydeTs0r6aLKF31Ncnhs6zgdK4qT81gF2G1rO5H+LE1P+HDw
oH6pymt5FylfY4kvoZH4ZozEZ62S5ynwk2RtHD0AkyxUUiBx1uS73sg5jee5yUrrVtVbR6W+y7gD
IHbryEGsirDJfzJVehv5xv/g3yaJ/5qTgnq+aURSeOndX3L0F+9IPW/wNqxMnIuTmsH8tHGKapQz
gkVeJCi/nkSbDm8dRZFFDEa+2q7eOY0BrH7qRZRE1yjos8wQO+o7ML544j1al4tMV/hyQH6GuGNk
j+KO4ZTq95bMAfv++FLJaMchc2CCNnHZ1chL3XnTOotGeEzxKo/jKmYeEjC4gjEWrRAXEq3GStHj
LRnVTpcb0XSIDIO3+o6LJVAoss640pk+3bZuNHnXVsOAf+d13z/eedalCEPajQFirkvqeYeMhbrL
cZhTEVoBEW+JWLBsWDBQmNITE1NpaoET0BuWsiUUnD6ryIYSDaxNupeLDWnqdMUGUnTH1B6XiQLt
YWgrLwPUHIPGpBOXZBjENhPYewZnpIURfYo0J8ShSXtK8Jf3pF+c5oSAjW6/EDA5Zx3N0PCLEZYs
Jj1h3UHG/GxcByXY+L1l0f8HqQGblOKSo2UVtHbJ9ujkY9vxw35QbEb7yvWjwNMGRanwVHryvaZ+
C8Z/CkqS2I2TPVKhSSGEx/rRavA9jmF2VbUWYolzxTednGfuu7iaAIWOS7RfdDyx4i+xoNTVrJLA
IhbMVMrhoBo7hz7Lumtc0hJ4Bv6hz4uXA8fondJVdqBzic1H8T850mrKEnK/RSU18/pCr1cxNVCh
ul5NrEkicRUnkgLDmxmNUBI8uK89AgXNUVT/y3fOwdw5J4UuZbm1ychklMtXB8afVdtXc6kSq5A5
aho/ZgtIjuXlyAjjANvrUmRW2xCmdz523x00nliw3qs0SqeX5TZdY/VFiLmxqnSyyD8W/+k6wkfB
TUXn0+wzBH9TtPQ0h4lSjJVgBEnRDQT8bRefHI3ISrNAYLGJbDLBEGAoCsdmYu19mzaaVD2QUeEo
dzKPEZMsKnSt5UDWsdg++yLUPrX9PbWvynzUDEKGXJXhUhtQIZzOWxos556MqR5Az8dVPeWDqwFf
c/7gbR9sd1L96Jw6y5Y31UvgonOuehegs1Y8int0TziF2Ndz3lfitaUT3HaHsFfKuPm7UNuZfUuR
OIxMJbbdTfYH34pKzgNG7gjlWx8IxZKLj72hSkjVbr1Omww3FRzwSlYv6/layMWILxpUTItHLNnt
UyjofQCb8iuzAOfb/THFOI92kuBnB/GFjlNxC8IMRz/E7bwnkYbuS4rHZmpsWykf9JX5zyRi3ZEm
1HgGuuzyEIX97ms4j1PhgMaSOV2ZkihKV1RTY3BVL0iFSU6XeBsU5HyUg7S6pU2+m9gzrhGCB1bY
UDF6zgsnfKHFzAwLZsg9Jjpo68Eg+OwIcQG8zwGZ1r7iU2M4fuZfL9By1QiE+Wjr5iDoAD/Kv+Zl
+K3RfqVAWvEacSL71e2cJJtI19bbCqbgCTOD+b/2jmC7cQMxD5Gdy20s5n1RdAbU4XLxdtllRXGK
Pdt4fmwtzqr+r2ra1xHpZAlFZ7RfSJuVBAET0lEGmDLiJMLQxqf2rcLzqNFbSQ4kHefTSVCvfMyI
27PNKCm8xdG1V6w7APWjjGx4masKRE6nM6EhhAHafooQwMSddEWgoYCBLxzE19qdIVxMHbuC8WpS
af04MVestBzaAeZELLjcREICbJt94xGSJhO4gNM70ISqodws67swhPftuD3I6XDe2TYEklAQQMZZ
YetXZ3ZNIY9ORKRqhma4jK0jvbelGeivslSPFX1OCEW3lpHwsOiZ0u7OFLyWG+vE5THdrCYGuDKQ
NWT+6lL2n+aQlmcITrPW1uGt71cziki59bKEHBAHawgcg7qVTffTLgIdM3TdERCnMb0SZ4/vVIk3
ytt1tyd+GqUyqsD4IZHX3o0ilKA+fRD/TD8HqsFt7SVGJTX3DVS0xXSTx953DJlAZeCGLYgSM0WX
6LMq1w8BVPrF2zwEO2X0CKpvv7Az4yzjITj0uo5/W7qKGnxv+Nf3CdLPtCHvYhYlAVcr1BC7LqRM
Fh+oIS35BLre1ivvaHfMW4XFNrqwCP0/ypmcT9LUbXGDWBq5OmxWYvtnfJT2/4ROVOfvLMtVP+UV
27QFCOt8huaunA6j9qSywVs49+7pTNavyB6EbtwD7SVDH60j8qFgw3Txo4yWK100dnsSfftaCg4r
HdJ7Dy/lfLyovvV4/py+7voQ/cetRdwfsSKT/rYfCGjsKNxwGrlgDoCwHedKqX/7qRgJSX0+mGf7
kVQZSt7ce9ebgsLhILDYZWSizKU7h7TKcvHV4JTSdY1/b1wSxfEUqTDeDU17Nm9IIptS/99qJIj/
uqqQeoeuHyTg2sNV7QBVx3j3grsZPnCgvgm8+d7SAsxzG49b3WUIPzej1mswkF/GpCnqbR5+kW2C
3naM3V1ECXJ8wsxnyphaj2PuaHcZ07GcWFbwI0ubDkOVDajkfJdWk20HvoginWuk68VJE/6aP1Cv
MnSLalEPJgM05QzaKUTvVG4dkde59Xe5g9WlYYcOyFUeailRdWgyiIAIo98EmypT+U3KlaWGiAZH
bSdHnA4dPTMNgbED3eKruMEcvY/Wa2RK3rbMlt+GT8DOEWGq8sm4uZ74UN1PAbgdOnKM9tlFg620
nvV0ZF6JfvyCc6D6RwvT2KWPi0jIftugpDasb2KTQLg4Y8asSo0FKEsHDkTHs5GqI0GMREMPIAiq
oAusmnYZcA62CCB4SgAndOXmk6q43/iw3kKK8J0TZwDwyUYhewzg3oeuFW6F4InT7Fvl8l52SDb9
daeRwgIjmkitPHKR8ptbdZgUPdglDfZRcF3RZDkPb1bVGbeh3c2qqUVtKVN1tB/OQlX5XMfN8VH3
6y+mnGRtnj3q8kE4LRgyWyNDpDmjm1x3NIdspdPqM8fQrNgJXedA1HAMZ+LB8P8vrC07SWFaWzdq
2m5POuuOU18aeHLPNYvB+p0VBMxIRhTSaxjf5IAfo20tow/+7aUMQ0+x1QAwC3Vm+rgqhRqn8Q1+
o+qxErU9KZcuiTQW7d9MKtbVQ5oiquLfTsUk3vc1jsuWkt/x7VDbAlzyH+ejFmbAKJzcD2yq/Fat
xfqOTJzJfyZxFayoZR17TleZTS/PJmTA0/WTn2+TDV+MmP80C6Z/k7dLgt70aWJenw13LVVJHogb
VCyxiBcYrjjcaN7FpkSC0wFUJEHvVqE1a7NNYKpY9XuU84kK19iscW6SxStPkTI30/ENkFC+x9dE
UtrpuY9zuxNYx8xUIJQWiJcI6uyv7EUTjTgkLyHnT8yL83Z+zcvlpf1Mqj3aIe26NVrLwiV4ryPH
DueZfHS0VHOwP0g+MYkNGxQh4Q1XXK4Cfg6ni0mpYqRcAWm+zs7ccqC29BN/eBfazphG6zNzaqXj
gDoEdUukbYqMNnqbzpEI2PAFHHyYAI76gLVyaCumB0qHUX5nLb/Qno3dFUEVodW51jjfSqho3c3l
IkNEe/ceq3PvU3BL6fANiQe9ypZSs52FrOgmhoONeNsap6WbIAETpOkRNtiDF8I4OHdVomZGz4A5
bimQTiqRdiox3J3VoJiLLfKoe2xk8O6KBuRFdH/y+7OoJeIY2ptNJ+F7HJVDRQogqyQLMDpPgYNG
fWgdq6SeEREhqDqOIkBYE80UkIjPG/KVZHQkD6iyWqasmhJ9rD/G7x9BoaVND1qGqOFaNVBghaGu
ws3ZpPcXYljaRf9i8KNi5PmX1Ak+tmSTJMyhHONp9asr/A6gCgPSeetImnu/ajrvmOlDD1SDJHAB
EXasevK8EaTqVdOEJV0IY1EgNI9eRNUTlsKVDbe2OsUbJ4Hu/1CNGoi7J4tFS+mZk0okh0OTppJq
9t/US4uUmvQdRIjRwNSRPNSH7tp7dtQeflB4MniyKJ4ON8bO6gIp8eT7vIk8z9K1vVw6+8nd80uH
++YFgoeT2GpPLTuDKtmQ6F0xzWdP6Cu/JBshS4Wg6hoB8U5ah+x7K2j3jtTNu1vfU1a8ehFCK+Rw
NGCWm9l3kG+gYCJEip43ocoL9hPyQgE6Vq+1/ErLDTxNgSPHVIz9r7cPsA1z2w7GMsSymzQzyRrZ
GtildVuKyBjCSaMWTqjFxsOSb38BuagkavYPH4AhIQYhVwAWmvvdikEatLPAnZODAFGep9mR6ujf
I2h+LboKMalILnEgFMm8aKfH8zGQKMCbTQRLGpcCys1DjuT4jUs4ElXHQ0csQrw2LnSXCYw36o6e
/D3yRhKfaWdZJprQUMRIT9A58/LOkngPG3nVcg2jRrdRwRR9WB1wvNvJHh+Ezc4g4Lwva4uAdN8B
ea8H/aO/wffqwSqz/6Ihx/LviKGdCJYDjIL/7Ma5Ane2KxNyD1gmOusYWaKqgd095CRPEwt5YqXD
3WtV+CqQKRsbysWn3l/nsY25M3vMmKrrLPyRHXVx29H0/wUHfpcxrcx038I9AOSOm/bxKww5HqFD
VKBsG87HVNF7PHiey5/IAv7tHt5KeyQdTZgG6f5dKpuVDSHPfh0ZBHoGuTImZ6/egbqcwVWfm7l9
CuEOPg3dHwZS47p48C1CvCxkKxjEJqqPyHN1dVhgGi25X8qxmU5dRTWQ0WXV6RzR9Jkji8RIwoi4
cTwlWvX2Tv93bJyXZ6fas2Ccuqe67u6T+4mFVqwZVD+Jj/dboF012l7l3RvkNWEUcVpjTRfAQb7P
NBTWz0CHtAG9Ap9e4ECZGYwHfiFTA5TEep6v92QxzJuw1C5Oq7K9QlG/ZH8yZdNsUqOclhaoUx4v
4jO7u/j63cO1sNc1r91TTB2IuBk9AANEqSTumvzel4VfDeiAfndfG7tjSPRsdGRUl/wgx3Bpp18v
4u4IkzG/wC8vq7NXofd5WGTEvsoWsmrRu0YQTFGPH5N4xD3WDYDF36Umz8tWcl8JitVHRajCs7z+
vBu1ijonJABCrtWrrCSMGc7zr2CNHqUqsmSGn80gkjFVvCB1ALph4suDcjhgB7aExvP1FilXsO5Q
98OeCBjK4PMDKQ/BVv8osq/hP7Hrem7Z3xtZDH9YA1uafKJ7qUWibkvWgCpgfXzq1LXB4ZWaBcnV
SxB0+EWVIxn3Y1/E15DUGFuey9N6+PkZQul/uaCYNxwE8/wKWQ7Khyelpkkdu3wPx+8BK+JB5VIU
tlt1eARYaoGt49Co4GmZgWhb5dG7VmeeAbC5VozmirKUPXHxL59iiJfGkOMPLYShHDG/rWAYN47g
Y1o9IIf+xNWvRdjmNKNFwrjgUDXf7jinc6w+0FSpvRu7HtcVv5/iCdWKKOinhGYHnSK7vSx2tF6P
9kx3ZiZxw4QDkXNr6SFVrAlYptDyUwfiV11l4yZNss6N352JFlhBAjySJZtNFvqeP8lFI+OGnpms
0Wewf/kbG1mtWi6e3FUP14onB3fXlnmtPf79g4J6+rE4y3gDlNsxlBbqjbC8Igmz8rSmDTCT59cQ
nRV0m2gmm07LPUjm+UGYtG1rc+0NCpNAD7K+52gbZhILGNsyFTwDAXBjgnc+J858s0rYM/BcUdlo
tAKrO2KEAaJ+Zc1Fl1rwhH2O5wAw1TRHeyKXLhvNY39FU9aioQq16l3P8G6p3sZ1o2wA8zwEjQ/o
HtZxSF1aWAITHvIfFpMTRtsYRR4LJXyw3ZL2AePxifBw4MiF+Z3j7qNswCSXP4TVS11C7cXfDSAa
Zc0wKDjSxBbU6g41xUwFgLGyiH0Fnc04eIxxmAI6bMZYZtCD/G2/raeSdmMUL427BIM40eApH1Tg
5xmje156wncjEzvZo+tz8YwHBlnkGgZxHIR7y7Dux5jmuACtBcQ06ELX2+hazAitU5ZNfm6TaUca
V2RE8+FMJKoD2D7DFCIL+ERnefl5XgNBM4ABPeKHZtyv7fM4GhJwO6+PMTN8egByPrsnZNVgumpp
QWjZK+XfxUIp59bfMH1PZn81oyFxP1ThJzw10s6hVnzg2ZK1yXWkJKQlckJ+TBXelZ93UHlb6qdE
SRoWsk+eURzPms1VmVUNblJZIttL/+wu/nsXgF4U/4mXf5XICPXyzpHme3SXTXXrTXhxfmvX8It+
Kv/JUhuyW8WBfwJ64KCVrlQhFE5GpmRo2L8VQ27nEqh79SOPGCwvNvkBxA1UwpmIIrozNWC8bzQQ
KC8+yhxML7td6X4kyHeSUfk0y2Tlg5fiOctOSCToHDtHDxuLPoAoa2M752OLZlH5QEtOqhrfVwHu
V3Fn9FlOjmmeomFaKc7Lb77ss+l6vB3xuFu0waYi0nxIjgVdA58U/TbChYg4/wH3EZ/LTzmz0UDm
geecEEe6LGw2uZ5IMJHHGNvxJ39NH8aG5KcbtbGB1VmoeJxb6QuvCIa/eRbDDuDVs2sAW9BgwSZF
7822qcAm2qEWuSwj0FEgE7AX84l1tVaBRcMTL3ufq5D2DOSEKjB4Smn+YN3JBfbuUSQOqzyaZIdC
/dRoEA9qhOVW1vOoB/bm2ucMyzi3DcmvAQYyHg9P9OzY9UGHi2/0NOm0Deq7KAAqb7Rnt2qlJdjd
T8KO1ymKt1Uvm0SQyVnbB++z3sYIkcaKqFMyco1Rmh1m5ukF95yBdFiGBZGX90+T6oX6Pfw7HPyK
gCENhqXZZMV/5eebxKVPQby+KSj3cr0igw/XCM/AuHembGYUseLMYEW33+rU5ORjYdQG24bzJSgK
FvFfc63bmWNJ3RfnW5tl4My9c8xnpnI0ThQheUffr/a0d9PmkRDBe60m1VwKfz/uCUGAlCd7U5G0
jGZYDT37xcl4QB0el9qHSGusi+JW91sR3E/fy8+phWQfw8UJDeNDYv2osyz//eDafjKcima1Kwu6
D9Dhs5eqh01voDI4/iLI1GCziDqrqglHsA4QOKsZNiWaVijBEL61eB1GDUNOi2oMxNZlfIeJTboU
i0u5nB8BWmsLed9L/m6dmw1xf0TZDqByTOwl66UtvEJHbUUsHznI5JUQZT9pMN4pZwNlNkrZOStw
FrFeTOoSIGeRqDjxJ2+ip6O1bJ2kztrQ0Owi4XBu1uV99umQw2n+c81ll9XVFQFYC03AcWUvq4I/
1AlMvf83QCYTv1tVp6cf/LCVqrPkihO6qmKpQpMNsjaTkoh7jvYyel2CuEPgXzYMz27Zn946sXya
YPeNJyfduUZItfhSRxyEv4r+JkwXRkDaLzlsC5kn4Fz8t2jgniPbkvaNwEE3DmumXi3G6mJ5vbXc
1RgiDjprURsO9mHEhkxCdgIidipqrXAawGK3xKfKKTNf/PT4Ur1hvch0gfgVedapF1gwTTnS9qj9
49NH+94oOHwXDbogxwgu/+eTRYgRXHHnkJnWZnNX13JeYJooroMVOeG+0XZx0myEFB0y6vX3nLsw
/YKapK3fzqzvzTBMocEj0aYnMdHu8fDL7rmnzMS8j7QZ3bJvRGjPf9ZrEXxASOXtDAu3AIIKyX9w
Voa0e6slUGSxH3w3e5ksGWIC1DTULbtnxMapL1+Bo9B3LSHOdZwjRBZ7HguyM3Nb7mxjxnRh28OG
cElILmcXGITksqahHT+xLxx9l0KcivBBHWdV4psWatjvjmexyJpMaWW8/cFf3JJVXXbBsBIMy18M
adtUl59yta5cQBd4rZCuhm25ocUn4gEUd1cgvtGM7e8CXNmVH6c/hDUj5QvS3cEQIcDptI0/9uNt
pR2MlZvIQhbTAQ0lCrq7NacG/BPHTdk95rlCJ69lpHMBbLfOr+IoPQE4dLqfxrENsxd1HV+8Edya
elKN7ynL/xhhIUTRjm37phJSIzWscIAE4SB8R7KMKIKmu3pBJg9lataUdd1yz8/OpMx5OeZfNIDo
OSrtQq3z1ND2s/gltmsYzFM/wWmqpp9+wZg6iGjEUdrdFmdfDce+VPalb2LYAJUqNFd2ukExWM/t
RAZ8yZx+ZoMHENzlfIpP6SvfeqvNJd6ueZMGrhDbYxjbOv4c9U/4yow3EeVcKZjmoPl+0Xe/UfvS
Y9gKRbXkDp91+yacEOu8lh1wKwAgnwyqpfq/gHQFLnBVfcBkB6B1XWre49P/sHkW5ddu2ZNLFzQd
FZsknMWEjTqe6jU4z1cVvZ36bEtPX4UH0+Lh1MqbkKIkTNRseZ2ypj84r+jMj8yo6Ios0zXhGA5f
/dDpvXw7Ti3hd4yPoHu0CuYcZcbPNTjHlNP9ySpVFdPXb/V4OOcG9QX0yafFIArDgEdX9nDyV469
WyBp8V2lBzlveNphuRbpgqrOJnwer7cM7g0k4cDZ2WOVpMapkTXu9J523JCJ6O/N9+cQ02+v3XYq
qnNS+IoMFoXsysWzdKqTKLet7dazyRlDM5M2GOtSioe6BjNxyOFZy+VT86FFcHbRXhaex0o731xE
JUi5coqv3R8Qrtf2zDlHRLwRXvjcFgQtvY+/j6/bQfKjRSHUI1GIUwhGrkywXjKlC3ui2w+JmQzz
PYoVoqvEEBGuwzKLG2pY0NducFfEZ+3s6bIZwKGb+UfWIv96UJQQcFP8T4nP4untZiwu0Enm/AnV
w2eR5WQ27OYJg//Nwt4iaz75MMWU9j7cBhhfagoeAhh9qZzuyQ9KLJ6NwbnW8ueQMDMi7jOMC6XT
Iahgley2kolsoV7+OU6mNhDKsZTvA0INSno4UAlTfyr9EYXOgm2s6sJRU3g+U5T6bC8MQwkqf7UT
NJMumMo+Nyc1xcBLlkntdDvgc3viRRxW+03X+PUD1kCjYfuNl7lKZSCaIZNypeKhSIULc4Mvum9K
VeVFe1TMmvaZQWb143Wz6bgLOwWsRTIbz36LI1sury3h9rX0BFKXR0wxpQjrGe0Lu/e0ZqKZJoV6
XLvyxLezMXPssssn30FEBqUH2JPH2pS28shNGhbHvEXr2qorLXZOd/450e4EHZ100+RvVymRmspz
YKzkrcgwMkwB5uPspvWcqhMOjFg40PPtW+ulaR16bcpasGALuGwptE6Vt8rVk7KmwhMYAKnLbPZH
tMRleuw6nvV2XbOxllDFSA2P2VD/QN/apmMRfWGrTKjoE+Oz5ezQgsQkXhrm5mElRnDhfMtzm1w3
PpJkbVtcQslGqb67YXCm+98RXKi9vQT9RYH+9R3zqJhw7JiGUYJdur6C23Fa7QbF7DBz/L5R9jKr
vVB8vDT+uCeXGHTbk9R2TGVdoOe+KixfwS3HR72AEZLUcuqEL4sL5MedcDYbsKsV44wyWfQQbgfO
oX70mTqqZcQcl+1ugGbYEDkWRbOpisRrnc6CSEDfE7SzcECU7j3IConFr3RWyl+w9n5BgcDwAnEU
Cr8SvN1rYBETo50fytJNn3KM2jpvN1DR8bOUQUCwUSjzMGSzM7jw/q3T27fKKu0sulWpru93el9b
sGSMfkCn0aCppLX+Zp9alX+2bRzWORGff5cZtlu1aQGYHp6F+3eyB5HxX9SV+h7KWxiJJTvRYYir
lKm3IMijefWNiG/LCWOx7fY7CGvAneSTbtxM0K19SU47DBsT+r1xRQ1bhC8bUH36yDHNAu3GM/Ui
gUqw+OXjo6EH2Aoiqb9sVaahilMqTJcLFjYGRf8EsSfpwRdmZee0aN9RrImFO8tlK2MScie3opBG
GJ0gyabgbGMe9yCNU12b90rR9mTEV2wIAscuc9Lf/vcqXwKdHmndtZe9MQGCtmlEWILUin6YRUvg
+fDoO8Mu4WOPFcDJyu0gJuI6ohIS0oW0Luq5Ljy3yuLxqvK+SIrDj7qDqTvT8h4KiI07JezJFkHQ
auUd9lw4u77NLtr/TOgs0P1eTEwmCFUwaACsewSghbkn6t8PgoCqkYzZoEqp7Wuf1RAGeP+t0/aF
amRt/omfigiyFBF/RcjdRBHRKotyNQk+Ti/ToJj8GaBraElCrNauioeMKMSwPAjJ75ZNG5hpdLCw
fPqUMxVFbEWUcRO0WLZLDVdeFE4Iusmr2W3Y6Q8QEHxLg+i5ynqcD3u37ed81u19efGyywdLHe0e
brfUhfJz8b40q9aHCxFO0w0dhqybzhfchCHLmhCfG4iUkMokxwYYuhLl6QoGBkJfKFyCacVNT13m
aO21EH5m8o4Whqz4Ef0pesiMN/Xy9rUrc3N0bYfFGktg8Qf2EXjwm7urWy1ZBOwpmAtmog8PfUFh
8WxkO5uzwTvSw4zYbKBCHfuE1qwx6DuQLS2PVkRZuSP79nOq1/GzSqLPMMwz9I2S0O1hpCUm3/C8
GeGkopPdrHWRkX/CRvnM88An+CLXSc8I5ocDFSVpmeHb8UFz0YFc+sQj2kLHQ2YOHxhgPX1DpsRP
EYRblQsuNbxid6rSevrgAY1DcyXD0OP60IXHvphU8FclxErd59c5FKmse1ErUIwGpWe0ZxnRePaC
3x32/J/ZiLwzDJ9ug5E5DZ8Hq6Zu2ih7pSOHaMoVG/Mrpiiot7Hbg5i8hiD4e2MYlXQ+eRSb0k0I
loS490Pxfef0/2NZ+ce4udW9IuHQu8h51N6/bLkt00SyXOPWku+x6orgKowmwPXs+4aSWUfBtl/L
4+IFq2MpLUWNVwwbSG7HsUVb2+cC3ZFcwgnuap/mEgO1pOptyXeSTc085Ekz2QZM+/zxyFeCE+Sj
Cob1944s9DIJrdLRl2QBAXfYaxXHwwp6E5+4u+DTtcy2NqL8BBao43EmAX0ocF6WWNDycvcf8j9C
KE44u9i8kLGA228gsAtVAcPHUyEJhZE0iVNNrFLMZQRMR0rTmzmzo7Y5bfBz97+tbPAiLycjm/Lq
3rZ2eb0wEIIVgn6i3bH0oAQq6migol7yHfTK2/VUumlK5rTYFYeTo28uWso0FyR9xeGEUAn1mpRj
f9wB5rmgnTI5tESoo/TYYXLY67U2RCUUKSz0SnqGlbkiQtpp/vb8xQYkTCCw+gDdcWxwALxJw9xE
wwav9B65do5AQnIO6qo/EMNvQn23XWNpkkx8uYXvypzNfVizAil2fNEsYqKZG4pzHXcfr8zHqUIJ
nqTlK5mbmxkcH5mQqUajMWBwwOeCQij43F9W1g/ACxozZN9/c/Djh8eHpQvkepl5JE6E2tqu6h+3
qsvvF70M/zgNuIwh6Hzmr5sMMZbrW5el40Ya0tMUtDOm9nSSa3FZ/Ilw5XosYWxIOkW2ZreXclG8
b7LW3uxvjTrZD3iW1gcF19IlupctJOjC9tcGQbq0IMV1C9csPqVdgo7IA9QHerR4vxQ+0sa9lO3A
l088ACDF79rEVwpPbdQeq1/neoHPFfxehtU5RaJyqTqTWkO6b9W8NFt8Jq0lA9pbRz9RgITG9Sqv
2+5iBzbXmduLN0PzYwSUVKeKq21lhh4yEj+WTOOtt8pnMxh2ZkMpUWumtJDWFlsOZgGuofnEYF9r
Ujh3hOFNu9AMrt8XbjF/GQo+gEmq+JliI4pYF/nl0slPyr82IpPUqFivpwCU7cDV9hHC03lV2IOf
aO0INFZOLsX6lOzEMaJmGgD/0dtfgeqTmSe3gN5/08hrkCeoemLxmFVE9wVEVBy0TsmUf/ABjV8v
fkhsCG7xUIByMIrQbsV+am9TqYAsNo8fUoL4HzpTMuop/zIcn4kMYpIxhx/omEepo9yC7NnV9FkA
vFG1eflKBZOzdxGysXL5X+YVFZz9viku6ajmCBcGw8MQwHpb+0lafgx9izw+VKBpc9aU3Fr/Gy71
AmJ0hG8Q/1XWZlFE1BkyIijKKlyGJBOFQF9As70idTC8evqYvyC3T60B+gRA8GgGAyTZwWjN1seV
uMtLAmIIflPuWGEnIYffmVxRD2FLT0K02cv9HtLCReXeHrqySUxqNF6LJ+zgknLn47Nz4XPnVOOL
Izo+bc6Q8sVT8Ce6iIeUZVZObvV48Nl15kKiKu8ANHwc8eKZWZg83gf8Br1rYWcVJzUH8K/StEha
6zDU99peyaRp/QgQIrZRBmHWPIXnW6zrjoj6aNgsAtRnutTF+zeW8Wu+kf5omJQkYpLOSBze5j+S
PeVu6gsPVHGV7OwaS8S03m2IIHQyjj0yVEzDhxILlcyZeh4qD0gJzEpqGzkKKsqwcuAgooCoid5E
7C8yvJpIjI3ytmADHB4UoCrQBowTyogXEs2Fx1dOWy2sumvOlboCheZvOEiHWTOnqOoakQob+L0y
Ez7qts/HHqb5i9fUnMEQxGl1QZehErvldVxwHpf9qAlXM0sP1jCu423Qtfto2B+P/hf7r3jGJNU2
WvnEviMQpHhi40MXRJ1kGI3pdCe5b3QLot8FJ8hj0xmxsVVIzBueduAQ/CGQ2X3XJ6Fod9GqwZol
cYqklcynvDSVPmG73KHpqscPBGawVxNFWnxZZHPzQsepMDmCn8S9DvyKv/LeRA+Q9KPtnWmGd+XL
mYaUcyPI6dWt2HZ/d7VIzCW2alpV2I3fkh6yMNMcYmRXWY7bQ/sougQ3QOgjsaGt1j30Zi8bxDfl
jTa2noyXIUK9VSynAOO/q80NjxHde/CgYAubQkfDLyrcz8ZMuF/4pjCVU3dikv/MSOx5GFKpvj1t
jGNpRrOQh6w/KicnynA9Xw2rfCQN6ulzNdxzig/I3xQhd9O0bagjxPkupcF59XpvY3J0AB+1HNkD
upx1MdY03VQqukyuQdap7irigvAt5iuFHvE6gUAeJs5zTdRTCxv3DvdD02kxxZJdEHrEMadFFKfU
71Kh7/iuXHaooUt38P4/b+TVONHh1qnmWfnxhLG9B2s8CHdnSI+5BaRqXOXkV2CL85vW3dkny3+0
eEgsY40N9zFvozXYiJKfSKGnFRi7ZOIgoxgmYn44AlUJfbpISUoRPkLTaWU4wmJsTcXmlMc9Ph6U
pYLL4NCRu7iftYKl7R7XTsuNooPH+veeKD9JZ+DIZLegjKXXOxkQ6OFtkiELD8KlN53iWoXFWpDU
1uE0yEv5NlzO+5kvxg8jriV3kVq2h2TdMQGNc/Jchd6aWV9JEIZvpuXPC1b5zUOdHo/VFHmKt6G6
pnSyqjI+83ds2RFS/A4Fuxr3FOvpCRUvS2kzRuYtXkP0y+uxgRrRk5vHHHJg6fTRcPsGlyOx5Ct9
0cE8l+c0ewgiMW6jiPWa+NlGTVlUf5JPdey46lmQq88ogeWaEYHfvYBVwM/dbrXoHY4Fhdupqmo5
mI5J71m+NE8FIUY2/yNF/lFnqDo9AQvfiCNAxQyotu2o8VEmL2ZKptL7VobAtxWy8uV6+fYuO3MB
9FnQQhxxVxCuzH3aOb1CxgJGKX4Hr9trhwbOhr2FknhERAEDkRipbCBm+N6jbbxc52IIarXnFVtW
a4Kn04sfFWVR/X5IzZUTKzX7vXxzLZrXoQfPFudKdFcq9Gfclk0LzbkpUixXwpje/AEoYzYlBVkK
lzTuV8lirM6DgaSU+1sUQjChevR1wQy5OhdBiG6wFT5I6IkGd0gLdE4xnKJkrkiG7BdER0ss88aH
cFElKzQggloZ7pnQ58TXsCAhz18GbadkVkhXBkP80h54tez3yirR3eNNnHqjb92fBMBakhB96+4r
ofVB9Be5/kM9DWo4j48fgtPHYH+mP1g0Gd9NvOV35PquKVEdO4S0i4RqhfpMOTdGOCZY9csEKXbN
lIn0ewAV7H3PMK2wWTGqQhqWGbaaOYXizItvUR3Vh83TJ7fbmiB4xv+Fp4DElhlRpDo9qJ40OTia
mPgW/j1kxy+FBN9aZIul90KC94THBSrCh2LYZyN3QtpH4/m9rKDO/aQ+IwcVqjc82s+E9Ihwb4Hg
T3kTRb+2FEysC+vVr25PkedCpEjLGHShmnK/BXKp7glhHvaxohB0p9imezQYwyD6srnNbhNywnLc
g9JVedNaUFOM0IkXm5STs/iiUzoau6gZ5cgKc2pAESAvYUOycnLMTFv1iII0AzPtDt0xJnaFpSKx
SKjrp2Yd1MvGpLuBDPm89BGTzrTHbe7i4+MSpRmvzcxoLV3Xsw2TuRbG1YK2Iyl7V9kpbX9yJMj5
92XTm8jEyOuNu8WQTos8/+4LG7nV1RFM7wxyP0x7NA69/R9JJTiAUizJh8ae4hn7mpFlL/JlzNP4
/v289xk7hg5exN0T/sR0ZmUR9z8jDoWwxv4ClqjmNZk+OW0JZFj2EEgKBPIt9g1WWA5gyLElubRo
pLZcXLAZ6n1fMeiF2s2GYthYXC1DlTjWElf9GNQt8KIZoo0ajYW1Za8kuvXbI93vJ1gE0FCSk9I3
87kC3v4KnnUjjEAJ3i7pilAt38ELnhfjRF1lKIj4kzbNecf8vbTSd2m7NWG/elfI7gCAq4t7rkkg
7PwJn+V04ZEE7CkChs/2OBETuZbXeFhp+rPMND4QQB6jKXf5+gSJjAyhmBZendwMMGyd8FNdRedR
z6QuTeCKzFgNgPxcmi23UzV3zzCftRb1PDgTDmseSGBIzbNSadhcskoyl5OZ3phEB2TXHdm8li47
t5RJcyNdQQeFzEcgecgneSep819COTJ/YOqLnvu8rKWogoqxjwSEvILODXQU52Z3X9p6l1Uh4kUi
dOGQuwmS68QtvGMGw5+IG16YvkKuxbOAEUlzX6dsp0dB2fXXaiBTZa4uuZKXFN9OzDn9GFJIeEl0
bacAwAvUm02Y1cmT8iYKV52x/9SlCZ8Xif+HJYlvEguUZjL7k/fKhmxRe5Ne+3cJsKx0qiZt8CpC
9V4xehlTUMl/CYauBE8lH5Vn/slBPNH639VjkWgebQ1AzJ72E/wMUj9wqg6VuRSlNcCn5QsKZ3xa
IqHPwk8Y2GQpyBwvyH4kkSh6m0pgwC5L0Qx3li2sdegIVN83t51lmMmTdsa0FJsnhnv3AqoXQt7Q
Jon5f2EzP0ZX3e5KVt6eyoLL3Glq2MCfBBjXQKT3DxV4d/5HjF6ybhrlXnjYJ6NbOkdY7ltxVRVR
S8yrwhEJlw25WMPKIIVD5kg3KITvEInez8mB3OWxHCkuDZ3Hyqr0CVUVUqqVpSAkJo/0+eYLIpMN
XSGTkVzSMbaQIdPEeCQy2jhMZFVvOsBuef81VOlX293+b0+U+aXfmyqUle0bOrqsH90ZHmKI4u3K
2uyJwiDuKFYmhy4fuASvsrZq+dX6gQIS+J1Czsm5HHkNz/fAc/zlrxwpExKJSl1d0Z94RoNGqp33
9IfaykfAI54+EA/IF4x/IMaEK5nEXte81mWF2ApN54/vRNsNMPrB3cO7fcj8KT+lRBn9w3m5hPph
+HunWoGu4D5ePhHXQ/udf9Y85mm4tc5yr2s8Hf0mX2mQKTJlqFpfKrYUVTscANQ8dcfaWkjFAh4=
`protect end_protected
