`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MClIjjPUf3yfhiE+m58bqUtvc2IksRotikQaMkRwRUVKudsCE9ooMe37uEVTz6W9cSaaoSwWws2U
Cewb0t+WHA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ix0lL4O/9TR1v8ZaRnOokgRS1usxNRx0dmGdcEINWtlm0f+xl3PeanD4igVumZ3DKBEANkzDE923
yJGqY9Aibd3bOu42wjVKRQ/rXiGDTV5MjbPHUozbcLSob5dYNnNMPf0WIrdtFKLrALZ7GnYai+D4
Jaf030nznWwHDUbz5yA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pXC4GU84Hy4OQhCt3K5fKQiwx4+CRBx19XEl/TBOZCMbB0aIP1ySAxiS4klxd2VubR+BPyBuuuEW
JamVq5EEujFS027xx+l8nqqRmiG24huDZ/gGmrgmlFk2JfFW5QVZ/RzbgzKLg6i2KxNwfL1wdw9k
GPw8CeIgxjgrR+gezpQ7JuamgFnoWuHtZodiRKIzlz0pOacI0EKyEddf0gZlhdcbRQKuS6WY/jku
CBk0rDkXVmKNisj9XVe9LiQopjxRwyp6YbGYYrwK2KsUWzbOBk9PxR+70jv1NfDt5xPaTV3ymph+
g7zQKian9wbL5Aeonv0RwRFQgwrjsKkCxTfZoA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SWGIzCEQVdPJ1rd3aRiYLOdXloFYRJG6wmFlc8aB/EhDv97lwazKohgsRl7gEj11nWcydRp/Jeek
MHPQUkIqW5BU9S4E+9jiMjjCd2MLfKs2NPyoEjBxd/9fWNxjPAmFUO7Hl6fM9MP1aK1Lp9Xk9SX2
GqNsuS9rbi5mfNeA0SY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NvBxEHP0PCX5+nAHxlEPg7jHzsxDs5XJSHdx9lmqgeH7m9ThnzJKhgIuCfHmPQ0cJJswF2rPdJc/
YABIPjrbcBHfdH3yrT6lccXbOX+I6gZUZrPeGUboEjqSBj0ldh0EILWEfhQiULnFZvCDgIxod7VV
8c2yeayrYb70/dLWaekzBZ7r43gz4VtqsyYNsIMyFdzxdN6I4dk9q8OoR2HPTpkWV9ya7TWNjIJM
u5lrr3kzupQdwcdzf/9SbFd8qahg4SfAOxaZkf+EiOYmmQOe5N/R8kXErnoj+EENzAoO8wcbMyz1
zaDOfO7VlCxHvOVI9ZhwwIGCPCtuhjCo3aG6/w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4672)
`protect data_block
wv0KW971qzQP8PdF+SRtg6iIuSJStvwvojv39XD7XLdY8PpslZr6MAwqNMVRZgBOasHaiFDNRUNI
8mF/iwfMeGEOHhI9cOBwft3cIyhknYT7XvGh86pqBuVOtH6MmruRClWVt0PWPAeo1Z+md/11JKcJ
mKs5DC1uEEgk9DS0W9UHwj/8cFLKVilfViM+0jEkCMcwmqmZo++DLYCPfcMJ39/Y8SI8hr69rR1J
Qy5ZCNJTMY3UbZabQpG4m+foc9Gt6mB38/fua1z8XlkhVuvrmXKsK9s+m2SPw1+0aaAI73YD40Gf
5VJaCnyM0gzrscGTk0sePqU8PJFnAPxZcUYzmI7bLRpTNFNhY7M25VifsTce3IbNXgzRqMobFf3D
2OhA/+RuGXGtCVo+ULyCpMk5mbSZ6YZpBlDJujUQ9Z6CtZHOnSKyii8l4FjpX48AOEJ776Boe4Ph
RIHtYmvDJZF0KV4w03s7XYBVRcVSVpauqwcXpL5eRv2XsUfY2uF83thugG20ev9nnrUezhlvN8tS
PVCzQLxaP7CnsPot8ybMyZANo48oqwGYScdTD6qWczPy7TEXurYefLsn4kL9/QQQMneHt6YlLdA5
bdnKtTyYHp2POtIIyNfr4C+3mMk+Tw11/jvCbTfFqbVSCElIpgLOXxvRmvQLqTGzdYRzL53jE4Ny
RjnIvjUxJro6CGWlB5bbRpueabmrM6IuMfqRMdMez8z8y0v3bLR+5YDdYfdU8KbdWs4hZIXFE7/c
3ASAJYA1i+H8x98/VpjhcwgfJMVzNPb5MvR8ykTUdCTN/GI2inQVMvBJq2TAS0YHKiXsx0KgqRFs
IjpKFGx1dQh3smbnUqOCE+RJqR6PA/yRmFv/vJtoUfTga3I0pRclpibLgIhhIurqQZ58JuZTZ9Ea
hwK9waz6zB6m2ItoMmjW+SCtt94dDXREitdLYhh58iZUG00azVWQ+MVEsVtVc3ljSmM+cRCHLCEE
eZ5ef/rYFr4U1FBZjY1fUsPpOmqcrQNfUveyupSD3kvewILM8hMsbF6Oc4qgum2GKz6XAGemFXU7
vNWr5VbXO89aHPuB2S5fWFig+sosRoay4xAfRpMXBV3a6OHSA562/IsGwjRZdBr5aQx69bOYtkmB
3iEevKt4M9BkfJxdokEx9oZtkXKagNtKOk0cdlXYc7Kc8cToDgLmPQEysJSMbTfWjijP0VleWcOP
f+xsPPcMHOpYwMfd5/LEBzR71puc3f35IFGRLNahJ0KS+XCGKkIJTAj070lnvZMmmN8hEkj7HVEp
T204sM/3DeYXHAclh4tMYcmHr6k89pgaFF5tXUnvSWknTW5CpCBXoUJdZ8ZTrOpRruB4P2KbKUw4
xzXTPMeBhltWHT3e+XdwpbJGE5y2tDLKUkoJyZti9rfzCXRlonZ8WUWxdMY14Dm2oFbwqTSj/voM
6fuz93gdCcsJvmyAWZbM3joCdXlT4VctZzdNcXJIA3ZiKIu9ib9mv2DJW5V8cUsVlG0uDDd69yoS
X9pCcd6VOuCECujykqGSN3cdJfmEtKyeVqA7CxjkJOWZz/NyyBw+k6+4qd2Or8z2N5/8Tedd2KqK
WegpjDxGZLBe198dHH6GCoQsZAQD6vwtF49Zx9olakFIlFjOVcrHh67sa3KttgreACy/1HHzokiu
aWlmJHK5AmiXljSNjNObVcFt+xHXs3NGuKyF4kCLPVz05spNAQGUIGFyKnEIVaBrb6okGfQ88vl9
iRJZd6RNjuoYulJiCUsb2hxODtfW8b19r4Zh3MO3ws/a8btUZanst7Wj4ojmPNEXtuh0GhmW0oJi
7HoRQpdITl6F/UaoQ8q+KFU4N4ubMRKfgL/4ag/1/er+t1J1h1ydWg4MYIJcv9ZMWu5xS+vDhffe
UfiorpqFW2sjOyQVWxJrwBmaFLNvoa6GCaBl3UzGZv/L3UUmHnOQmpJm0Xz/A6KGjD+v0C2g0EJW
SMYqyFUf2fzPVtPAhYOp8jGfx3jTZgGGUI1eBRXKPJbeKj/pzygCy6+3/IzKdF3DXcJOVcdqexVC
pfTE69oigpNBjoYV9TOOuyD6U6MuJOATOC95oYhYkkm40C50dVG3XVaWnniWPdQgzfv645upuVYO
fLExnSJDk+No5WY7AsPhLHf/prX66Utfp9SQhhA40bO6niBw6cijYzfZCgXZx4Y7d29GSLTVZDAq
8YuSl3iBGsH1p9xmI4a3PR2F8bwAcGpaLpU9lLiG4ASJ4lWDdfqOkRlhefA1GHE3pVF+8/UY4El1
t0pYOPINCaGCGe5A/Um98+6+iTYRYo94dLv3ABOYXhRoy9obkvdFFmppAO9YURS+trZlsL0V0+7g
nYyY7Hh8rShGGQvjj6UYNRwMbsuvQ3jWbMzwaLP5YJ92IyEIkTuwimK1cuYYf89Rci30LqR/ya8I
CraoDPCHuQOgQDqaH5DwvXV3utnXxWhHOkvTmy6M9QTENTbAhnULGhh26f1ixCSv5uGp02gVVfGH
vXML/Uj0HfY3NNOYWSHF1ginskAsv6FLwKQFtIXh5/rqbrzv6Hcg2zS1ei1aZ7aXjBrV2HP0wIrH
QV3KLf6J07+1yB7r2kLDIQP6IX0R6+W17BmyEgqDNTZRlzhMrdQHNbtqx07YnYC/2EdZykqrwtR/
Kn9zJyp94HrQDl2169TwspFlEjGuorK9k3PemB3k4UvdcYGLijVR4+nYvk2+jrqaHWX8iKow9aal
xtI5yjQCSxmmxGQdCRIhnp9493jIiTqawXAfcchqBPF6dZ2nlY6cIrT75mSt1D1p4nOKAZdLhmme
Tkq2RIYM3K7ZY8tcCz12CSMgD6hW5OJfSiSWInBF+uyYEtO2N3vodZhm1FuOj/wD+zbEfuHpCM5w
7sSOPoetboXNkbnRRm67K8I3VyzlnnkDkvJQh86+DpMjm0hscK5UjNPT9aJ44BNHD5+Us4xxb6Dk
dIIvC2K2sGnhphEfjlYq4qGuhwYfYD4XhuV+rUtqcxWMBELoBZKrAqYbN6LCKt3hJUW4in2lW+Pp
lbi1NU7/PRV6brqhrYSR09grmvfrJgm1Nwp7+5xOiWMfPz7USBL522GoAehiUZTmeFGITrmdBmUC
SseZFxG+HgjEsZlhEKReqF2xG/vYid/aN2HcFvPTBjJeUr7Ytt0OfkbBA9sS1Nz6zIvnsI6g8LLI
RKw5ZYhth4Q3J5EAPsdQriVDFIp0VuWIgj0R3Lo8ZIzr/s1p1+3Vnb/I8xZWkO1MGxJt8ANFUVEQ
l5XF4DNOvZhQJdu8sA42YiO41b01PSKldTXY3NWYAtzTArdr3FBUk4OT1o418KpgJbod3P16iO+q
O8jGe4SjEfO1B5zyeptivO96Puf8Z5bjX8tGT9IBcCMJrP/JTmschq5hj7A8qLtYxliDyRU6hDwx
fH01Nr68JLv9ktveO/0zU6LgvxwMTNz2xMj2+/60ogibGc7ZZUnHDSpmx0PUa5zbUPkaXtTecuHz
sYT+QjBzLCVJlL1RRw2slfstyN7cUIisT2k+GJtlnmatU9WTBt+lSNRK4ZqI1bht0TVXM3B6lIF6
ZdXDf6msSmYKkwqKbYRCzRfRDGFutGMn8LpeEtmx4laKPR60Vg13zAcdsMDVOqNhjNd8izxPfn16
H+X1jbAOMZzdWf0SOvpSSEB2d99SJCmjOtP4YYdfAgztpraUY4CaEKKzk+qYzb01iDSKemRggSJE
jq0TvKNmPea8FpuTkwrfeER4XITsf5I+lvEtLrMbHICtTQO8qooZp/iPiERK8dEIFhSUXpD9mbAW
jRu71GUMqbCjScAn9gvQsPXPK78GlCtZ1AzAqKNcFL36r4ToUk+FFGWs/HgQedCb2JRHKfrSjcmX
XvfIa5rQfCwJcGkAQ044iMxRUJzmqmYmBioDkOTFRmdOpNwrgyTcQAZ48gsUPw0Ig+BmKO61XcHw
MeuHA63jJTpCvM/akrK1SOcq8PpciUW+1Hv5j2kOEae/LJH4S4pxbvDP6LZ6hfHiIbvxC2RQO9VG
oeuqMpI0jBRMnG+by6NHovoMKh6J0J2i1SGkZMHxfPoDaNTwHBIoVyUQRDQFvxaYWWSB2i3IxAA5
TTwhNQRDbULrFLoHUWpOLjzcbPYfORsekYzNjLFl+yMCBQXSo02gKcdcd/WcR/C60zqBbUF6LEGN
n6DQiIdUBasIrCoSydx+nOaiCRiFsN6/N4wcGyVj00eakbVrDSmP9Ux7ELlpnRmJI4bGv4OrK/6l
J+dnbo0fAgiMqO/J8XLBEtUiq0hqEXgPBRqZ4g1FrvPv6zyidzm7AlwdPBJNWdrivT5Rgt2j2EmA
3K1Mf7D45KFfUy0n5hvQas6JGiYwM+nPjp7cdlwqLl1rp3EGqDwaBm1ky22rUUMjuPcw8A9eGy//
VHjknDv0SupPE8EA+sk/vUwnuCJ+YlLeyrPDj1w9Vho45EeYx+8nZSfk51b7+I60cYUKHLxjLoO0
e7KCbauIsHqMiH/vTGCcmPX1DWip0nIYaVx7UBEiQp9fpHGjrCavoFEJ1iDRnbUxDr0WcVKMnADU
UZTWjyxKM9O6pB3DpBlKDjdXmU00tq7G7yB+UEFHXjP9+v4dS0/coc6QeHs5IO3QKS/UoNQOYC4A
M088Q4nuCtQp54C3BenoIWytrx9OIfHAVqAjqcWFbf7WGqFTDBE6o2lZNui2YK3GCyG817gnSHh9
bOUH3dUrC1rw/+xosYrY4HNToFJzEb9iznlSUJh3lkljb3LkuZyfwSSSpM/TK6ljSG6FwLZD7akW
oPj9P/kQh0XZw98dRsMS34H+ahaCZjKAceVVfEI0Z3JjwTYIb2kq4p51TZqGXwZjVTJHGkfHgumj
StEAtoUoVsGgsRzrX2tGXvprF4t+xO6AAb78g3s6EBzh+0ceH+v+n9S8MDbC7k63NuPzpjzaNMZG
202xrqByN4rvkRx7lsU0SnJKF+J/iB6kCTsJNnvacvQLdLontHgYgJUhv/SnO1/Cs/rAQC6GQjKo
JYCXkzXEUXA4ylPDThlxFaQAtlLqCZwMqU8G+pZeVuH+u862T4bjYvN4KLrMw67QG9Y2ICUYzZjl
KYbYWArSHNBhmKJiROIlJ15xbuAcOF+77ReNzaXv3GgzBEyavUWrwiHTd6fFvNI3meD01FiSMto1
+kmVcQrx5qB7SE8oBAIj9pbI4S6c/hy6BzIuynWVgHXpfQznwz3zom5yCERI6SDDCOHZ3klHuzAD
+vMg6c8n7HQYHmA32qkJB9t8vmTaBScgqufyoLqOk1nEP9oKlsfvuAyh3mbO2qxOx2DMcNUVT4i3
KOQKbT/p9vHtQ+4hxTaSPF7YawXZAD0XGrWAHLOXJoBBaa3h2e93GVWJMbbTqlVEsDmW6k5N5yX5
bpxdLamk2Ex9TcBQqnkoIxGm0yh9l6/B1da14j7QeDgPMYE/UWSegwXduYOhYrgWSZntwLeNbgly
jX0Af8hVCN8dZXa4F2Br6MvYgSBoHXcylXRIJWf8mOdiVc/3h14f7CbsmM31uHipticXuvHAwtbt
yE/DD2ZPnEUoEPz4C24SmyCrckIeEFBuBD6NK+Nja77kH+hR2EGVekaePiGKk3c6X2fdziJ4NO/z
FadV3wkmtgfPwGGDpTPT4iWWuzrGU08YKI/dTSpN+ybLGmFJqhkeS+BeqsjMsUv9uE1LbHFhifEd
vR4Q4HhCaHWAHakVjsOB4mG/v+8oszorp2CrWNZdEe2DSP6/WALU4hWFnFy4xdz20Vg2H3sbhPHO
nF2iBiPR3pU3EcS9mbKx3y3bEKi2TakYwaoQaP6aV1y2JDoG0Cm3bWyGuZUgA3veuAo1T63t6Kx+
hdA+hQ9xQkt95wTC/+MK5mXjWoRSAOySG+e34XheOvcSRX8hbwYbN1o7YyelrS6eJOjaQNyTh5eT
EGJ1cqxksm1JRm7Ff6wqClWmZR4RsLGUxu4yFtY8xDtGRbXV2wCIx05ostN1UTckxffOTbrR8NJe
PtDEIY7ScAsjh2+eJpZkclJxSB+jNjudRII4ct803Ua1w666KJKZw0SqHvdz9DeWt9/zz8j2GhpP
aSxE9t78n78pzmQNaHj5neENOJJ8XLwQk3hoT5YfC8PPluz9R3OmB3zxaWBwY3vHUMocYt8vC4IV
jSvJUkQaPy3Fi9wBoB7oNShAG4z+jUDtgXcttAKVdboJkqyOIcuWWzguIUlAX0HfeWw3UoSxUQ==
`protect end_protected
